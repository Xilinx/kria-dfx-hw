// Copyright (C) 2022, Advanced Micro Devices, Inc. All rights reserved.
// SPDX-License-Identifier: MIT
// ==============================================================
// ==============================================================
`timescale 1 ns / 1 ps
(* rom_style = "distributed" *) module testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R (
address0, ce0, q0, address1, ce1, q1, address2, ce2, q2, address3, ce3, q3, address4, ce4, q4, address5, ce5, q5, address6, ce6, q6, address7, ce7, q7, address8, ce8, q8, address9, ce9, q9, address10, ce10, q10, address11, ce11, q11, address12, ce12, q12, address13, ce13, q13, address14, ce14, q14, address15, ce15, q15, address16, ce16, q16, address17, ce17, q17, address18, ce18, q18, address19, ce19, q19, address20, ce20, q20, address21, ce21, q21, address22, ce22, q22, address23, ce23, q23, address24, ce24, q24, address25, ce25, q25, address26, ce26, q26, address27, ce27, q27, address28, ce28, q28, address29, ce29, q29, address30, ce30, q30, address31, ce31, q31, address32, ce32, q32, address33, ce33, q33, address34, ce34, q34, address35, ce35, q35, address36, ce36, q36, address37, ce37, q37, address38, ce38, q38, address39, ce39, q39, address40, ce40, q40, address41, ce41, q41, address42, ce42, q42, address43, ce43, q43, address44, ce44, q44, address45, ce45, q45, address46, ce46, q46, address47, ce47, q47, address48, ce48, q48, address49, ce49, q49, address50, ce50, q50, address51, ce51, q51, address52, ce52, q52, address53, ce53, q53, address54, ce54, q54, address55, ce55, q55, address56, ce56, q56, address57, ce57, q57, address58, ce58, q58, address59, ce59, q59, address60, ce60, q60, address61, ce61, q61, address62, ce62, q62, address63, ce63, q63, address64, ce64, q64, address65, ce65, q65, address66, ce66, q66, address67, ce67, q67, address68, ce68, q68, address69, ce69, q69, address70, ce70, q70, address71, ce71, q71, address72, ce72, q72, address73, ce73, q73, address74, ce74, q74, address75, ce75, q75, address76, ce76, q76, address77, ce77, q77, address78, ce78, q78, address79, ce79, q79, address80, ce80, q80, address81, ce81, q81, address82, ce82, q82, address83, ce83, q83, address84, ce84, q84, address85, ce85, q85, address86, ce86, q86, address87, ce87, q87, address88, ce88, q88, address89, ce89, q89, address90, ce90, q90, address91, ce91, q91, address92, ce92, q92, address93, ce93, q93, address94, ce94, q94, address95, ce95, q95, address96, ce96, q96, address97, ce97, q97, address98, ce98, q98, address99, ce99, q99, address100, ce100, q100, address101, ce101, q101, address102, ce102, q102, address103, ce103, q103, address104, ce104, q104, address105, ce105, q105, address106, ce106, q106, address107, ce107, q107, address108, ce108, q108, address109, ce109, q109, address110, ce110, q110, address111, ce111, q111, address112, ce112, q112, address113, ce113, q113, address114, ce114, q114, address115, ce115, q115, address116, ce116, q116, address117, ce117, q117, address118, ce118, q118, address119, ce119, q119, address120, ce120, q120, address121, ce121, q121, address122, ce122, q122, address123, ce123, q123, address124, ce124, q124, address125, ce125, q125, address126, ce126, q126, address127, ce127, q127, address128, ce128, q128, address129, ce129, q129, address130, ce130, q130, address131, ce131, q131, address132, ce132, q132, address133, ce133, q133, address134, ce134, q134, address135, ce135, q135, address136, ce136, q136, address137, ce137, q137, address138, ce138, q138, address139, ce139, q139, address140, ce140, q140, address141, ce141, q141, address142, ce142, q142, address143, ce143, q143, reset,clk);

parameter DataWidth = 32;
parameter AddressWidth = 8;
parameter AddressRange = 256;

input[AddressWidth-1:0] address0;
input ce0;
output reg[DataWidth-1:0] q0;
input[AddressWidth-1:0] address1;
input ce1;
output reg[DataWidth-1:0] q1;
input[AddressWidth-1:0] address2;
input ce2;
output reg[DataWidth-1:0] q2;
input[AddressWidth-1:0] address3;
input ce3;
output reg[DataWidth-1:0] q3;
input[AddressWidth-1:0] address4;
input ce4;
output reg[DataWidth-1:0] q4;
input[AddressWidth-1:0] address5;
input ce5;
output reg[DataWidth-1:0] q5;
input[AddressWidth-1:0] address6;
input ce6;
output reg[DataWidth-1:0] q6;
input[AddressWidth-1:0] address7;
input ce7;
output reg[DataWidth-1:0] q7;
input[AddressWidth-1:0] address8;
input ce8;
output reg[DataWidth-1:0] q8;
input[AddressWidth-1:0] address9;
input ce9;
output reg[DataWidth-1:0] q9;
input[AddressWidth-1:0] address10;
input ce10;
output reg[DataWidth-1:0] q10;
input[AddressWidth-1:0] address11;
input ce11;
output reg[DataWidth-1:0] q11;
input[AddressWidth-1:0] address12;
input ce12;
output reg[DataWidth-1:0] q12;
input[AddressWidth-1:0] address13;
input ce13;
output reg[DataWidth-1:0] q13;
input[AddressWidth-1:0] address14;
input ce14;
output reg[DataWidth-1:0] q14;
input[AddressWidth-1:0] address15;
input ce15;
output reg[DataWidth-1:0] q15;
input[AddressWidth-1:0] address16;
input ce16;
output reg[DataWidth-1:0] q16;
input[AddressWidth-1:0] address17;
input ce17;
output reg[DataWidth-1:0] q17;
input[AddressWidth-1:0] address18;
input ce18;
output reg[DataWidth-1:0] q18;
input[AddressWidth-1:0] address19;
input ce19;
output reg[DataWidth-1:0] q19;
input[AddressWidth-1:0] address20;
input ce20;
output reg[DataWidth-1:0] q20;
input[AddressWidth-1:0] address21;
input ce21;
output reg[DataWidth-1:0] q21;
input[AddressWidth-1:0] address22;
input ce22;
output reg[DataWidth-1:0] q22;
input[AddressWidth-1:0] address23;
input ce23;
output reg[DataWidth-1:0] q23;
input[AddressWidth-1:0] address24;
input ce24;
output reg[DataWidth-1:0] q24;
input[AddressWidth-1:0] address25;
input ce25;
output reg[DataWidth-1:0] q25;
input[AddressWidth-1:0] address26;
input ce26;
output reg[DataWidth-1:0] q26;
input[AddressWidth-1:0] address27;
input ce27;
output reg[DataWidth-1:0] q27;
input[AddressWidth-1:0] address28;
input ce28;
output reg[DataWidth-1:0] q28;
input[AddressWidth-1:0] address29;
input ce29;
output reg[DataWidth-1:0] q29;
input[AddressWidth-1:0] address30;
input ce30;
output reg[DataWidth-1:0] q30;
input[AddressWidth-1:0] address31;
input ce31;
output reg[DataWidth-1:0] q31;
input[AddressWidth-1:0] address32;
input ce32;
output reg[DataWidth-1:0] q32;
input[AddressWidth-1:0] address33;
input ce33;
output reg[DataWidth-1:0] q33;
input[AddressWidth-1:0] address34;
input ce34;
output reg[DataWidth-1:0] q34;
input[AddressWidth-1:0] address35;
input ce35;
output reg[DataWidth-1:0] q35;
input[AddressWidth-1:0] address36;
input ce36;
output reg[DataWidth-1:0] q36;
input[AddressWidth-1:0] address37;
input ce37;
output reg[DataWidth-1:0] q37;
input[AddressWidth-1:0] address38;
input ce38;
output reg[DataWidth-1:0] q38;
input[AddressWidth-1:0] address39;
input ce39;
output reg[DataWidth-1:0] q39;
input[AddressWidth-1:0] address40;
input ce40;
output reg[DataWidth-1:0] q40;
input[AddressWidth-1:0] address41;
input ce41;
output reg[DataWidth-1:0] q41;
input[AddressWidth-1:0] address42;
input ce42;
output reg[DataWidth-1:0] q42;
input[AddressWidth-1:0] address43;
input ce43;
output reg[DataWidth-1:0] q43;
input[AddressWidth-1:0] address44;
input ce44;
output reg[DataWidth-1:0] q44;
input[AddressWidth-1:0] address45;
input ce45;
output reg[DataWidth-1:0] q45;
input[AddressWidth-1:0] address46;
input ce46;
output reg[DataWidth-1:0] q46;
input[AddressWidth-1:0] address47;
input ce47;
output reg[DataWidth-1:0] q47;
input[AddressWidth-1:0] address48;
input ce48;
output reg[DataWidth-1:0] q48;
input[AddressWidth-1:0] address49;
input ce49;
output reg[DataWidth-1:0] q49;
input[AddressWidth-1:0] address50;
input ce50;
output reg[DataWidth-1:0] q50;
input[AddressWidth-1:0] address51;
input ce51;
output reg[DataWidth-1:0] q51;
input[AddressWidth-1:0] address52;
input ce52;
output reg[DataWidth-1:0] q52;
input[AddressWidth-1:0] address53;
input ce53;
output reg[DataWidth-1:0] q53;
input[AddressWidth-1:0] address54;
input ce54;
output reg[DataWidth-1:0] q54;
input[AddressWidth-1:0] address55;
input ce55;
output reg[DataWidth-1:0] q55;
input[AddressWidth-1:0] address56;
input ce56;
output reg[DataWidth-1:0] q56;
input[AddressWidth-1:0] address57;
input ce57;
output reg[DataWidth-1:0] q57;
input[AddressWidth-1:0] address58;
input ce58;
output reg[DataWidth-1:0] q58;
input[AddressWidth-1:0] address59;
input ce59;
output reg[DataWidth-1:0] q59;
input[AddressWidth-1:0] address60;
input ce60;
output reg[DataWidth-1:0] q60;
input[AddressWidth-1:0] address61;
input ce61;
output reg[DataWidth-1:0] q61;
input[AddressWidth-1:0] address62;
input ce62;
output reg[DataWidth-1:0] q62;
input[AddressWidth-1:0] address63;
input ce63;
output reg[DataWidth-1:0] q63;
input[AddressWidth-1:0] address64;
input ce64;
output reg[DataWidth-1:0] q64;
input[AddressWidth-1:0] address65;
input ce65;
output reg[DataWidth-1:0] q65;
input[AddressWidth-1:0] address66;
input ce66;
output reg[DataWidth-1:0] q66;
input[AddressWidth-1:0] address67;
input ce67;
output reg[DataWidth-1:0] q67;
input[AddressWidth-1:0] address68;
input ce68;
output reg[DataWidth-1:0] q68;
input[AddressWidth-1:0] address69;
input ce69;
output reg[DataWidth-1:0] q69;
input[AddressWidth-1:0] address70;
input ce70;
output reg[DataWidth-1:0] q70;
input[AddressWidth-1:0] address71;
input ce71;
output reg[DataWidth-1:0] q71;
input[AddressWidth-1:0] address72;
input ce72;
output reg[DataWidth-1:0] q72;
input[AddressWidth-1:0] address73;
input ce73;
output reg[DataWidth-1:0] q73;
input[AddressWidth-1:0] address74;
input ce74;
output reg[DataWidth-1:0] q74;
input[AddressWidth-1:0] address75;
input ce75;
output reg[DataWidth-1:0] q75;
input[AddressWidth-1:0] address76;
input ce76;
output reg[DataWidth-1:0] q76;
input[AddressWidth-1:0] address77;
input ce77;
output reg[DataWidth-1:0] q77;
input[AddressWidth-1:0] address78;
input ce78;
output reg[DataWidth-1:0] q78;
input[AddressWidth-1:0] address79;
input ce79;
output reg[DataWidth-1:0] q79;
input[AddressWidth-1:0] address80;
input ce80;
output reg[DataWidth-1:0] q80;
input[AddressWidth-1:0] address81;
input ce81;
output reg[DataWidth-1:0] q81;
input[AddressWidth-1:0] address82;
input ce82;
output reg[DataWidth-1:0] q82;
input[AddressWidth-1:0] address83;
input ce83;
output reg[DataWidth-1:0] q83;
input[AddressWidth-1:0] address84;
input ce84;
output reg[DataWidth-1:0] q84;
input[AddressWidth-1:0] address85;
input ce85;
output reg[DataWidth-1:0] q85;
input[AddressWidth-1:0] address86;
input ce86;
output reg[DataWidth-1:0] q86;
input[AddressWidth-1:0] address87;
input ce87;
output reg[DataWidth-1:0] q87;
input[AddressWidth-1:0] address88;
input ce88;
output reg[DataWidth-1:0] q88;
input[AddressWidth-1:0] address89;
input ce89;
output reg[DataWidth-1:0] q89;
input[AddressWidth-1:0] address90;
input ce90;
output reg[DataWidth-1:0] q90;
input[AddressWidth-1:0] address91;
input ce91;
output reg[DataWidth-1:0] q91;
input[AddressWidth-1:0] address92;
input ce92;
output reg[DataWidth-1:0] q92;
input[AddressWidth-1:0] address93;
input ce93;
output reg[DataWidth-1:0] q93;
input[AddressWidth-1:0] address94;
input ce94;
output reg[DataWidth-1:0] q94;
input[AddressWidth-1:0] address95;
input ce95;
output reg[DataWidth-1:0] q95;
input[AddressWidth-1:0] address96;
input ce96;
output reg[DataWidth-1:0] q96;
input[AddressWidth-1:0] address97;
input ce97;
output reg[DataWidth-1:0] q97;
input[AddressWidth-1:0] address98;
input ce98;
output reg[DataWidth-1:0] q98;
input[AddressWidth-1:0] address99;
input ce99;
output reg[DataWidth-1:0] q99;
input[AddressWidth-1:0] address100;
input ce100;
output reg[DataWidth-1:0] q100;
input[AddressWidth-1:0] address101;
input ce101;
output reg[DataWidth-1:0] q101;
input[AddressWidth-1:0] address102;
input ce102;
output reg[DataWidth-1:0] q102;
input[AddressWidth-1:0] address103;
input ce103;
output reg[DataWidth-1:0] q103;
input[AddressWidth-1:0] address104;
input ce104;
output reg[DataWidth-1:0] q104;
input[AddressWidth-1:0] address105;
input ce105;
output reg[DataWidth-1:0] q105;
input[AddressWidth-1:0] address106;
input ce106;
output reg[DataWidth-1:0] q106;
input[AddressWidth-1:0] address107;
input ce107;
output reg[DataWidth-1:0] q107;
input[AddressWidth-1:0] address108;
input ce108;
output reg[DataWidth-1:0] q108;
input[AddressWidth-1:0] address109;
input ce109;
output reg[DataWidth-1:0] q109;
input[AddressWidth-1:0] address110;
input ce110;
output reg[DataWidth-1:0] q110;
input[AddressWidth-1:0] address111;
input ce111;
output reg[DataWidth-1:0] q111;
input[AddressWidth-1:0] address112;
input ce112;
output reg[DataWidth-1:0] q112;
input[AddressWidth-1:0] address113;
input ce113;
output reg[DataWidth-1:0] q113;
input[AddressWidth-1:0] address114;
input ce114;
output reg[DataWidth-1:0] q114;
input[AddressWidth-1:0] address115;
input ce115;
output reg[DataWidth-1:0] q115;
input[AddressWidth-1:0] address116;
input ce116;
output reg[DataWidth-1:0] q116;
input[AddressWidth-1:0] address117;
input ce117;
output reg[DataWidth-1:0] q117;
input[AddressWidth-1:0] address118;
input ce118;
output reg[DataWidth-1:0] q118;
input[AddressWidth-1:0] address119;
input ce119;
output reg[DataWidth-1:0] q119;
input[AddressWidth-1:0] address120;
input ce120;
output reg[DataWidth-1:0] q120;
input[AddressWidth-1:0] address121;
input ce121;
output reg[DataWidth-1:0] q121;
input[AddressWidth-1:0] address122;
input ce122;
output reg[DataWidth-1:0] q122;
input[AddressWidth-1:0] address123;
input ce123;
output reg[DataWidth-1:0] q123;
input[AddressWidth-1:0] address124;
input ce124;
output reg[DataWidth-1:0] q124;
input[AddressWidth-1:0] address125;
input ce125;
output reg[DataWidth-1:0] q125;
input[AddressWidth-1:0] address126;
input ce126;
output reg[DataWidth-1:0] q126;
input[AddressWidth-1:0] address127;
input ce127;
output reg[DataWidth-1:0] q127;
input[AddressWidth-1:0] address128;
input ce128;
output reg[DataWidth-1:0] q128;
input[AddressWidth-1:0] address129;
input ce129;
output reg[DataWidth-1:0] q129;
input[AddressWidth-1:0] address130;
input ce130;
output reg[DataWidth-1:0] q130;
input[AddressWidth-1:0] address131;
input ce131;
output reg[DataWidth-1:0] q131;
input[AddressWidth-1:0] address132;
input ce132;
output reg[DataWidth-1:0] q132;
input[AddressWidth-1:0] address133;
input ce133;
output reg[DataWidth-1:0] q133;
input[AddressWidth-1:0] address134;
input ce134;
output reg[DataWidth-1:0] q134;
input[AddressWidth-1:0] address135;
input ce135;
output reg[DataWidth-1:0] q135;
input[AddressWidth-1:0] address136;
input ce136;
output reg[DataWidth-1:0] q136;
input[AddressWidth-1:0] address137;
input ce137;
output reg[DataWidth-1:0] q137;
input[AddressWidth-1:0] address138;
input ce138;
output reg[DataWidth-1:0] q138;
input[AddressWidth-1:0] address139;
input ce139;
output reg[DataWidth-1:0] q139;
input[AddressWidth-1:0] address140;
input ce140;
output reg[DataWidth-1:0] q140;
input[AddressWidth-1:0] address141;
input ce141;
output reg[DataWidth-1:0] q141;
input[AddressWidth-1:0] address142;
input ce142;
output reg[DataWidth-1:0] q142;
input[AddressWidth-1:0] address143;
input ce143;
output reg[DataWidth-1:0] q143;
input reset;
input clk;

(* ram_style = "distributed" *)reg [DataWidth-1:0] ram0[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram1[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram2[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram3[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram4[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram5[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram6[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram7[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram8[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram9[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram10[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram11[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram12[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram13[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram14[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram15[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram16[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram17[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram18[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram19[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram20[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram21[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram22[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram23[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram24[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram25[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram26[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram27[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram28[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram29[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram30[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram31[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram32[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram33[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram34[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram35[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram36[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram37[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram38[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram39[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram40[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram41[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram42[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram43[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram44[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram45[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram46[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram47[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram48[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram49[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram50[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram51[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram52[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram53[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram54[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram55[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram56[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram57[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram58[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram59[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram60[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram61[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram62[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram63[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram64[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram65[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram66[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram67[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram68[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram69[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram70[0:AddressRange-1];
(* ram_style = "distributed" *)reg [DataWidth-1:0] ram71[0:AddressRange-1];

initial begin
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram0);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram1);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram2);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram3);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram4);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram5);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram6);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram7);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram8);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram9);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram10);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram11);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram12);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram13);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram14);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram15);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram16);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram17);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram18);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram19);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram20);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram21);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram22);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram23);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram24);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram25);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram26);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram27);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram28);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram29);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram30);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram31);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram32);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram33);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram34);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram35);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram36);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram37);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram38);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram39);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram40);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram41);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram42);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram43);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram44);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram45);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram46);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram47);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram48);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram49);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram50);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram51);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram52);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram53);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram54);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram55);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram56);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram57);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram58);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram59);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram60);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram61);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram62);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram63);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram64);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram65);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram66);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram67);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram68);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram69);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram70);
    $readmemh("./testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R.dat", ram71);
end



always @(posedge clk)  
begin 
    if (ce0) 
    begin
        q0 <= ram0[address0];
    end
end



always @(posedge clk)  
begin 
    if (ce1) 
    begin
        q1 <= ram0[address1];
    end
end



always @(posedge clk)  
begin 
    if (ce2) 
    begin
        q2 <= ram1[address2];
    end
end



always @(posedge clk)  
begin 
    if (ce3) 
    begin
        q3 <= ram1[address3];
    end
end



always @(posedge clk)  
begin 
    if (ce4) 
    begin
        q4 <= ram2[address4];
    end
end



always @(posedge clk)  
begin 
    if (ce5) 
    begin
        q5 <= ram2[address5];
    end
end



always @(posedge clk)  
begin 
    if (ce6) 
    begin
        q6 <= ram3[address6];
    end
end



always @(posedge clk)  
begin 
    if (ce7) 
    begin
        q7 <= ram3[address7];
    end
end



always @(posedge clk)  
begin 
    if (ce8) 
    begin
        q8 <= ram4[address8];
    end
end



always @(posedge clk)  
begin 
    if (ce9) 
    begin
        q9 <= ram4[address9];
    end
end



always @(posedge clk)  
begin 
    if (ce10) 
    begin
        q10 <= ram5[address10];
    end
end



always @(posedge clk)  
begin 
    if (ce11) 
    begin
        q11 <= ram5[address11];
    end
end



always @(posedge clk)  
begin 
    if (ce12) 
    begin
        q12 <= ram6[address12];
    end
end



always @(posedge clk)  
begin 
    if (ce13) 
    begin
        q13 <= ram6[address13];
    end
end



always @(posedge clk)  
begin 
    if (ce14) 
    begin
        q14 <= ram7[address14];
    end
end



always @(posedge clk)  
begin 
    if (ce15) 
    begin
        q15 <= ram7[address15];
    end
end



always @(posedge clk)  
begin 
    if (ce16) 
    begin
        q16 <= ram8[address16];
    end
end



always @(posedge clk)  
begin 
    if (ce17) 
    begin
        q17 <= ram8[address17];
    end
end



always @(posedge clk)  
begin 
    if (ce18) 
    begin
        q18 <= ram9[address18];
    end
end



always @(posedge clk)  
begin 
    if (ce19) 
    begin
        q19 <= ram9[address19];
    end
end



always @(posedge clk)  
begin 
    if (ce20) 
    begin
        q20 <= ram10[address20];
    end
end



always @(posedge clk)  
begin 
    if (ce21) 
    begin
        q21 <= ram10[address21];
    end
end



always @(posedge clk)  
begin 
    if (ce22) 
    begin
        q22 <= ram11[address22];
    end
end



always @(posedge clk)  
begin 
    if (ce23) 
    begin
        q23 <= ram11[address23];
    end
end



always @(posedge clk)  
begin 
    if (ce24) 
    begin
        q24 <= ram12[address24];
    end
end



always @(posedge clk)  
begin 
    if (ce25) 
    begin
        q25 <= ram12[address25];
    end
end



always @(posedge clk)  
begin 
    if (ce26) 
    begin
        q26 <= ram13[address26];
    end
end



always @(posedge clk)  
begin 
    if (ce27) 
    begin
        q27 <= ram13[address27];
    end
end



always @(posedge clk)  
begin 
    if (ce28) 
    begin
        q28 <= ram14[address28];
    end
end



always @(posedge clk)  
begin 
    if (ce29) 
    begin
        q29 <= ram14[address29];
    end
end



always @(posedge clk)  
begin 
    if (ce30) 
    begin
        q30 <= ram15[address30];
    end
end



always @(posedge clk)  
begin 
    if (ce31) 
    begin
        q31 <= ram15[address31];
    end
end



always @(posedge clk)  
begin 
    if (ce32) 
    begin
        q32 <= ram16[address32];
    end
end



always @(posedge clk)  
begin 
    if (ce33) 
    begin
        q33 <= ram16[address33];
    end
end



always @(posedge clk)  
begin 
    if (ce34) 
    begin
        q34 <= ram17[address34];
    end
end



always @(posedge clk)  
begin 
    if (ce35) 
    begin
        q35 <= ram17[address35];
    end
end



always @(posedge clk)  
begin 
    if (ce36) 
    begin
        q36 <= ram18[address36];
    end
end



always @(posedge clk)  
begin 
    if (ce37) 
    begin
        q37 <= ram18[address37];
    end
end



always @(posedge clk)  
begin 
    if (ce38) 
    begin
        q38 <= ram19[address38];
    end
end



always @(posedge clk)  
begin 
    if (ce39) 
    begin
        q39 <= ram19[address39];
    end
end



always @(posedge clk)  
begin 
    if (ce40) 
    begin
        q40 <= ram20[address40];
    end
end



always @(posedge clk)  
begin 
    if (ce41) 
    begin
        q41 <= ram20[address41];
    end
end



always @(posedge clk)  
begin 
    if (ce42) 
    begin
        q42 <= ram21[address42];
    end
end



always @(posedge clk)  
begin 
    if (ce43) 
    begin
        q43 <= ram21[address43];
    end
end



always @(posedge clk)  
begin 
    if (ce44) 
    begin
        q44 <= ram22[address44];
    end
end



always @(posedge clk)  
begin 
    if (ce45) 
    begin
        q45 <= ram22[address45];
    end
end



always @(posedge clk)  
begin 
    if (ce46) 
    begin
        q46 <= ram23[address46];
    end
end



always @(posedge clk)  
begin 
    if (ce47) 
    begin
        q47 <= ram23[address47];
    end
end



always @(posedge clk)  
begin 
    if (ce48) 
    begin
        q48 <= ram24[address48];
    end
end



always @(posedge clk)  
begin 
    if (ce49) 
    begin
        q49 <= ram24[address49];
    end
end



always @(posedge clk)  
begin 
    if (ce50) 
    begin
        q50 <= ram25[address50];
    end
end



always @(posedge clk)  
begin 
    if (ce51) 
    begin
        q51 <= ram25[address51];
    end
end



always @(posedge clk)  
begin 
    if (ce52) 
    begin
        q52 <= ram26[address52];
    end
end



always @(posedge clk)  
begin 
    if (ce53) 
    begin
        q53 <= ram26[address53];
    end
end



always @(posedge clk)  
begin 
    if (ce54) 
    begin
        q54 <= ram27[address54];
    end
end



always @(posedge clk)  
begin 
    if (ce55) 
    begin
        q55 <= ram27[address55];
    end
end



always @(posedge clk)  
begin 
    if (ce56) 
    begin
        q56 <= ram28[address56];
    end
end



always @(posedge clk)  
begin 
    if (ce57) 
    begin
        q57 <= ram28[address57];
    end
end



always @(posedge clk)  
begin 
    if (ce58) 
    begin
        q58 <= ram29[address58];
    end
end



always @(posedge clk)  
begin 
    if (ce59) 
    begin
        q59 <= ram29[address59];
    end
end



always @(posedge clk)  
begin 
    if (ce60) 
    begin
        q60 <= ram30[address60];
    end
end



always @(posedge clk)  
begin 
    if (ce61) 
    begin
        q61 <= ram30[address61];
    end
end



always @(posedge clk)  
begin 
    if (ce62) 
    begin
        q62 <= ram31[address62];
    end
end



always @(posedge clk)  
begin 
    if (ce63) 
    begin
        q63 <= ram31[address63];
    end
end



always @(posedge clk)  
begin 
    if (ce64) 
    begin
        q64 <= ram32[address64];
    end
end



always @(posedge clk)  
begin 
    if (ce65) 
    begin
        q65 <= ram32[address65];
    end
end



always @(posedge clk)  
begin 
    if (ce66) 
    begin
        q66 <= ram33[address66];
    end
end



always @(posedge clk)  
begin 
    if (ce67) 
    begin
        q67 <= ram33[address67];
    end
end



always @(posedge clk)  
begin 
    if (ce68) 
    begin
        q68 <= ram34[address68];
    end
end



always @(posedge clk)  
begin 
    if (ce69) 
    begin
        q69 <= ram34[address69];
    end
end



always @(posedge clk)  
begin 
    if (ce70) 
    begin
        q70 <= ram35[address70];
    end
end



always @(posedge clk)  
begin 
    if (ce71) 
    begin
        q71 <= ram35[address71];
    end
end



always @(posedge clk)  
begin 
    if (ce72) 
    begin
        q72 <= ram36[address72];
    end
end



always @(posedge clk)  
begin 
    if (ce73) 
    begin
        q73 <= ram36[address73];
    end
end



always @(posedge clk)  
begin 
    if (ce74) 
    begin
        q74 <= ram37[address74];
    end
end



always @(posedge clk)  
begin 
    if (ce75) 
    begin
        q75 <= ram37[address75];
    end
end



always @(posedge clk)  
begin 
    if (ce76) 
    begin
        q76 <= ram38[address76];
    end
end



always @(posedge clk)  
begin 
    if (ce77) 
    begin
        q77 <= ram38[address77];
    end
end



always @(posedge clk)  
begin 
    if (ce78) 
    begin
        q78 <= ram39[address78];
    end
end



always @(posedge clk)  
begin 
    if (ce79) 
    begin
        q79 <= ram39[address79];
    end
end



always @(posedge clk)  
begin 
    if (ce80) 
    begin
        q80 <= ram40[address80];
    end
end



always @(posedge clk)  
begin 
    if (ce81) 
    begin
        q81 <= ram40[address81];
    end
end



always @(posedge clk)  
begin 
    if (ce82) 
    begin
        q82 <= ram41[address82];
    end
end



always @(posedge clk)  
begin 
    if (ce83) 
    begin
        q83 <= ram41[address83];
    end
end



always @(posedge clk)  
begin 
    if (ce84) 
    begin
        q84 <= ram42[address84];
    end
end



always @(posedge clk)  
begin 
    if (ce85) 
    begin
        q85 <= ram42[address85];
    end
end



always @(posedge clk)  
begin 
    if (ce86) 
    begin
        q86 <= ram43[address86];
    end
end



always @(posedge clk)  
begin 
    if (ce87) 
    begin
        q87 <= ram43[address87];
    end
end



always @(posedge clk)  
begin 
    if (ce88) 
    begin
        q88 <= ram44[address88];
    end
end



always @(posedge clk)  
begin 
    if (ce89) 
    begin
        q89 <= ram44[address89];
    end
end



always @(posedge clk)  
begin 
    if (ce90) 
    begin
        q90 <= ram45[address90];
    end
end



always @(posedge clk)  
begin 
    if (ce91) 
    begin
        q91 <= ram45[address91];
    end
end



always @(posedge clk)  
begin 
    if (ce92) 
    begin
        q92 <= ram46[address92];
    end
end



always @(posedge clk)  
begin 
    if (ce93) 
    begin
        q93 <= ram46[address93];
    end
end



always @(posedge clk)  
begin 
    if (ce94) 
    begin
        q94 <= ram47[address94];
    end
end



always @(posedge clk)  
begin 
    if (ce95) 
    begin
        q95 <= ram47[address95];
    end
end



always @(posedge clk)  
begin 
    if (ce96) 
    begin
        q96 <= ram48[address96];
    end
end



always @(posedge clk)  
begin 
    if (ce97) 
    begin
        q97 <= ram48[address97];
    end
end



always @(posedge clk)  
begin 
    if (ce98) 
    begin
        q98 <= ram49[address98];
    end
end



always @(posedge clk)  
begin 
    if (ce99) 
    begin
        q99 <= ram49[address99];
    end
end



always @(posedge clk)  
begin 
    if (ce100) 
    begin
        q100 <= ram50[address100];
    end
end



always @(posedge clk)  
begin 
    if (ce101) 
    begin
        q101 <= ram50[address101];
    end
end



always @(posedge clk)  
begin 
    if (ce102) 
    begin
        q102 <= ram51[address102];
    end
end



always @(posedge clk)  
begin 
    if (ce103) 
    begin
        q103 <= ram51[address103];
    end
end



always @(posedge clk)  
begin 
    if (ce104) 
    begin
        q104 <= ram52[address104];
    end
end



always @(posedge clk)  
begin 
    if (ce105) 
    begin
        q105 <= ram52[address105];
    end
end



always @(posedge clk)  
begin 
    if (ce106) 
    begin
        q106 <= ram53[address106];
    end
end



always @(posedge clk)  
begin 
    if (ce107) 
    begin
        q107 <= ram53[address107];
    end
end



always @(posedge clk)  
begin 
    if (ce108) 
    begin
        q108 <= ram54[address108];
    end
end



always @(posedge clk)  
begin 
    if (ce109) 
    begin
        q109 <= ram54[address109];
    end
end



always @(posedge clk)  
begin 
    if (ce110) 
    begin
        q110 <= ram55[address110];
    end
end



always @(posedge clk)  
begin 
    if (ce111) 
    begin
        q111 <= ram55[address111];
    end
end



always @(posedge clk)  
begin 
    if (ce112) 
    begin
        q112 <= ram56[address112];
    end
end



always @(posedge clk)  
begin 
    if (ce113) 
    begin
        q113 <= ram56[address113];
    end
end



always @(posedge clk)  
begin 
    if (ce114) 
    begin
        q114 <= ram57[address114];
    end
end



always @(posedge clk)  
begin 
    if (ce115) 
    begin
        q115 <= ram57[address115];
    end
end



always @(posedge clk)  
begin 
    if (ce116) 
    begin
        q116 <= ram58[address116];
    end
end



always @(posedge clk)  
begin 
    if (ce117) 
    begin
        q117 <= ram58[address117];
    end
end



always @(posedge clk)  
begin 
    if (ce118) 
    begin
        q118 <= ram59[address118];
    end
end



always @(posedge clk)  
begin 
    if (ce119) 
    begin
        q119 <= ram59[address119];
    end
end



always @(posedge clk)  
begin 
    if (ce120) 
    begin
        q120 <= ram60[address120];
    end
end



always @(posedge clk)  
begin 
    if (ce121) 
    begin
        q121 <= ram60[address121];
    end
end



always @(posedge clk)  
begin 
    if (ce122) 
    begin
        q122 <= ram61[address122];
    end
end



always @(posedge clk)  
begin 
    if (ce123) 
    begin
        q123 <= ram61[address123];
    end
end



always @(posedge clk)  
begin 
    if (ce124) 
    begin
        q124 <= ram62[address124];
    end
end



always @(posedge clk)  
begin 
    if (ce125) 
    begin
        q125 <= ram62[address125];
    end
end



always @(posedge clk)  
begin 
    if (ce126) 
    begin
        q126 <= ram63[address126];
    end
end



always @(posedge clk)  
begin 
    if (ce127) 
    begin
        q127 <= ram63[address127];
    end
end



always @(posedge clk)  
begin 
    if (ce128) 
    begin
        q128 <= ram64[address128];
    end
end



always @(posedge clk)  
begin 
    if (ce129) 
    begin
        q129 <= ram64[address129];
    end
end



always @(posedge clk)  
begin 
    if (ce130) 
    begin
        q130 <= ram65[address130];
    end
end



always @(posedge clk)  
begin 
    if (ce131) 
    begin
        q131 <= ram65[address131];
    end
end



always @(posedge clk)  
begin 
    if (ce132) 
    begin
        q132 <= ram66[address132];
    end
end



always @(posedge clk)  
begin 
    if (ce133) 
    begin
        q133 <= ram66[address133];
    end
end



always @(posedge clk)  
begin 
    if (ce134) 
    begin
        q134 <= ram67[address134];
    end
end



always @(posedge clk)  
begin 
    if (ce135) 
    begin
        q135 <= ram67[address135];
    end
end



always @(posedge clk)  
begin 
    if (ce136) 
    begin
        q136 <= ram68[address136];
    end
end



always @(posedge clk)  
begin 
    if (ce137) 
    begin
        q137 <= ram68[address137];
    end
end



always @(posedge clk)  
begin 
    if (ce138) 
    begin
        q138 <= ram69[address138];
    end
end



always @(posedge clk)  
begin 
    if (ce139) 
    begin
        q139 <= ram69[address139];
    end
end



always @(posedge clk)  
begin 
    if (ce140) 
    begin
        q140 <= ram70[address140];
    end
end



always @(posedge clk)  
begin 
    if (ce141) 
    begin
        q141 <= ram70[address141];
    end
end



always @(posedge clk)  
begin 
    if (ce142) 
    begin
        q142 <= ram71[address142];
    end
end



always @(posedge clk)  
begin 
    if (ce143) 
    begin
        q143 <= ram71[address143];
    end
end



endmodule

