// Copyright (C) 2022, Advanced Micro Devices, Inc. All rights reserved.
// SPDX-License-Identifier: MIT
/*                                                                         
*                                                                          
* you may not use this file except in compliance with the License.         
*                                                                          
*                                                                          
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
CaihNQWwu+qKJWjcmdIgzgKIXQ8l3vMImmWHnChjYqoa51yMcErBScyiE64YZSDih9WCUqsVfjEZ
HfdPZ9ljuyASaDAJWOBnJBbhrePBDPO5jKkFmPbv80QoBXSWaNMFc5sW0Ulg3lCiE5qq9SVr7IMd
vkFVewJkI9IJKPXIqEiYLMio527A7EkzJrjUXC11BQnTYghbA5n7/6q2WIDOwjQ+BdLZXxGdIUKi
ihIieqBZEgdd6vwETSGv3sSorIwnUPSueC94L800xEEoFQmghwgPGvLA3IEIqt1YNZfrY4rcuvTH
rxE5ve/ar6tMYP0QdSitAf/UOVre3EWtsP+Jcw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="IxINXwVvXQ/n7KwTaYrPoEaEACBK27oPy3cRIdl/LOI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1219024)
`pragma protect data_block
EiGu1ShDtOnFp1/lwt6VhVnr89cfK8CKMJ2UPGIzilxEuTwiEDclURCinPuSr4AeMArg/BvgN7//
oHUMQ6ItLPVJK+DBXuSqEx/nVO87wjtL8hTSpU3NGRWQG7rUNDwFHYCD4mJyL+w4e3KqStsscXGU
GcxhG47ZhKGm818YviW8QCLcWALdMz1Qya9xTqt3v1yNs4V7aImopMHL7GkQ0MrVGMz9AItNoz8l
OSy/o18gequ81DqC2cT7XAMMWG7nMKBZDEDxTBcEV9gYstVm8+cpjyfQFJUdeZKNIZkJBxYzVM7V
z9u/Ii3xhjODAmwP9IAMbIg9Ex7w8Bhh3SoQ1YG4MvB/cUR2nWRMNnWcfe+rlJe+VnIJPb9Q/jNQ
10naNt8wzmWMNXwEbbR1TYx301r4/vekmfgR9kxpH6A9f8D0oL08SnLsBdVvF9GeJfCcR3ESqNjq
Db0KsCG05ak5ge95G4xumYzp1sbe0RfVBo8VnXQvRhlt1CsL54B9fl0E8RrSwsbyfbSzkOfks2dr
8qI+GzyjPSrPbLsi+FqH37ohPndyb92D8mC4r5d6jK/pv3TCC45mOVdy2d3Lryb5qOOfpABhblJS
QihuSXq+YLWi1u3Na/KsdJp5sGOzkPMyBQ3F/S4U6M8zeS2lMtvY3WArWRFjQy85BFPFt4Qj0QbS
EXG21MXDes1BtODd8kTU0Y4tgVbix4N4uqD8dZcR3xKXf9aoul3QxdtlNkNuPMfLDVwncK20V731
pmMmSYy7Py5mHVlYbpcjuuqNv9sOaCxWWLWubqiadKgzsXqVd5Td4ZMdGdSXfA81rVclkxWn7TTb
Or+Hnx2VuMzLqrlztIH+vaqEG34j3jgr2Kn2fifj1pKDpu/2UIwsDSjhXh3HR3L6HuKlo/PydtsM
5Y2rhVAtBroT+RGvCFQW4N1zdegpVn+3PaNLOFZomWUh3rx/n9/mPVSna7a5cKTzN2Z4Ab0VuI4s
O0BziEMKONCE62ZCDhO0Mh5aFnm8it0nS66SKNOxM2mSygf+7SPtURM3HN3oNP677X5Brnlb4BWt
QpMLymT7zAlM+Dq20nGeOPFbMD8hxjC8T76hKvBUh0UCP8FBqJhuiY+d66gabbI/XB8GYOzS+Cuq
s2cxvJ8AgQMEb2z0LT9fDkThLdBHUyHdZ1fu0lkMJ0g/LPaMz3yRv4IeGY+06s4+095UNv5Q3i7F
8g60pdsdhD9YKbp9Pf5Jve+6Tla3ea1XdqC2EIKfxeILsf0arrd87jYzd5/ENrJpR+aL9w/mkcLU
OS29cHWVwvOCRV7r/Zgs/q3QhL9OJfwvX0phyU0rjwkCXdIC5o6Nsz9pFjoI2nf4D1wGAqEBRxJq
0vpJ0UY6pHKbX+4E9QEQZ3AOkMTbhgmaQvimGLHArAtqh0osCu2wY2ZSQ+OoNDNSKgOq1/+S/AIs
R4Cv/iYXtD4yEXat0LZNBzT6Abu3+2BqkG+CCYYnKex682jW8pw8Uom+z1/f5w1mGMnlGiHR0fJ1
nzu43q2oyMqkFzMXOmykBJDhvq+RopjbZ6bdB3zv4WTzA6Hc1fofSDHY97KA28XEXrLqYXt9A5HV
Wfl5gBm2+lMAI5zuM65T5vFeytKpQRivh8cNRrmwPBr+51uTtpLkGpHM9zR/U4KdrjPTxSd+HhCB
zH+emAlh3yfZQbw1j0EFubwfVERJZbrQb3CybVqYRIx8A+pyIFVqRUixnskds4dngG32wgybJqwr
M52yrNfNYrW8aqxwciQbifO5MN8btFvmia2027yZ7TWezBRJ+7C062NVpwWSe9+1eSERp0BrXf5u
tSIkz9/8lVT5Q8Xea6u6/qtC/G9zf9ifPL260uiqSRQ/5awMUqMaHumawqCXZ0WZGkW2G248h8aY
OQFlSaArxpntyKZ3qidx/lzL46HkdZVvFCN9aXA6oBVxnO1v5Oyk9MMg+n5oujrQZ8yT0j6DgZYB
QkEjpzyWCYyVVmFtTjGw2WEjoCEK8O/Pb1PvIfb1OnnUxv+yiYKkoLnTphaVctSQW1mHUxrT1IN9
2hW3sxXTvamN0WC99TefdEN/pxHg+9VnO903ZdBdlmQWEEq+pEt5SpuorxnqY3HUBwOOiRYYarZH
f4HN+LBwg3aTZTA90nDXkWlR4P9PSw7dSE96A8u2u37jah1Qb1VlVOlMp6Iz/oO+f6VZRI1oNmGO
O3Tl5X5OjHZHybLavFb3BgBoi2qEYxu3ekqZIx7lZCNMxcex5AX5P0kkj7y8IQNx8a93TigAGCzi
XgTgtpcv697h91fClU8BXzuhR+0xP2Z3uhCcTaqE+5CDCkp5vdKsMp+wSBedsnTFLOf7yc7jC36E
GAasybLEXifKSkaskiMI6llvnfuvBP9jVtOHTtzpcseodZ500bA5pDagIlVORfY3YOCzTZ0Ynnx4
JVUMhKjf7Q39ss47QVOKITnYO1/VPQHFVlDvcCAJNZcSy/DBwFa9YtPp1riorkMcDx0iL5wY/VM7
Dw2WhoUyMJnE/ZLXezSvDPG61zyo23M5/CMGWx6Rgi6lTH9ufX6li0mil/mBDUgkL/Uew4iYLuXO
RKYoRTpBKbhXe7bhf/tKNzTeaePYUStaTvfiwz12OKBu1NhhFHWRVn3zkct895xZmqiPTtfiPqsK
aLw1vH9SvMGW7W2qkW0zxZQX2gQBf484ivxKxgb+VyixwwSpvHMgjf8SDBckomOwDdJd7uSeJZnM
fDrTR8Ssqrq2pkOZ/s3e+DVsTcuKiFhHO/JrEzIXbmENo0URSfawbMrl10KOYhxV9xlMNndqJOqu
ZflcS9GdZZCiZh4BvZeb7vQQx1HzzJT6ZJJDIwfLGx80o6iV2LSdw2Le6Obh2Qtyi8ztjQOUMJCb
AG7bsOY0jOO6hzhbtSPS6lBVois9wa2VKuYj4MNqii5Rc+Ntdj7snlczas3hPB/HMTg4h2A9a5nd
N+d83GwKOZQLPnIcQk9+lBBZaCEtiAnH7hXZ4s3txZZLIMn6SZ2xPAoRNXjN4XgKglipDwB7gkZH
4mfOeet2iR+KObQU2CxD2Fu3KyKwc3hhmhPO/hEoYjRahtrKbGT3TS1xdrqbqn1AIby7qayiG0Bb
xk+93VBKug/4LFBuIBPRhXlv8c7wXje0FqbgeNI7doLDXC5OZZdaj7YaoL7gvMoX2pAw2DxrRhMI
fReH+H0nvkBgC6VDX7aceFTyi8FDuYaB00RxOg8vsbZWnZ8i41h6GbxuYiK8TxvIoGrNQZwTi1YC
K1S8GJ1InoZM7HZOH/hfAwRvDVjgWjKHqgBt7f56q1rvAHjDQl81xTf7nyKk4rAt8ND+1Yun+Q0e
twXqB3ijZ/EP9NTxyUFkfiHl84liZH+/ndCOTY0WL+cT+CcEmahqe7nB80k9VM5GFv3UdoX9wuBY
x/QiRMXJ6F6NmKNWzeYOEfDEVYQzFXFepGQoLczlF+njjCDK9OmnK3/O0TglMACRC1pJsbspBO3F
25IH9ZNSu3qmEPharTTHuybubgxDWkoXxvpaiBWHZUNV6GzPTznQwyVcirxgj8TuDcPzsMsXlo3i
hvfck7FIRyUWUoMDbfniWU/LzjQo8ZVkUZQva7kJfkwx9Q6YPT6NsDhq2FxNMA6Vc4mNpuc8qVwQ
/RTeTxtdzufjAXchZc8f/h7lLEWrqzYWzv9E1EUeXe6BtRndBFwpN5gm05zzrmi7YGrWQfFHnBEo
O7jFufxw+lIXD0tjOMDWBP7+6B0Y8viUn46cKd6MSU5GMwGV358HZi+zRBHfef0kJcxUcCF4kU0o
EZQ9mecIbT7/9ch0mwSrLdb4rfn1I+ixbnbbS0rbSf7dc7ykWusT66+sng8Q9/rbwV+wBaMCilet
iwP30010iTqkcCW2SFILwJrUtFCVhFD0/Y9wd5sxf+h9uPsuNM+C1TryBapPz41r1kkC9RfTvYxa
Nmq+pnesaZ8RPvBgtk4Ha9qjZ/0SoBBarBdRcJ126R2PFG6P6NGuKJVgbAM7+hCLWJ+0dZCanM2v
f83C70svi4L23kzzOISZVq9AV6/eIIYoCWljGtjRWnHu45a511gBMF314WWxI9qBxViTnbakUrzM
wq5lHP1vwGLnrCM/Yu6bGGOvXIPS1ZJXAgl20AWrLBdUWIaFPPVWdV4wZzGeyz1JNfMdV+xMIkAZ
JoCRq97MVdh58zVS2ec1Lx5hCI68Ov/NO/CJvYWhgb32crqzvgy+clwPPInQlf9Y1i9VZSbmGJZ7
FrKphIu+938ZYYa1RtTwlayKY8GjpmKIZ/IiPp2e9VQ6DdClJ6xPxTK4p6kCV+sBkChn3bAea5S2
4TJe36VxcrZccDafncolVpwTndBTFpaI1echjK3xPS+FAelSJEN7pZ89/e9fdpuUMZFdKkY+/0yj
ffM+Oo2wcUBhR9GAPaPcstkskpueXL+Pxu99AQhUIDTGQQU6Zk1PDqs/2f0wyGzv2o5s1qt3ipRD
6yTPM/+6bPx7h5xKBNgSgbJciUaZl0GZwIkDf/dKowE8u+FQwSM7W9nLFUnKYOroSp2aUJFycT/B
n4Hj0Nu8h3qc6LTg4m5hrsiqS+92EpW/h2dCPHdQvtyvGadwty6/YXwpuIJPJfuhS/8hV2WpWlBU
M82EQYARlEaScgBmWJcxMG6sIxT6lMR5gK4XRIneQAW8fzJBmtR9Y43L2kQBKKc9/D4eUZpymshC
lHZAhkRWaLsLjLqAr9ifUkjt2UyOnTmv75jKBVYZbdtRcoCD2hl7j/yqqbK2Xte9ebCgh4rAFLM2
xeRs9kp1FxPEtbR9UDN5JV2+erLk0oyEzdbAhdShHOhQPSd8Bc5a3wGhHql0yqCYISRiIfHmQExT
zFtmiEQtiNB0EgMFxiTWDB+6QX+I9BMKl4Uzj3lQJ1nbDJd1i7SiMeDNNOC1Nwg1hWxlbU2la7dO
eLEEj/sM+IvLr05bTkIFXJpI7oXiCe5dgRIWIeBzYc02A5laldwXzc6uo2oVGtnwsrUDRRF/Jd69
53osNtgoZ30I2IooHIHjPPaz9hpp3+YsEeTfv+CeTMSXHClrYutby4OXGfvVDFRPcoNSSEj7DQWf
70jZVQgv9LMcbkj0/7LXj5VRb4ThSafOzYCjtvdHDenVBrShrgc4vSedO2q7RVZN/XOnbfgablLI
+CXW9gNsytMFGPYvT1hEWVl7xwRzgyRHVZx1iVZKX/snbYCNyfBqQofvE9eCTkVdYnqeAEdJwb0u
YndGpuXCYZNiu7AvEONbX3qj50ibx+WuuY6wPR+VmW0OamYeAPu2RQWiUpT21o5zRiOFD1u66WqC
oWuLxOX+r6rPJAhr6IourobnCOTFyHTb0Qlu8dMTi23gku46xtcM36b6FpL2JQ90OH2OMoFB8efm
dNIkDTBW92vFKt9ldEf4I36TAc4/+iHZed2KRq6s1UpUA5Jxa8WbVREc+UaQWdnC4r3Y+bktHRVQ
vxtMo6xuSpY2YDlHeKTWZTenZS75EYxmJvVRvJzLZuFQCaMgCy+fVgZ45l+1k4gvbdrx2MQdR6Gt
IsS4tKdn6pipKDsyXOTitmlJdp8dMiezFAzxHfRm6J2DDWWwtKte5xo/rpPa1ztdcZ9XxmKaBRnH
dpC7I7TlmPmWB7grLUdQtw4P+rqDYJzlHzi7fnBu2Ebro9jhC40nxxg23Cc42TikSvJAe9Q7Evx8
ym5/PiOyXFUrl1csDM9jqPRZu0CU9tn0wkxOXtlk2D+zWaFpYSqUWqpVRlKXJvDwk9iqEfiLsHRl
OLArG7R1LcOK5ia7JcPU+RwtwyJJ61WMIOZxME+TYEWGefRJttbBzodRwGFceGUpcgbbn5HdGtN5
KET+h+2VJX9mC+8Zc7pQ3fFgtccjvL6rOS5Tix9/Dru4QdkaK4X0klE/9gedIyBEi4TwTc5UTEU2
P672O62IMjrdl+GX3qEXo59iwzbxd2+lqTZVKrPNDaOJp2r66GLp7ZM7aRqGiDDlRCXs5E7gOeqT
0GgGj/VPK4nZFyjauozniD0PFkQcpvAQBL3dPc8govc+k49N6bueVIqGGR2Z2cEuM0mYb5gM0bmN
qETt+adqHrmGS5nmjJRE8K0sUMQ/zxs+AVcKNCw/tCKicpJRBBRq8WVMSJNNoIpy/c2hLsaEqcID
aJ6ViOqgSV4L7Y2N25E6BxqbP45gJJ+X8fMirmSPBySeHwokkiUs++foOY54LyXQsJ9LZzB/+Y6P
4Sy6R8/S1K6tbJl6GxBN0TTmFQhUxyOJOC0m8VqU2g1Y6TP4G8MsQuuT7FmqJ5nn0I7vIAGfO6rO
BFJJ+Y3aCRNEsXXNUNhb4RNrVMBTKGMgCo1D4p1ZkPPRe0+EWBnyzYv/8vMz41gaXNZmMu4vckm2
OUVCq1hzzIWUwTpDJ3+kP64sXRXxi4OD+W2ltPSEcuoKbaB18lzLv45jfTFI4dcYgjCD7obvmH+J
aMN+f7tdnEs4KqeCJd6mOH9g0va61iXnU0n96qcf6Nzlaw6NOOyRO+CLbd1PtpzThSascJkGkvv7
ydl0VFhO8NJGtrAP7V3TlFdKyvIcR2oaCQ6g7B0Y171FqXio/9BTXwSrJAPwiGm5F4IvFejVz2SM
FWPYKktlN3JfhPH6jZ8hYafTyKlgm1aPFupxd9LjhdCRL/iy9D3ur9zazVB02Qcq2l4kjHbkZKuZ
VpcsvAeujazHQPIhtqfY3x2sqwqma3sc3I+ReZgCE/whvalMk8j7YfV8shR+EKk5rpvxfkNIk/Hi
WeCWWgJJVW5pyuDRTHsRSqA6jlGH8jhdiqDW/vHRSI0eJDr9YlB2RN4mrXjE3aYqiRJg/g9JznB3
SSAeWqw7bJoENzu4c3RSCRoKi3AZKylqQ8tArk64RN00mLB9YuXEL+yyRSdoFB28MQgSvUHZ9i+P
Vyl7Ytr7W+5tFrBm4GgkpZk2HX8QepnTckLQi4vUTbWui8w5LMDSu/KcZJAdUWHxYZrl5zfyB2O6
HpEmg/JcsfS3dzpGxGf1MNMiLVdGq0wMiSVZPMf11ZcF6ZegUCjFCIT0b1MJs22FFz2Q9tCBv9gg
Ur+tQyhdHqH709ZmBskiZpReLrDU0F4uKwd7C8UdmMv0nJnzlm5Rd/2LxdUEg+YyOBhh55EKa70A
+ZJU9hqRg4QYoshQnMQtttbGF6Bw6pr7IlyzTwW9BbVjBDe00NVnm0htGQ2V6d4e91guis2Lh2g0
k8X+DmKE2m1jKjlhpBmh7wZgiQGvepvR4qoIDTErya0z3tTFN6gTtOtbZMYIsmgfmEmmjvzENwj2
nDQF3XVUA4gHuk+jxphb9XYrhX/v34k70srYmURRCl3o7Ww0/M0OW45qdcNYPQL/kvykDzu9yFbJ
5m3ilvfgItgVZ9v3ENTLXv1WG3X0Ldkve+j8+cuTkRg/rZ9YiZnREHGvNuB2iy4qetndWUvpmB5R
J0iTGnDZiE3jHsvyzAr1/eeUpGuq6sXTCF6j7wrgI/+JrRdloxHELKzHEvnfvZZjnIR8sFPDqJSN
uu1FRyqCJIPW42ca4g1KK/NnFtodUnn4FFOjBYkCR8sF7I/OutS0Jg9imF3+TkK7z0NPd1tcxu6f
OHtUXqRj4wOSIIW/9GOPdPInLHikdszHsquk0pfH8WzdY1aNf27/AjYj/07eO9Ev41zNr8TY+Mrw
51ENwvwRso+tHscdqQT1hYROD+xS21a9Ikv6q7h9c7lUkZINXkm+WfTsQovz/PwiCu9LoSQb+sLw
dyJc38HEWjltcBZCmM2+hXxLV4HyigysULgnectDfqmrpLE5CzrG+oUjbTtztKy2Y4ZMdsygB5B+
GM6Tj/mXfQdAq8maoj9yjEN9AuJ3qFVeDCuXPWlJmTXcdcrm49VL3Z9z0+hqOMlFfhRXvYAvRe4a
wb+IjE95B2XIPFPTdZkahxxx96i7ZhbGj4y7bAoOeqvZc9JVasNoLbruw77x0bONdZRcsdh6RKOR
kX7AuQp4OUm2BMGT4ULAFidBUltZT5FEYuxE4dsiRyEGZvOYjWAfIF2MIB7q+8IXTacYzOVC6lHh
N9mTGL6XmnvIjXnW78+IifPCLkRju27RfgMDrbY7+FmiSFuJ6dy38W7QxxVT7nXOa0D10hyc2IXD
wzOXUxfYN4hgX9rEHyzoiZCU4eLUfqA5Bh1no95uIa2qzGEyRj+ISKbiDZitEIV4UcLBJH//j2Ea
I/uA8l4QeNqinZ9yKMR6pTahXaktgbkQUrTnSnSuT74BlzjARAbZFyuV2Y6CSAf9TuS+jEjxDcZb
fP/UbBIMEsdkfgMFD7PfqyznjW2P5liT0Ly4WA/u73fQCsByerrSZ3fOUSkwyXo8/VC0drCOHf9l
aajeBuRvl2/n02boWEBb+6wJ3ZksYmHb+JbEJfccsWhOvQh6cpH+omMmARXPtamOKsBJag2U+7b8
bzpfLw+P7m8kMa1Te9fJqFVamZgH9kzLLTxsgXIJct9eWYiyubBX51R0iRPSaBGKvgIbshGChrua
0PgA19q16moDPttD2uhcPamXMIJl2aggPiuSy/yHG+GQbMWT0APEpJyR5qGz0bQdfT7bROWbJyVk
XBbn1oWNTLEIowHKybtsIy/AjvOi3qB3tRQWA/hzuKutEhk+TCpLv5h6FzRtAy2mn4vIDHeYJ1Cg
E50sQIuD/+0jSD3KmmnwaCdAYxdjz5xVXqDqQIygke0hg+kHRMT/FAj78zGXYogusieElcbFizYQ
X6EFv+26XsH4ZZNWrhbybi+KfOivJLHp5mUn3Pw7AuALYWVGl6ziII47LPnSYtGeLgZbzGF34jB6
qspVKD9Y1kpAhmNJ9Re4d5lmzi4OP52/Y8S3iRBMHpo9wRhKOtHQAVBni0yktpEKM8gql0bEPtDO
coOeQtzsjhPw0gq9w/cFPWlf0juJfmokxbZHFAq7o6+WNpWJVYLv9KLWIvhYvjIQ5Zn0Ix/xRTer
XAqfK4zLZqGGyhTZvs0DEFh/uC2+ITl6ZFqHSvvvqZqo8BLBYZbdPuPibePi0rfXh9pyk7J0xSLl
3d0t+pQQDk9MwW/auRbHyFPYDUv4321nv6QXf6YkqBD3X0va1fSUg532R4aHMKHowSPreeyKCyK0
BpIGjIIkX0mJik9mpzA9DQN+Nfrh7FknjXVyWUI/sqd97BO6jBbzEMo6kN3LBqztv4wfjtYxuGvi
sBkJgLOaGMNDMGYDO1lIooEVQK4F+sEc9+QNG5x33noZGsH5Qw7DLikKGtLzSjyN/lyTVBN/I3MF
//LemSUShf2b9KkkDebWInsyIIO8jr4dAFamp3jk5OVCWDnYLbGyVCqVIi2BBEMKZY5ygEa8MtkQ
eu2BZcKqI757tsMKREs7EP7zkboTWWZjUVNDK3HU8UvrnkcV8ituzV8/uIvDRp1l2RgoLN3Y/vYr
YAyw1rmOvcwK9SBFw73FS2h3ypxdO/AQA2fAKzS76fjNpgab2vxHcbQoSF9FFSsorHh17I/WT/GV
+ldmHsTdjYwvxWydFPupXdnEdN+c1ZYPmWTP2V6KwogZuufS6+n3QzyNtsBh1TRj56QwaIMvF0Mc
QqwtLBTfdi5+hBq5e+NiA5ug4mGi6ERl0C8tHzxV2vsm8YE0Rn6kNBXZlxXb5cvqqn5BtfCxpxST
NUG/x4xMoNuY2+pwPX4nMqtQ9gaprQAz+mDvf4XiQTONX6WAhR2fGgteJB4M6KD2dfJcmgjlzMT7
3ew+4jS4ssH6wYKbbMBreBj324XapcRvIANoOdh8bN76y9NNKFhwayEEOChab52Mv2eG5nDQSZK1
moXGeXcXGVzQA8Q/KCX9eX/rIQcdTsXjfoGImnCAxOmc4SMGaaI9RhOe0OD8dWGTIcTOOsPHKWdy
eLanLCizrS+szWrk8Set7z5I0nm7BsGVeZY6KUvDv1gDYdHmQuCDGZtKdLefzOFsNJ1y76pNvNFa
cxelEeUVqIEPibT16z3aSYL7xw9j4qJ+1bManqAycxfFntAHn0nCSHUcztfgk2FeIVbEGNqf1Du0
82hrVXhb4f/tFnUmhjN61NN56WxMvRJXaip2DamTVnGzq7rdsueRpU8q6U8YVBts3axZfBGkr5/S
byCdeR+ZJ1JcwGl0/WbRVp+2xj9PVZlp/EvQpVvcy7+Bg32WyZ1xnvqGM/SU/9C9IZlTzAu/deRu
yskHNPh0AuM+plXq2wz3TKR5o6MXnR9SmmrsUT+w51fXUkM5bqmJw/8E5VYP4IQ8TTrJR2//0nTT
KuDMJAaLh/msl3ztXoOhCi9zG0jzTSHaVNbnT2IsVbiiKPP/AOxNliIBVAMDfdTxJDyXFEEFfdLu
5Xo3DEJgGKWPjoX5mYEvbXqrwRZWYDEJXdj5ibJ2nkUP6lkIBAzXEXLB3ZjW/KVgkEbpfvHeJEmG
vV9buzViIitGg3ImaU6+a9Vt92utovO0vMLykNDltEmVLPSuMWOlrnBOU2l18AKOFCHocfqGTq2c
sgySHS2y8XasBqcup83HCXZb4Ucd0ssxYFTguTj5ZXRDuxWOv8Jy6KuC2CJADuti+X8oGIpKUOGK
a/FFGa5HP3u85cdd56zfHxpBLxH7VXKh4rhlhMaUrrFteIKIJOnz3ycQjUZ0lcDqKO8fzUKeTha2
cm02kCnKJkCfEumJMeF0QUCdeMRNHjdjKEQjJ5Ty7Qe89WPordwJsAaXw28mM+74k5y8pJhEfyU5
5cP/bd4TYgLERy4HxhMxPj/6gGZKdZlbkjc8kTjRZroFIz5aQ82dvcLijWuzE0tdcujm8Gtr/hV7
fS01QleD9VOefHrO/CgEsziHbu1rxz1OJKQnJpMRAFXOGm3B8KuPQWCbtcySB7mS+WZKdcMtesig
VGINBFg8AG2Lm/EyrmmfH7h1q0560l4XxhNxbHxKB9XsfmOJBlKG6YiWqS8jWDG3IlMiwLoHIDjr
05Alqq2/u9YP34Etmr4wzyAAkVQ8Rtv5+I6zpx5gK7v7ZB+eNRmHwap1P3IdzSv6+6HghQFazYMT
G/uBwkTFrpWYx8qzzCtNatlDp1FwBZX+gfvy8pjifgMX/Eu0MNIbdOH34pxAQ2y5B90lzc8bqO5A
FY0uMpqShYOBkKO77pRuNnmiN/iWAUUitP638xdzhVphmZrdlK0yNdaOk1LP4pB+QVsZhz+uglsB
HXQWXHlLIpbWFFPxivUHqyExFEINpVUJMgWLWOdVSep/eoE6JSSDVlVzcUUzLuYcPoz2zWEAFkly
nkaeJjf5cmgn5QdTCeNO26lo02FJ73GHj3po2eJpDonVi7PzIwHsIL1f6PSV/UbiK753rT9dT6nF
waRPeSxO/Ume2N2KqO6dX8wFak2af3K5P/rqnbgqHOLHQ2K1BDpft/rDtk+tMntgcMuLDXEdTHUV
w+DDXA/UP4f8lfW4LT8j0FzH7qLeksdn+eWleExAP2IlSIGaqP0vs1eUGclLlicjOkZXjd9tieql
KTaqWTuvAl/pN0N5qTWZKezk7ZdGUHRepF/JBZK8ShOKhCkWMhlXFFcaNPvIk10YONFRli45YqE7
6FYeIn+5TChJF7ufByu8ROV3pvZ/drz6qxEIEXE/UFqilHqRefL4mQpKa573JgCVIxncY6HS7bQq
EEw7OdK4k4PaoXIw/Roj0MStc1jP1B1Oh1FZ+4I88T78FX7wVnWts7zGtb4ebSiaGlrVW3bVRvpd
bJ3KdHNLup0qCPpAXceIPUnlzl6eqZLfdBtav0j1f9qKuwkezEnioR2OTLeVKmX7hErLaofp1OI+
zx9ca2M01Q0hlGdrFzHgncA5FzM1WHG4839AHZFe12UhGmrkCfXnIVcgaXpQrGQFM7tM2+OvgwCT
gsWkKqecSPSJj6a1z7/rhwupAkaWsgiwLcSWnWBexiIPg98Owod69EIj4tsL/k1dzI2YV0xbyX/0
DVCFwag8Br4LTCqED9p8wfuOmzBehO/ubXg0FjDjRMwzDQhkyFRQxV+N8AL7dP29siqyMQXmOPir
RWvIHQ3ad0rhD272v5yUUo/Blp+PzXphH/2HwpI6jHPrrEMGEbz+ti0zcPOzVdTgEy7xWVlVHX2+
gh3cS3S1bF+VnfyJHrBsFH21VtPde4Z/tEkD9UWpE9hJxEVSviKZmAG/6NthGyNrWfomJU8tvE9p
Dh7BmaaFWyd1stwuSLFvvFEThmjKwUHLxNG4AIObSZS/ekQon8Tgfr0ggK8pK6lemlI7yPsKrci0
dkft+BxKobdKnA4g9e6C7ryPA49mKCV4VoqREIyU9JH8DmRsMlTour/AqC9OJxxlud5KFhqGQ4vp
xZImvKSR1sKpGs0X5W5vt18i4XD22G9JpCC7ZWOgsByfeuxLGYfz5nNEFZAhQkQIN+zaKwdrRUG1
NcxApXF3ZkKZuLFxBJtAeLOL7V9matrEPo50vc1l7JfhA7oKNJsCfXRkZzV40t+gJdcUPmkB7Kye
Es3KcDqddIjChblXmG9CWZksPxAGURgDSx+AUx54Ofze1HdpBeaaPeDCnPwVcSujcoF4lnvdn0HW
bKu9FnDrXqMvtP5EupcwOB7Dfawn2qhCpqcYt4U6N9nfrsnlHbNm2QuSuZjk4WYE9OWAfVHGuvYm
akVrr44xbZaJPGxUlrWCxC6qPLMroTSFj9HCsaWMANlSjLrWV7tyXTcPLFZvPhxCx3tHwanmwFxR
MH25WGZle6Mf1AoOD1YRiQmvK+9nmUk1J5MnHR4xXwahyq4v+hKKGNk9WdKy8sKh9TFUyM/7T1p9
dIXn9sVhApcWHSlGsZMitVv5shlvij9HBK67pquYjPpjOdnoub8/k54KWXI2vDIjadmQ691LVdnw
yeW1lqWRdecc5AilH7JznETyQPD4o682TA3CyeVBD0S/JxGcPlh0CdZLWkj5MhRxfxQpgHGz/OY+
DJxBhSpJD2oNhc786KI2mcRdCLm8bHw87b1jFOt8oY86X+ddfechG2s805kSveUn0mT0dRZCDSd6
UwawIcCcYGjA8l1mjQfsrt+uUjHoCvb36ISySGK8XYDPtDHyP8UsxED2QDdL2i9A+ozBA+Kw461A
OAXcs5qIzEmbHWFTMAmfDXc+aq5XfoK+vdul00pE8UoKebFC0R1aCnpkFZC5RqFQARUYEvy9mIN5
l8As+zmXNlB5zRZPfF8EuXwEQZqP4HhAAHrpQ3r0wzW5P7SNKVj/sfWE1a4e9bU3aMHzm3g6VS2K
wd2tnyBnUMAh8XVwkOFL5lZ/Lf4kAeh0SM7KTyjy1naWgj08DEAsBbdhyb7Y0sy0DMtz4JKUQ8W6
WiEJEhHqdIG9IboKkiysIApMN+CIoTqRGNCtp2YpNeHr42s++K4kqubq73fbwXwosti1OcEALni8
MkFIYwmZcS8g/wixbj+A6+l+SS3kdQb61qxRdxfhJIO2eP//MrFZw9k9DY8CS0PkPuwW4StZYRfO
yXnjvWbHHO5z9N5fwPwN4TUWUnbMT4M7USNdM5WwmbuVkAuhZ4eX7Z+OkQQK//oeuojvZe3XSf8K
wVjgCLfyVbyotlM8niD9KmOFV/CYf/cK4twp4rffkKkAyQT64XmKXCMc3Ma/L1l2Fa8MgcsOtuyy
dhuIPoj5GYl/LAx+sstVyRazRL4JsLOvunuBUDaYQqzWQsz+gcjKotVT8bvUI+dRiFEfuhdnZdDJ
1TuQ84lvAxstkBOF/zSCA1MD0d4QloaLI0UMxC8ly69oUO8ldslFmXSt0RplEF8fK726eTAZwg0r
CWG4PDTgmUHT0m0CIW/4vejJZp0BKfJEKcSn5OlVx/oQAm8pIQPwSkgCXWZY1aMOkvt+C4Taokh9
MRG0e3y1M+B4tnHhLEMmEpO6/WxCuVrWBKN5EvTsMMWxeD48cxVYvd1bct49YQZQrYmLrU478Qr+
vwk5NN9mi7wS3XAMCTUa9xk7/poAC8NA8rhNfm9V1Ll8Ey+U2SpJgMXPMj59Cxyc2BakQxBSU0w9
QXs33jUo9Resdo1OsojcRPW/X6b4Ducfq+MfKyF0rGOrXomAXJ7qj6K4KpdrInyWcnpkwr5ljLdt
qD4zULbHDTIXUNuab9Xlk6/LPHirvQKGTF7N8SqyFQ39erwE9GcAjUIN2cz7POqxNTowQyVqgWJ0
g712yJT38T5sVC0+/jFTm8y7LEhN7nSlHqGykjGufMPUGbK+dZZHREUygvJuepO1ioVIBGLqhQYU
rg3ru/kup9ulz2S9JddQ0tMnmqHyBqqMAsWnMKMaBuNnjCd+el/pJQlEoFdnD1BF68V0LPi5aTu4
172h3tSI3bXORBgb8jMJj4c+Uqf9j7t1GSNgoeXeJSZeJ7XI0H15sBJgm9TsNVZ6Lg4WVq/6PEA6
LyShy62T6DrBOgEp4W4FKj2kCP4gFfcMc+Q/ZCAHkGAMkNhqFjcP97TkGpNGk9/lkUPtBLHZw3ZH
KIHvvqsGvWEnvzthcCmASUk2is+ctd2sqZO/Uc6bsHGpxVpP1FPEPKUbkXUV+e+90kus7k+01dE7
S8RCqMnRziXUmbuDNegor26jX7b4Sa1I6Ei1Laf5cfd69/+QWd/kkYcaTUhNEn7/rF870r27Qt/T
Nr/6a9Hp3RgI60x/pe6fHUmJeBX8TYx6cGf0xqYdgFFObGpIGCUJhe/RlsxGq5QLbmjtd1oa0DAV
/U4j3tPAssPt5zfOzhQNEFY2Se2jWA1lBEwddKxhRoJUH2obn9+96cFdEG7FWdJEvCeEODW4tJ2P
Zb4bQ985et+bH/Sh0l4iT9CaKCanWQnRujquNy603iDKY9KQ8/cxYFx+HuP5ZQphrl00WsiRLgjV
p2BpleuIxM8xXlGTJALLyi2n22MpN/3rbrynWv8oUHbzmULlNQGWRJTZh33wBsefEK873uq9USU1
+2z6XNTgW2cRAQjOpW4l4NHFBJEvEXLFdUwd/KW9UFUJaZtDIzs4zTehHFN0nMXfB9fDMRandB9u
mGt9J2iQ4NPyHG5ET0+nUELvikUUC4dqoISPaq2YzBSIWDwVL87zUAymlCCtFge9c9jLo9gdQGNg
N2G3/e65o4qS1IbzA4Z486WKnFGrRJvqaj3+w9wpJZEq0gCOcx7BW1eEijtmjcGIIY7uWn7JVLRJ
nJgWHPe5AxnVjdokFujl837qptPqB7EvwqXCOcDK+w6dFPJgw5GyNBtt896ave/lB8bOkXsKIt1Q
jnb7I8S8L64LGvbDXZJ0iQtA6P7jeiq4G55GEUHE8q+YHCKm7nrw/D83JqfP/9NoOgSjnDnOVt1B
EXW3PYDbTc6oChswaOw0iNe2eAYyJhlHTzlS+5SRofiOyA6cns2SSYxovWOMoe2vrvLysVdeI26j
7KoZQOHedIBuRPR5p7rDYimniUc6o/JRANELFcZfYo+uec/kuPDb3peZcFycdM5A3MNXvQmyY2La
hmlpsu3qqzHMGB4w9Alh/s89zXCMz7M8tjVckOVHA4ggykvh71TQ/NXV9HtVgEBs1D+uxY6sKk05
aINj8WbiWtqk2dDOs7i/0WeigERII6Qa/YeCevlJrE6Et0XesJg4KC8QaIWE1wQZhoygLlaEkD7S
Z4yu2SwZnxALgb9CZGThtKyA6GnciqXcgsKUAuMEzSIMZ9g1UW5wwNhIKXVnH+jZ9QunPNGNtf5O
ip+MuEvT9IjlckplHUR51OF/Cq03nEsQYwOOaYxESOlOPnGo8pwGx1DAX5aNWOTVNyz+pOECx0eX
n3judvfp6LKb7KbiKeCfnmW9UwjM4wSw8DxvzNeGc+o6FK04nkipscGShRss9rB5wfRRmv8fnwjR
e6l5oGYwfVyX021wD2hTU4duqsrtiruKQ6GiOUgFJhqCJ4JUAiSfLWFm7BMXpmFnz8GGjnvmU0lv
gmfdfw4AJ4b9wAFXATD5V5ujcWHOik4Mt8y1W5V+j710EwM+t5VK9UxFqQVi5p63qDolqRmFFLgZ
7sHfdImEvorVrgammhB5C0di3oqKa+kKzHfs9Y22u0ktUJDiTNe70H63i0vvHCYNWGuqZNjUly/a
UvgWdAPP2K9w2OgyX52+Nw/UcIocjWpsRaA8HbYv1PaszPZ6/ETnHKtCsQNW8t/jUnN1CY5OBt8I
6zikZKhFDD131qKw8Qv16UH1eh04xiKuQ5XueoA7SnpX25GnHjMJy9fBsBtH6F5hbGhuCK6j75ld
eO1/s7natdjyM+e9P//E087SwGYSylCPMwlkzOrGvqSH55hkw0TIycKlkGS6FaAzukoEThBLkO/+
erLlKhGih5hxeENnGIYA3vnpDQr35xbvna1rTPXSgi/0r8N/BEOjguVM68ADrKI+jATSSowSpzeb
5glmb705U6RTqBZjtbifsSU27B/5EIGX9Rp91vetyaybbPN5alfPkUA7fFgArGeFZcRn9ad9/Gsj
FUfyoAzrEICzh0hjyVLWW47/jBs6uTDooGAnNBRZ/fSkieQ0GJc8/pFc1pmAjL4r/SZpKri8gXvR
uYG6AIYtVrpFNgahJKdHoJ9qjddFx0G9i1WoHrTDXLdbo1MErqJvCETqL7viGcP4bJvNvgJQeLK9
53McZIUJfGt8REyOmXiodAb6MM9JC1iVPp87paHbKMPQud+A0gFgF4iy3XFp7GO+4+wYsu9lINNq
2I1WYoMEeYGaUQ3zqccUfNf3kMmQ3Md9lFo5G+5jEDBSI7sDRqpZ1f3AorCAVOE1akVf2Iq59o9s
c2o59Y8p+TkCht4tiCspG0trirj78YyC+mTmYc+g6OOZ4/xVIytfhiwTH+sr65rtTTYmBXy0OJDh
LFycwNHTJLWa69z+6ab9GGXFIrZvNzb8IzflkuIxsOE9qYRFA2jLwyGhcCAfeXw6S45O4AfEOZ9r
pDuFLy3E0t987sTqCpNAtcHM1DqoXnd7d7wapoUxowhCLVtoW9k6kX98FYxuuRU3p7+X1FAmlIDX
p/TcRejRz+N989QLvUF19H/uDRAgWRjiEbQzOgoTgA4iB/WZuCCek4kEVvH17/LdXj5ChQplrVf1
D0dcF4xyBnJJu+NDGkx/VIwVUYcdn5e65K+sbGEakMNrVZ11k+84ND6dw6spP+9aVrg/48JmIZZI
BMJBb9jRQ3yl0c3kUzqKsBW4DbRWReab5Zd6h9Zo75O+vvR6aeRDZPZhLecg+NUhwjvhgZzl8p29
vKJ3mMgk+qeyPZLTryRpMqV7LCEQ22hhEK3ZqYj1T7iNANNHTbAzIpJSwziTufYjl9isimqyEKm4
D8uTEcaNkmTDFMHXzoYAeAUoYFq60dWuhE5k03rGyNnaFT1AWhiwerEPBh41niJxTNMRKHgXjGj0
notUIH/oAMQ7Z2rWTGr2bXIH1IORKu9SXko86VUgchRnaNY5RyvjTiZ4SkcwUo1mWzk3jCX1vhXk
Eso2Tv6Qo8rjRF+hlBpRTUkTdtDTp031OnzvbE25w1Uv8IkkHz3cPh+/UHC9C2CHyE0ZhOTWmc8P
C/ElHlAKsmuGuRPrXlwXW273oNVcB9dcyVWJvk3oG9Ka1dqEas1mMiVzs9znDmVWEP7AlysRbsmo
M03cJn8v6QcubE4TQtJlrGhFodXQknO7YkpN23eDN5ckjzPCAaHCLeEkCO8jTeRvotKHA0qMaBxc
E6/09pLlQ//hmAa/twHUJYaBx5ASpuZzPeBMQmVl3GkPnLgf8nkuoH6cSunCYvHeQGjvyr0N6IUr
3/U0MH+oVpPTBxm7HwpnSYat2xodGgHpNT5BY8I92aGaNXAW7HvBPdnYLatO6YM4Unneg8toNebV
Wcs9cL3TtuoQWAFIf0GUm8YUWl8r3QoWK12t2kQZo/SvE3CbcwQ4fF+WNljhOdSVacRdqfGJ+dcP
qiMVYdAru71dGeBVS2HgBbU32uqufnZKcvcMkBPbk/dNIPT3vDjYPOVBYTi2tcFyBg6VCkWF8q84
P9V8xsYWJeoDAbQipSFDOctwKquM4Tu4MMG1FGbZJDB2EA1u4QBBKekFpdwnTSBgySUn3sLUWj53
SCGrLvjwk1WxkjWqT1U21DQhObUNZjYmB88F2okSFlMzY0bEw2Vz0d0q2huEjr0DKJvdvpDDEm8H
2TCdTq5FT3O1jzWe3EFuY2I40yfeTlkmMpCUNIjA56DDPCVhUB/zvvtG08B5o9Op8gL5hyBsEvpl
FgMyW4mXQN51VVyu2dco7RGjsZqMOSU26+dP1ADsT4LtxUbgLdyW6rt9Tx8Pi5h4b7apb9gzp9Pp
pslkgFj/TM5HSbMfn68RN0UgUh/jYLq/sKkUcXlab6qqFxM0UhKF9RXYWOMbgh5ULXdeIlBNtyV5
dvlqnrRH1c8Dy0ijX0ckQTFgIQ0vquVEUZAcmkg4DfGx2zmCnx0q81SaFgoLorcozD+aitr1rfSV
vcrUfL2nSuFQB0puRg5MrHQND0IHfIpKF4KpdCUOss4UR3G/S7w4K7sfcLT/NLoG37tEHTLNhJAM
kTcRsPjQTqcLhqSzDL6OFa8JJiVggmYcjxo27XOeNNd3FxI6ckGIW6XFh1rIDnvdd7yNyP3SmHr3
M7PI6FnM/A8bikuBYiXLN3bjb6McIWMkuvpS2Kdhl6THpJWXY82JhkRKwB6Ob1Re6k3neGYiMoAg
kzyTS/jDdXsIQ4wmEITcYdMzspxVXeiWTXiPCQGk/k6sLGBFw4L6Rsh8uyG9m6cYiaecrN1KrV/J
i8wTlC/dNIli+dcjhisLgjZkspvfMXYyA7Ur7o1utWl9wUwuvBrmEx2sf7l+Sdp5f5wKRf+2jThk
v59W91Sh248RXFdJscE2Qc/A0iNN93/uAhWO+o2V+ibQHXQnx667OhL6sHDTnI0cF+Fbj3MDsJ8b
zQUKGsTIcTGsS+KzzkLZAowbhTnq2X3358qai8qjVcO4MubujvEAbNqX53aJoL9ElPxn4kr0Gd2E
YPZMeJVhuBKpQOnZxjKJeWbqmfBmdVIHiumfmoJIxDUUvSlFYWG+p1hTXGx81kZn+yAddyzWeMTF
NU9xc5Mc9jpagtqI++VIA+tG6D+7KwPNcT9ynY8H2SlKzy7BoPxGMqJJMZ9x9AYGwYfMzvxCiXZL
S58OJekD/S6ZVr0XAsFUPSiOsdPg9M1WPHg7HnqxjR7cHsAL5tVRhAn7NrOslvmsSne0avV+TQ32
SHdt9dvtUwZzLbdNC76SNGBXS+nFodwAn7zRN3zJY/rDaVKV+IVAV8la9AAeQEkJM0W7Dv1YN/d0
mqI2Bk/hes1mQL/OkFsGaytn/XbTotFtutpL2FQbWM4x46Tv3r3Dewk4B7eEckzbvtK4umqad0go
zstzuII8qS1Umpzoq4xE22A0hjQqGeDHc+C0HYd4kNdtc8rcy0luW5TfCqjaU3cOxFpgUlNAZXd5
Li/QSWoG8DeWm2nDfpfK99q2Z9yXHSaM/4UhdpTpxa8/QXXjLALDy/u5+FYT+l5JbG+qENxs95R6
HBQ1tzyVwicLfsGInoz9GyF2i7DQdPS54B20C20FfY+Ju4NO/apYz8QaGhQsBrH2wQv4WGSf3yuf
cBcPDrQbPrP7sqiJScfVnTeUICZVX8EUg/KJ3IqCzTbh3jAB2axMWupfpGkqa8/NvpKAkOyAiyB8
6I7eUwVCwRCTdd+5eBN34KMXPwPaqblPrut3Pj6/FOT+Jr/0+Suy3aXOWNC+9BCdwaNiNJtmc5xJ
JaqkCA56HX2whAxmx/svCF9yDP/hp5bEySt6XAhTeFAj/T5nf3VKjrUlmlR06vsB0xv2D8oWMSYd
T8d0EdFXybSo7I8fpwq68aqJ37Viu9j95ALwYUpcNMkuiEflJu5E7LmuFI+fUV3N0hnJZRxK+BPa
TiOq43FxHTyn4G8af1yerspRM6m/9GaA9kzK1tceGXznEdzNl1PsTuKHLy+F0dszYGfqxkruk6vE
6WTL35ifcQJXlKUwBnSOF36y4NlKOE0uuVBv7Sze7GIwRJeZfRhCYoa9xLa0XhUU26q14MMLJqZR
fpNWJ2OuXH4UM3nMEkSgD//dbqgM1GSb/uYAfzoNaG9IWvSuOr7jDBCPvQWBnAV2uOKG4WR3uCHU
IZhXn3Sy9rtfWfAGh3wsX+X27oTZdWq++klYGSuw5dtoDyqmnPfDZu1rZX52MvSXto5W76pAHrS5
kO1Zqaemv1MyHvovSRCVmbdCeqd+d3njETFpI7tMWK765pbKC5iXjfbG8js9yE2YDTaPtKEX4S44
kctNoyrPRtkGCeY2hOq4pCgw+yI0YdDu0GIS+d/dJnKshUfORAQoYC9AkmBAtoNL/eCutUzXSPQV
uz4EP/8FL1PK0Si3/O6W9LUqdwf0KhXwM34/Ci5q5PUeA0sEWMF90DfJahnXsJ6qXQNvy1uETThw
TNBY+pQ1MO3sqxcy3elbQYwBEEMLxKnonCyZZKgxwA9QYLgDKSNkj7V91gdsaZnurFWgOXHre6Z1
kMrVLq7ErCg0OhCRkJWLmgdFPWASOvfrxBaSV/jJR9JitRGj2EQj2NnxGb8ZwrvcrfZWCx9ml0Uh
ICrlCCuaj2dwBDXZvYzPLbxZCR85umwiNjYsDqOqk0sLMXpMtJdeh8KMXiqmcj5eyO/FfiWevKLE
gk5My9rgjRK0V+D3WXUgJ0BPGhja51Z0Lz7++x23XrmkHdDKm0Jy3hUEDyU3fqn/OMka0DNvf4cN
wLmwSzeW4GXZUnd2K5aPanGxcUkyzJlLLsSh7MhSdWHjBGYOTJAv0cC3EUJ1AsjuXdHTv8iHfN9Q
1+HjXZ594/9XDWg1yygCMwab3KMhFBI+zEyCulJeEubN2lirwag3n1WV7eyv0TUEqgMjlQdsT78g
4Q7PqVtRTqfkF9y+LTIDVCgdzEdSsr1DZvdvd7cCk/xqh5ni0T7+KBESAsQIkJO5j2a+bkI8tYLT
vWMPxZFm1QEXHooCK4FHPPgzzBPD7XnEO6JnqXy1AeYrDo8yROF0GUNGDQ6IdFGuu3WhgyPhRJFU
x4Uy4LgivzNozuOrmnMyKWN5nOAvenecmETQYrcZovhjNJ3dgMH3/KeQYwxTITnO9uloA0FvyU1Y
90aJj22MwbxlCigD0vF2MeVt5Ui7SBuGhqURaLYS1Rclezb14D0/nulv+0kDoNLtIgZ4qPvFHYlI
+ZnOkvsybIa8evALwpScDW6PseWDLklWlsr9ovvoSq8v3ZIGeK6Ta7QiUJaWXUXXPcBdJeLXZxAt
2SuBsxGwKcPYD4HvGPpKCsasalvOPxxRM2vhhBD4FII+1/i7HSpfKMTz/rq+RAjBODEzLV0wwLpC
fb2sHh9FlXuPLmEqZgb88h57cEMi0K8kkA9jBwCWSTzzJGwNlQy4IWVLbF58eGqK1QPgNO6Tuiht
HN9wgxZygtnydAO+7/13BJLUxDpTs18R4GqOKxPaYDgGqeKLRkAEKE2r9o1MmPV5aceeNyfi0CBj
7mfD6gsjwkD5y9jstsPvOE/ZHK3YV58r5Le+OBtjVyuiacMQltEGPl5rxWCFSVbjld+K9+cli+qv
+VQcNFAIW6+SYnPUzJK7p8S/FoAlh1KQBLHCMZBk47n39+Bu6N0PGO8MbyFBLpn8uKZx6OMWo3eL
gq0dB855saVsLDfwExIdrO7RhdgPDffVjvM3GJXJojhbBt4sCe2sKmd9wYsTg7cq2qXwcjfNjs2Z
1Jb44xVyTPNRTCw7cPlf3XKbU90hgQjPhjOp8MbE9Qmv/RjlSm9YzwBQwIrM5XGfovMEzn/vIrG7
3kErx3/vTAsYc4dpwm0HfdWUUE4/lOr1lCmyO4+n/SiNFLNkPTsmI/EMLMhgR2q3Iy0Fb1Hwv1gK
ubv0wYtzEJyiFcfIR457URQhd/V0roLpnVAMpeNieBGGQ2+IyMbKkSGtCwjrsN3gd3EDgoESvpm0
n/RoZyZZ1XcRDYg66deTA6Ms/YAPKjpDDBehktIooNwblOR5R7Q3nFRonjpUp1FEGDF83Oq6sh/O
t7Qb5xaBnd7h0I65tVogo8jOO5NNBZ+SN86XdW7M6194D6zWWMewM7pICFmWzbJJdBZM1A8EhSzD
vkoS4WrLv1n5OfdAR+47QjadLgaKWb7+hiY8DRM2qEaV+bzpcj57RxH1mPNyIrrPpclplRDHcdqL
IF3oIK5ThiO/DJF67kD++gO97ScmNDzrB1canYzbTTnaCpBTgXiL1UgtruLteynn9CoBKWCf4U68
TtrzM/CwU3B5b/f4AxAKf2QsnId+YEePV4aOhqlBT7YTxreA3dmP9nIunjsiL5tjJlieqvCbL8YW
orETCfbpfhjs0x9NBxt2hr5+cg2ZY/OI3EGSu9KEhCfsZR4wZAzA3fWXD/bR7107S4CoZEOlGXZu
oJ8xZ/0xyIKlD8GQlr+fYuj6hwPlzdx6crprgAko/gtYLSyiOvWwZ5wz8DB4OZRwoy6svv12kHoZ
51pAW8saDWXgVi8OH9UH3+A0u1TfE8tuQMmn07LXQ3eHaBo+pKeJzzygA/Dp1/DO7XyBsmyFcil8
CBGUVLaFDKKkD9DOIyLAFlO7azcEq698PjCP6mELifEvUulUjQv10qOFVkSQ0jHkB903kCmLorDd
EICTTg7RMPQQ4hWU8JT3fXpbC/ZPV9FXOJ+BbsHiv4WLSk/dsAXvKtoAPgINr983PqD3So/fkfaw
NvsLRbqLAuFzxcy0s8yUjXfyIYYbaATDxrQNArU1wLMwJWRW+SNPimxlW7zuOCqlU58sOAU28nGo
etGe1Bii43wCKCNiiGDXjnX49qD4uOq39UbANZDVM+V+JMKSAZK6X2kvb69/HbS/VfzVctms1dO3
/kWC0ldJoDitTAZslO1LT0Us4pURNjCJCvLGBFIiD4MS4Vbh4W779toUlpoWia34w5KhiQMJtSil
XdB9lGc1BJCYkn84H3exZIHssfiLoiagAuYtN7w9tAl6egmSTSo4iY1mxoJ/hZGRnQFMQ/PF6GvD
SX+wZ3h1o7Q8wVZvnIKJbcuSiRPe15MsGmN9jj3X5VVrs+BUOkJ/95Atb6GwyKoIjNgK0GvXs7QG
RvaVaLmCwhIMKnpTZWvqAdXALoN0OLI+5fpLN2EGVIJHxu+miM8Xkb1P20qBJoaJ7TjrBa2AgelN
GIPHly93cHk5M0Vr3o28OaR/eghHCs7wHl988Gph457jlZFLqpVmSFNp1DYAwEuVsSQ3081er+SJ
O9W5zV1LzWYeZitAMFUcgpeJyG5R2rH1LICUociuTjSlwEjqT6/nh2XBv/fKAZ7I9IT9DY+yeM3+
nXulSZIkM+9MK2C3+NNiV6eZfXc46jtWrQICTtw4Ruq/qQh2wBxjlFzKjy4XhQH/VeYk8d3cohdu
BOuHcPWQ/WvMy9RX7KkA91G2rH7NtTxABya2CdJLPJiL373HLsV18g5Apm7LiFDD9GON5OKKh5rX
t1CwY8QFPienQVXaER/DkdvRMRE4Geo0eOwkRpP9xKLRwRQFA06nWDvZgTqs5IQ2k7yidr9hUeWu
GwX84QnQGVrej3d4JtKzTBJgMX7hRdEC3uIy9pQKsFY/x6xeWXPorCZP9mnDRBs2AB4v2zlGs6nP
pQEolkiyBhql7ll747NECh42w4Rmy/bqH9WaAVgNz8ycJkgBBsyy1MQUu6hd+BNhkJDCmxz4Gf6w
r9GtvyB6F++COj1qG9hSujZy9EH0ASzYJjV8EGpvOnW+AW2vkTScy3BG5im4msYHdDhjkt/alAkm
hpYCI2Pdag28PsM9lKAWHl2k4zCpt0ne7gpc4Nt1aA8bOm1VwiAX0SJrMBFfMsHP6YfniIR/A2XQ
MGL/Bp0AKedMUsrz7NF9QDxJBd08g7eU57K01+epgqne1fRtKZs6qnCM8NEZEJRf2M5j2LdZRk+N
zbUTRo4gg+b4JwCVNykBXDV8OEeaYemXkRyFqwh14ewiXRLSSXbHM8wiGbQ6t9/7jLT1k0MdoG8v
WjO+2rJ/EUPqmImK0FU5gz/5CPkoaCuk/EY/b3yK0foTcWq2vfVPFASAI5qNoz1/maA5IwY0cCbI
2+T1ISnAE3G3MqQOkLo/jUAhNi0v+NizSoEe/6Bf88rBjPmSMhDlpCGj+RzeH4HXczYFWbYVog6N
2m0yTNvS3DfW439ehshTQixqv/h96Rp4gfLT1Z+qaPaL8xgFQVG//B0gr+TYAv4IHefJPfgC9s4t
KKK01/idr60SY2U5eLHdHLgrCDfzi1h3CiP3uq65V/rZGvfGuHqaXusa5l5AcOP3y03mLRLEiVOq
7xKVXggl4hHMHEp6FjiM+Dvq+K3rQULkMWEBnUP5Z/9H6iQULAyHFvqMRh8Qsh8WW3gVf0JyMhfQ
oW8/o70Si/dXMZsEd/z/JUBF7ZKPkAgjCvpGRGy7IBxYOtJ1xxLGL6lQvxkg5JwD6+Bx5fHpT7W8
ALiC4e6Y1xIbybcScRil1+bOz1tcCpXH9y2EV5UO5NayEqT+b73TEORw0bsUoYdfivU6sGaLvGtF
I1bZIeZSqSbXtKgl7TpMN4L+9KYOy7fpPg0Ggdz0531v87qEufbykY/XoEj8bQ8q4oWfE0D4p1Zo
So5/ERUH55OjRokgftj52bFyi2cnr262ib8/9UAEjZr6pSD4lrsTDXxPJU9hm8r2lOX4u/4KzM8A
rhjquJCB5CoLEq2gCLBMCR53OBvDSljpWsu2yvwRlnN6ZOKuYRNpvfFpUPRpHDU4kJicM+uB4e5O
Tu7lwT71Vsf4c0V8dwjwVmaLhMgFMfcYoRbgUqw5KcZk2sClbeFnALtoHTiVvTjfaccfoFeZoLuM
THnOxKr6kE/zT30NvP8nROP7+9gpm8ldsBLMf5BQBSAxMMa4oPDh2DoWA0WMOXipScTM3o8bDmE9
c1V3+kkk7mN/M7gheAVYcTUFHuSPRAaOU1uBtN9QqaIRWC9TnvKrSR21y97W8DDuWUxUYbhj3Q72
TykEjmdu8PLK2Ta+249UGmc0/wnd51+wGYN8A0USnWYL7c+lZVuoyzzo8c59gRE4aai3ZIhKsbs0
teSYB+OIYcpy3QguvFPM3eHAd5KFrNVY09ucxEZKZiH8pGjD8YgVyRn/Wa+ohkItnCNQqpVkwB/y
+YQrnpTPktjeWNMi5JbaAxAyFgX7RmnAbGRHu5sO8k4+JGZR0WuH63raUreQ9e0OFltTB6lG2MwF
Jl6Bwgl2O03saGp2chPezXwqxi5uPqFh0A3jb/h1NB9jRC2228e6vOVy1c2gDykx9jAQyTdjvjyr
fiXkeAdbLv/HO0qtNyOaX4hvfiTfo2hBYBPepH2+9P11pY4ScqMWToU90MtdQutgaAq0rXungKXQ
p1fWsHtb0Sqw++dWzIxmuO02VniPSGFRG9MXV9FJ0J6fvkc8UaYYaD7QRsdrJrnq2disfz/Htv1F
Zr1zkkmQoFhQYTjwIldfLV0Z+KUIHTDRpkeWtv7WVxBJPohznPBo95KyIjoXImC4yEEdk2Ho4JdL
PtVYQk9AUNKkcGD3D3Lf0Y9p64oBIkvN0N3pV+dG9buE5mOqpOIyJjFfN98aiOLVQa7/kO0OHLGe
h4hKHelNlzz/nkTSAvytzo7o2cmvGqKa13/GWnZisVIhbokIkX8VOYSNmgo3OsNmLd5Pr69W29C8
pGD29kr56ivfnfVvYIRS6qTV8EdSD2b57lLa5Mx6zt4pJMPnw4zd6OMomAVmGgCQ6Dz01ADV1+b4
xOj9A88sek/ku+oCjigwSIgnRrdoJdCTK62LCi9/VjhYpw+XojS/NKRafWC+XHi+Q5z1OcdKX0ly
B/6f6lqXf98nx74SHUIh5gcM4uzpLDu4nnULpyo0VL7GqySNwGj/xclPUmsKpdESwWcZR7zgE0WN
WbJbsGq5KDEHKWSm7gM3LkWA6GAKvDI1MYh+4DCc5vGebL1k9EosWD6j8kmwt5mJztzNaGr1NLnC
r+RLJBvZljpBSRSGwTEZKUkmSUFvX/j2bYqYELauDLd4DmX2IM1JjvsBMSBuL0Du2N5W0XL65W6c
4z5eafWkzVeWSubrSkPgXkItRE/GCYvtS+brbPpKd55Ac6GCy9C8iWaqm4jQNd1lvnlWhaoTiWIG
b3tAIRKHM0G2v4hpg2jnEJ6rsP5RIiITRyw91CEa1i0S7W+ewb9PsImxje+fp99edHMtgpQwHVmU
0HpEjDY19TWnh/3K9VnSpqRlTGDW5+w/54XGiXCsogpxYlyiQhvS1kJWwTAoMLHhzLfrOZPCoKq2
GI+xFokV92OzPymW/iPlLqZ5V6nez5svlzQJKv32XA7qS3icHKCYwp16b9YL1mOGS51d81P+2aYE
X0Q1r1PLNMDGnJsq9l24b1oX6l7/t5wIZXFwJB0o+tHcP0mQlUBfsMM24QHFvmBTby1yYlrlVXhN
2O/hsWq+dUUZsm/D6OAEEgDRgCghcPokZMlAcnUMeSaOGQ2yvr3hDBQF29rw6BoUP/cym5K3UWuz
SeqvZ7m5NJxCzqiFSCnLwb03C4GwQY2rMLKpRIU1jwWKIN4tjkuB+zbLix/GVGr7yB7QXbtsibL9
p+AzEnSTBIBN2D0zK21O6QOAitc/3ZIk0yIThx6O8Wft7cIjRr0H+7twZWJLOeARr6uVwDbwRtbi
9X/Gf1In1PfVo2OC6ynfE8E0nPXd2LcGn2QWkZYE3uLqCKJLvAMzWkQDaRSr93TMe8pDCh38en5s
rg6B35m/0WaHs8/NLplj+C2WnTb14CORZFBg8svuANwZGCtKDU/w/54Qps6N8tQg9lw6K9Z40kZE
Hl29evH2rAbiEeRKWVNaZ6jwMpy0k5T3wySjzRPXf9td9f0dPfdFm7uKcQLRyjWCsUY2uYUHnhlU
DiQTU5Ko4ycMyas+B2QVCGHuzWujqRu9dmgZUlslEk64DyUykK6nGba140eK+TXW1GhAMdgi4WSi
r9GrswUxra1wasZpFbuffb2AUJVbjKJC4BTlyKq94g/iT5Jt3gdnNqH3Ds4VdZPV93gkPvNNWKNI
7ZKB0nQmpgMv9Gef84ormwqydGXsRNhkUM9SeiwS/tWly7yd575P0Yn7f9fl3Ki9oNRqFGGkqKbg
lR/OH/qI17WavWYLBmXhIptdoS4RYT+cl2P8ZQneUTtFJZLjLPL2/wHVQBM9PCb0v5MA0K5CC8tb
Sj60YBUNuyc2cIETCd9mMQp9bCYq5J4hoHD2+eRQU3HlqiKWUHVWY1Kc5Gclw9SE+G6MfXUCtfQl
tn4S5ckNm56QFeT4CJEHt/zGKrc7iTb2hznBrN5zYWSqv75ddd00SC8YYeb+dZyRbpT2/GAsuY/9
9PpBCOpYifNMiXuOcf19YFYa+hEo0+RFS8KRzXbXmLrWTwXE/RK2BnusxFjo9jIjyAIGDegUwhTp
RugkWBmD0SdUTOt7/5GAT/kH4GfWXOtwdRyndpqldW9+yOYBr+pPjmKml55eBZEbJC8wrFTApc+d
vEKYFSVC639ECI1RcLqenTKJmvKFvwxc04Oje3Tqi2wXDtKIw+4ZPDy2G3UBnN6d8Jxb3WLn9nW+
na/DLfeAKt1cdb2SAKPpzrpAYayU6HMr6XcElFwc26Eu+9SuHzLxZqhBIGbPcGOLnNI5pS3s0My0
bRsQ3x2UsGRKD6QPJfbDWdAVArTzfJyNGV14DKR8rVmHLRF3e1Ose0r35OgoioMxjwAA4eW2KIXn
nxbLPH6Ft5dRlRPCgsspxiDOoebqtfIDtqH6VDLcu5y5sme1qwzfpDwlx3Y917yy8WzhVs8wfii5
OTW91SKGykGYGztpT+5HJMldIsXlz5y+zUrp6ze3o8p4Z9FFc3N6CICWhoccB5+tK+dWwujddAjW
oDi8Ai3ttw8/W126zvk6u4UH5Rc6Kwa84lhLcb/DiDZ68PPGyT5nxGb4EV2RJ43d/myoR1R+brMo
eAC67/VdgcLYQDCAt5LbMcl1F1XFxcVAVJeym/iEDc23gltqpGitm0isCejA2aUFPeiX411I4Y60
aW2A8NVLH6MZYDKHHKwlG/hB/JaxwkBrj8kAg5NFrgO01DmM1XJjGA1N6VXvgTP682RuYaf5erdw
iOomP9ZTIdstLt+djrxlwM1H22S1kRYs4zWKdA64KikTWECuDs0OeKYLrxKTzYMTnF7wgvs5dmeW
zbvCEqzjdEJJafr86B7ZPOsuRMXKdhGNGBpoLvhkWCOW38dPuQDh3sjCqiUmutaPIaoVrT1uRFaJ
WLOwhRvJrv+ukkSpYYUsctZzPotp9UfiDpE9is3wtzSqTwCDaKo2q3rHzjNvBRWZyrN0Q8QqPaHL
OCEMM3yDkHzK9F6I1YQvmpTsoVZvuJi5K2UctbLiHZSHI35O+S2+OFCXYiZPJV32l6UxFjqdTug5
5dEBO5itSyWJM2TpvDVorp0FHizSfS+6yrDGPMRFwW3gPt4PilbZGz3nwSLGj6Bb7cOXErL3dxME
5q0FeXA2yt22iq0VNmgGEEE2wv3V8duV3RRv7dt/pZwv9TCHQUCKwFDUsjmzvNnMpymxNWgAEgwG
UmMallXHldBX7a5JuwQ2L3A0pB7v5NpeFO2sKbjoOVYNZNmvu0QL6sYNDh35u7Kva6xNkqM2Gp6f
Duj7F94r0Htn1cwnp6LyWEYWjvJDTFxLwfPlpjlR5PN1F1mEseNcydDz3RCAlu+aIghZJpuVE8ES
hR52DhOe+U+uzkXD+sRkydVgq7hzFAdMUxSqFntxrUnQbcqme8l36HetBnTSMSAXG6F0Id1VGN7r
vTT8R22/8l9GCdtPmspWu1LC4X6rgMjKWUWUpn9FUbKCnD0+sXGgTtXlQBhoXdpU06GQbKdvSCvb
g0CI2nEz18RRXBAgxvSzHpYY4Fx1BpKzg8YfjlGj4EJ1a6EdB5pP8SOj0hiLyqg3nB0p/4m6mVde
a+nA0ki+uVBWbDjskD4pPSoi1HYUYZYv9WD2+D+tbI8MAybmMvODSncvYEOJgy+KlOqV64tvvsEP
NpecbCw1GMS701aFGwwSz2jh1ARUQEeldH/ICF32i9jQxa0XoHCWE1MLy08R0nmYenVCcmRkjwc4
nODgvIL9LXfv0t9H3DTvLLJxzv03bb8fTW7F7UnNedW4up5/HpccLPvRldREFRf+hH1RomOH4XTl
O+R338EbpyJNAVD2HE9hy5EwQmWLZwiQH3zPu0UgTs26xAjNn2NQ2U3/wwMmeaxT15GQW3z6k2ML
m9n5nCd8HpMsSHsBzdJkBv0a6+8h37zI3kYXZPTOe7DlWjjjOUdFuClxkD1oBb7D60aVk/1TC60G
Fce7YIM5tA8cwVS1KhyCvpLLsr7NNknsXzcv8EkMjcam1KhD1ZLki2lbka+L7K2xKGmfXVoELiaA
8pb1HBjnl3gjzSKWgmi92Df2ghMsZ1xLSa/qtUzbS7yoPtVRzncmiEPoled/0arVuzo7t2zZPgB9
gdalGEQLUbkIavsyxoGjg3wJjEunTcOo10CnY44yiIVBfvSfnwnua75yf9wM+YmypCdm7I4YOVLU
j/7OMW0Qha3Y4iMMEk0o8nWijUxRIqEZTJQC8k+L0BJyYF4e0a26oLUwyGWpwLy8of99K72NRobk
z13fHX/vbY5l/49VzPHpJdfe2F9pcfJdrSyzYdj02n5DnlMqdENJFAf7vSJuT2NjnJNw339jLGqe
EA4wPvav1mE7Iu9IRl1EmuZ75cpudw2OM+QD4EWySHH+1Sc7Bh62JpoG+/YokqWl/il7MLcHgngM
giJ0bkETgFBDKx+NbJCILoAC4vTCpUX/aeviQd9eqF4zY0d4Yq1DEbrWOL4+fCWUGBoxW3fVirL5
+QM/MaPJtee61EZHbBZZdGJE5R3Xq5qcDPT/A0VdazHq5DEikuH/VAC/8bZrmmOGUf3kQszLnvT7
bx/KJql7olXKBVBK5YAyxRiMFFhonmD5/TnwW4lG9G9saQwpdSDg8BynLQ/BS97Q3VwtDdCNZCQZ
GELmDnpvOu9Hr0Dm22AhU+N0PTZ0nfufnr1mXd1aMFu26Hs4a4GYrVv5Peeb/oAW05ADtazA0B93
f9lKVuduoVQA4S+ttG4+8Do9LDz0wmUkUCMrm8E37XvHxfBSzoon1skxD5dYmgwgC6YQeB3xdJ2o
iNW+QxoYoZ9neD3kse3xJZdCPw/cYi+OiytL/lRV7DxxqXjP1rJRNbX6u68yMnttKLbQpV9Co1bU
be+pAYkui49hy1QDjb9LJKqrEGzA04sr/FVrFORNvj2ZUGOUy/zRIlr6dmkcg+AIRhc01fK8Cq6f
OeDsny1bPyP4W6/AqmjB1w5n6oEMu863Pf8Huj6OCMB32o6ktGPUIEZEaZFn+pq6toCecwIFckrI
nd0MSkHmTZfaSw1KVCxFL4F9SghxKV4IkIt2vmJRbLgZ0u7VD0220MNgFehPm2CpjJ0oOEbk46m6
WSxaT6GJ/CIMojPTw6lzNACxImYexED+MnP8JQexioqWW9bTzbPRSTAOmjd6oYH2CHqqQL3+sdE1
i1cx2U3ansqkzG83cxE5Y39f3QuQW1g2pCXNCrGVc/BkU9/xYElu2VKkkekpIThpj1dLtTtSoR3P
35ffZsxWZ/npPEqlGDXhH3n+L33gMjlEGMTOye64NJjAqaEJikPxV4jA5qGiWCIomQ5vLpPTW5k3
TTahzpZF6LpvzltIHXf6UpgEfbIC1uF4WULWWh6x+4Yz5DIL4vhzZMuEDHAZe3qU6fRNAMLBRaCx
CidI6MZ5Jbjg0EsQk5t/WEQPRk27oR01ZVWt1k3JogwazsA97kTe6LnszbIXRrgBv1FZKH/r4CMU
CfkNyrajR1ZmEeU/xzXEhJutb6bOFZKgFHN3lKjjtCWZahjKzGIRqRB71DUywui1JPM2M2mV71A+
xhXZLbHvQMJ0JOUxHOGWjHz7b9oRsoGznEUdfWkF4v/xw6I+rSNiaabQlfqRE6q1A+CMWqJcwaED
uzupDf7J5Ww0Dyw8rFv0eZwD/ug2i2VUyWEEBhgQqZkoxehXAyiRD3ulVrCsyCAtOFIL2dFFlscU
TCsj70HVZ4pIB9KgVU4dcEWxWZLqOjSxp/bjw28KCSynJU5OlEiFUWu8BU8QXiIaDcE/+HC4/uKE
95WmrbYq+C4G9Ov/mGuJ0SQCYk2myIo9TD4RC3ahDNuAaqRrzd3c9xhz9NP6ONOG1vwrYGMyaKe0
L3ah/iCQKtu63M6jwdulbwyoh8yQVKGu1C5mqnLqPhhNRXQsmg48N+TliKsEwCCLtSBGliUnACtt
gnI36tIOd1PN7EFjR+BI6QhvJYDNuUVAQMXxGimMm9zNzpNeMgt1YzjkEDj1H61ul6AV18AMpM1V
i1HNDGoftpi9CQXdrWmoBioxuWO+SPTUPOr4ryClEfgakGs1GL3mVrj+m9zsEhzRPbwK3YpF/aYC
OhcieNWsP/lk/N+6IXq5lVmVyu/l0xISiismevPDrK4W/pvzKIjpmgLtTDOkQVspb1ysHWUrFAQK
lHDuZA5Jl/1PlgB8KaVBVQGavv9zgZcqpmIvwzN1d0WzcHZktLgc2fk+RCQghnW3Q0+ZxiuYXoU4
nZXuRELl+2ir2l/T5x8cPKM2MRdVKU7BikuxwUoQOI6kyMrpBpgs3ctv9wg8QzrBrssnR2s1M3P+
gqv1XjP6LR5m/hs1/Wrdy2VctxVr5udXqTsg/WOl7EPQU19QuQdXVARtYjHvQ74OBH97a3ffEVTW
+AnrXCJqBVhxcvMXsuyn6IoYgJYfV7jymVfOZZ7+NfZddHCusnlc9dxdjOx12HTTvuyGQ4W7BHk7
K5D7BNmTl4T8GxyZbhjeYSLpU3ThLhPU0T3UMMXqbNu7tjJLCTIvEfyOvl8SOktRgWcwCxiLdbaM
cRxy+gjnUtJBEt18y7eQntvzVgQyaeEUqnklDkIokHvYYBe6PU8v4uNHqibLn2xhBFDZh1RgbXRJ
55o/s+8uBPsmdzCWfIBHVOY+glpYEiEr6291km/itiK+79FiTQypsP4W4ilbyZ/UAwpA54Z2V49f
1yAc7Edr+Htv9JwKO6gypljh/ZP2aDHFJwVFsxJ1tmpTyOVEQacsgtwK2LreUu8hSisICegWEuJO
4OOBSldBvupzeolwyQpRUqS7zTU3+FNgORgmfXRelv9HJz0ngWwHQgJAugqDF3vr6PjdTM8yP3Pg
ZBS94eOXOmkNiC+f+EC0GL9/MtQhsJUjeZEtSRWFYyWbmwnn10m318u5v2ni8+tLdSMkrBFuwNhj
IcjWZqr+TVFj8aGt2SbC7pBHYG/Lf3quigzWUyH/Gx7kk1PCHGdPN6BKJ2WvIiF992VHgaaEI25x
y2I2EIzMr8y7tyVFeFrA+9U+WqMbkUz66E07ve4a/1N+AAcL0cuddy4BS+sna/1hLXon+pJcDBVf
1nocG2bRyUOwIbDKyAwERIwmn+xSGg9SkE5V1VfvbfJoRluIzs4Avf3fHwW0ssTIQPhBGlrQeiiU
eXcGZfQoNATLTCo35y31YuscbFcxGsJ10lpTD6ceefHOcZa8cVXKhcjvc/WGt6TshPYiC+AF8Aoc
wwX7dLMsCDQ619qfp+ytVDMf9XVsWyLFUKZtdeiN4sesy6CeunUTAvzAI2ILt8lv8tDrB/h0unYT
qfwV3DrGUDiykcRYsiQo235qioMCoRsxq7tMp+oMLnBUl+bcJNHzlGAJ3yZdgPYimFcUd39OTWKc
XiEjjgD9qug0KUVdMzehyy1vDLDziqn+fvCT9o0dsMDNVvqvTG/omoeUSWWDgLJtpfpnlhzbh1hU
Scp5+JX0Yi255Ez65ISH5TL7mZ+48HaZfyghxUoHh7mvcv3rFS24VrZ4pvKaDu6MEXUH2Dg5s0qJ
FxT/kdgJoyeoEQb8gnOjFivAEbLfSaZDrWL1YsjARCE0BgrZP9pZMFgbhWkFZYUpHFdwL+fBz3k5
oz35MR0vGAzZHp9uE4Wh3ywYxMNALBuG7dxnZ0TXnQcLIQQrImUMRLLOSuwZ+Ebz39bTnahkFYOs
OrcDkDJRphJUfRJWyGA99HI+Hg1SP+8eh8rq6aHka3sCZXO0K8u8lwqBNcsJnxxvb/8yClVta3eC
KocZ9bnHEpyvfwvxEhzVDm5i/F29WcwEr+fWBYj2tfxU6Kg/YfsnQoFX/mf0WeYQovy8bi+CSSK9
AJuKxjQT2UMZXytSLJrbosPKrWL+DGY7Ej15d6SSvDxsrAl5nT+tMBwAw/XJTS9/bkJWVWCS2N8W
HTBAAfElVeo/uhLLrBwIS2v7M5spdiFt2e7LTTrxsdZzzzGk53qqBi6SDvbJqiQxN3CLzkdLzOoI
JBq0EW/f1psQMK2u6v4DJmHvOJ7GcTcHYVQYL0gp7g9q2wX/ctXW+8LvWIvog6ArgqCr0xYPVUUd
/s66sxQ7PkUcjPWI/TvHinGRcn2ws+WUVBFvpICNTl4Esm7FyTXzbzKrC/kczsShstlBRDwAIX7F
fLWzg86LC9uNVdU95MxrjqYrq8Of6JszEsJbSg9auhErNa2OlIyePIrScPMwm9vgAkoEvqW5FOiH
jbXdTpKBNtX/sjs98298AedQ6ef53JYTXA4s671R39RgxxjX2s2nzYtaoac3sEHLorD+ri3qzkiF
NaIPbn+pQ2muwLzuW3KrFYKMyM6js7yiKUi/F4toPg52pgAggbX0HST81S3EAEoXnULYmXCVCwtr
RPTSDcAtaeQdprqmftXP2+57TiXiBSryEvfxauOY3OvizLTMzjRtB5kD/CuqfvrjxQAkLpxXkmBW
XX+2at8XSgteHhUG0GoHMon+apxjGy8itFrKNONr/ZyH5y2LFKf6tQMp+D1GUkixvSneVRn8K8+4
p+LZhcNvqnHBJn+kUO3/HSrOpok75KHBtu26+3xFQ4Y54hn4n+5B4dhccvtzZwZopG4d05wtsm1m
+x5/z6Ug7f6vsZf0GSuG0/HCqg+TKZC8bkdUdbCKjM4qbywVWrvc5IbD8Z9iFI9COPDd2VA8P3nk
JXk1CBo/hn4aiWiEpoxpah1QsSAVt6CBtbOVEQwLU29YrYRFCLdgK3sNQMFvaVqP5t6o45zykorA
ltH7zN+x+2yxBILGCqRJIH0Lq08E0I2+Co/mAq5yxEfNjI+MDR+5rpryqmFu0ZqsKgJ8mqBM//cq
TYApb28+s+Xe4+S4S1rQU6IIxSvbCgpXpvYoNA9U0H64Ng4DZyMG0EzCRoOx6ZM9IQzI79tbVFub
0cAtTwXXkQi3ilcBBrLczNqGfQSiEWwyQuvNhBfW9r2XgBGHRpERvehFyFJk0EvwBW4RcygaVq/l
ft43L+6J3ffAMU30XBzQ8f5ZfSQ00e6+kLUaURCKP5ZGL3eINeVIrPSdol+fuewTA6wxbqpi44Di
OgiBwj+d2NAeautFPDda3MlaMW9Na7QfD7dl8JYTpf+PPg0ST9LC24vGupxcqxE7i8c9W/pquErk
5BHwkQ3vjo7bmTOmH6DmFfKhcvnsjLOELw8KfOXSZfUwY4zdAF46c3JLYCe+RfpscTQb7n6eIazY
uvhxBcWovFASlB6WJ5sFyJjArMzzZibboCqsPne7hAdPTNaHgelDGhu9JRE8121KBz46LCeBE3dk
2Gc9gDjEw8lBugMvGYWKQX3wXxtd1LSRwaCWRYH57FtqALj02ffWUvdMdwxKYZ4bCJdBPVpV3sRg
GE9gn02Z0sWSM1HnA5P4Z8dxLzwiNsTE718DnwHFOM8gftP9eiK0shUOh3k6yV9yLB8mXBAlvffV
Nbqk0KOZsyIFSAOAYK2e1+SdAqymgw01RiWLH65/jisvMEOmYdIlzkCxMcg3brLVVTPXcmGhUiWv
reVlhPTfRSwebCk0IFon/paH7YvVwfC1x+pQFS68KTjpi7k+duTShHYO0n1UwK8m41NXNcn/BxcF
PtPTqFiJSGSE3XTRnjWZx0JoO0YjvnTzTjvS9d8KYCMe9R/pNFKH8XvkMxyuUFzjJJozM+uVKPQC
6qUsxlMR+SfDqDrVJoawPuQHcnBK4xIkoMBQ81yduXa4AX2mMiS4Kk8OQPhyOpFMBSu2hyz8GJQa
bqEJWlp3lbMrgHvv7HtXaCVW9dNzGyVoLoNObMhYKsNw0sZ5rmtEgaCDlP8+V6P+fZcpLd8f+aeU
EeDE2gxjyZrZiS8MxAeOw7JUEAe+KQ21ALyvBtqqZeaOdnh72kkBJoDjCbGqgXK29CcNRWymgUPh
LiYBZWb0MxFQ7/eKm1WDT0OSGzs7egTivdbLiy3fbmR0gQKOAoepkjGNLET6E89ISQnSLaEdGxGz
CqsnZN6/RfKhnvfO471Xf8KBgbQv68mLJP/5W6Hrw3enXMj3edy3Oc6xTfQorj6JFd1TWdJnzwHa
imQx5V+m2Y4JXRFMSaJkc1RiXoSPg3Q8LB69xBmbE4Yx/2hT0YdHK3rYOrm9aj0EsFGm7oMI8ioK
nBD/OsMwTBJoz82Izmf9WchT6jCoPhaepsYjFsFBRx5bwYKejQYxRU2ZV2no2zELjIdMJJ2H4t/t
HD5ETayX/izheX3HgphL3wkFYF3QNJmDqEzmNgNVySgV0OXMX5sSYFurgOF1QkoPQpd1HnPxFBnD
r+xDBIRF5KWCEC1nbG6y64hDzU0mLHc+MfUHWMwPTJbqqQdUjebriNAMb/1LAHtbvtzue1c3Vzb1
/4BS4bSRyUvzajY9RlrSAeK9bEKbq8zJwW16WFXSgGM57kGRiFGbDU45vzJstniqazhzGNjSIPuJ
SfJP5+CIqhFYQD9I2JIhbFXJauZcil0QYUyXGng8dwpVRN1GZJgjvynAzuUARKu33D4XhPvZSXlc
/95bmhUaEQiaVEwhaYkyKrtoeAB2qv7Yax2AWpj4ADutHxQx9bUiUrJ99CcLRVU6h9ad9fE26vrq
pSE09vs+n2ByxNGqc18LK7pjXoXnLUuDgfB/3XegbeTzzf6JOESM3fuKIF87tve4Fy3NdtIvxgdo
IL5R+vnDTjaq7uiqoSis2axJT6dF122Cr2bcgjkzHyhv+Fs1x2eME8LR8ScSHw5KWnz7LB6u/sma
NQUspgpXauI20VAjSs/uN8q+2Eydz22lByjI+6T+l9/4HexqPfhZ/bdk0f+4R1ce6yNc202RfARf
6K3wsJfh1vs2+gxmKNwp/xohapXGryCU7dQevohJg3U3QkIp8IkMdciZxNSrPQyPcBnZyHIoEDly
UFtpxfk0fHMDWismzqBaNSMiTTY2YwxOHgmCgkpzq6gkOge46TUt63rV+gV4Edj/s8hv1M4+SFno
QEcZBOSSkoBxtdIOvTLlFErJhTJUrwNFa4a3ug+Jy1C6ANO0LkUpIhb4Q1lc7zk3VvPAC8bRXjey
RciAropBgZB1CSpuqHKOYlU7102oel6MgIQt87GMxQ74ctORROvizYAazhpNaTS86JN8BZ4ebeus
+cfWfH2fOyZ4P7iroXhRkrMEEYgqZfMswop0b4eBXt3J/nsOsL5BaLp5AtgaCCldhBp+l0glrdoj
hGHP92RVkqMQzJPtml9FSvbhkYIHqr/vUnMJgqd4INBQpd62lnU3VCy/jnlSPecSifhWLMeAh9bk
VbOLLNqFSJ9bdmNn3EyqpkyfZxI94He2jvRfMMgt1il3LUVKDsoX6dAVeiOKeBySpr6xsCjvseyB
q3/tp1WnKDLYGg0Sqk/zGtRhbUZyHoWO7n34U+Z9N+yVfXmzE2Ejk0oBcHKlrhCDMMnhcSdo3I/B
J8ZyYZR/1ES7n2zNMKfcIkidnz19aeF1qJgKCmKOpONNEPN9WgR7k22iU+G4wwMH610XVUVFuoo9
FshIjdDEUveIRYiVuW9c3ah06crvYRJzZcGyE36fFNib0HvPqzSyda8BOLbq+j95t04oakNNHDzN
+VC9drf9FafIwWu8Yy2Qq4k/NKv0l8950UvT9CDsm/99oMMejRpNalebJJ0+Jj8HtcgSZi52SVF6
A8rC3aHhrpXnvcUE3V/eh535bb5HU8GS1zALQhrMoVl2uIzlaZ/aiIT4rf8QsXBQ9i+pwn8YdlpV
ByP9rs15HTTGXqWNlu9rtoc93YxQm7YirGRSD6bWLPN24OSIyIjnvBgaNbbKX0AeSm1yOx244te7
ofeFia/ojyKl0QOSY4J8yHWENxxpCEHkcxQFTKTXdGQ6dvoOPUtoCAHfxcbR7jpmKLa8VJjxIA8+
5MsBU/2fAn2mdxiFszoytwPGH5t8HIeLlU8FTMxUZmQBCS8739/rIx3lEqmqe0fP+oN4Gf2DmsmM
dOeRw554ndrVAvwUgLPLporJ+ysJUIUWOUauef2BrG9Z1XNWokhlx+5sygvgU16s5466kgMfMaDK
rSoNKsiaz34d4OhN+BaJ0sxvG3KrVCYn9OoFuHmdyaImNqWX2AYb28av/B4bfkB5OYhAunHWgJmb
RBv3Wu62+cQuna9kzsmPzfOQNM6QhBN5lW+c2TSaQBjfapkGlflBeMG6SymK5aybFrat73UnUg8i
7ozYxvW5Z/ljX/OjVckSM1y7VUIlS8Uh2nF7G6vqTzsqX5eCDIbrNOLgM+KgWYQvNlE6wWyjFGfq
xpBgGb6N2vCEVId4xTDaWUXcBCo8Zb7bofgDaUUjPNR3u792ZOneLlgesWOvkhTqVqJE0wqpMlfQ
DM1FdrPE2+6lUHbkuJVVLNdcm29jVHbDBZo+hpXfU3Iu5juATXO/lsfY2586BRIMWGo/QVMpKxCq
F+DRC9343Ft3ohkt2GrJOmeXf5yMzv4pLR0falbkWfP79d8+IgMmygAzcbDmEg5ng+lGPRLXSjL2
tmiWvaDsShY8gHFKbs6IFF4pxqFQ9cw3JFU4hznXtIg4MCLIV9IGgxYjlAWk/ClaBYzsTW5aK0ls
qBsaXNclz7f3R912GAMEjIOpcNR313O1Z4T5zvDYIsLsTmzOsjv/idOwdcaNgJPo0AJH7ohhi+N9
wtMmYkfiPjScCrfUuOgfQqCLjxRDu0kpdHoBWNcdZ2DUAEKsKd4I0p8AlRcKdkQzx+i/tmEsAs0L
Vns1ypsc0aNEMJAVyKQ63h6PqVqz5J3VZT0gvlAMoJR07cfhz9kELb3P6jNjuM5GyPJ4Rh/nzZV+
xDPnNsC8iXsTj7S0d26rhpccZE4u/8nJ6jx+57XPFCbRqXDSKRWNBcNu/0KnTn5LM+dcDMF0TQ7K
jmrgpPxKMdsJIV+zztNjM5yx8zfAAu/T7pYQnFOf5A9Mzunx8+O5QABETUt7aSIrchbUl3ytrlhs
KWcmm2b/SXg0GEfKLvu7Q7iVAFqDVpZqh18xtqEu5eaUbqH5lod1U9v2S5FOZr3c++FImqQpxtlq
4tuI2BJLvuAJRlhsDDr0WXWgRs/ZFk8iB3vRe90/ri4j9IlyvFtuJKcTD79RuTBXO8DikIVw9VdJ
W29d0kMmrax4lk+cJbLGhLV4lZ35DBgul2Rb8SpkxaLEk78aXkDAq+CfaKcinqCXTwi8dBR4lbTx
Xoo1LImfOLvjbpFfWkAmI3q/lNk9FCIkuj5v5kKzX5jCXubZK4UiXr68G1mMke8RGlK2Qt37WXA3
C2Dz3FpQFx1fIUCXrZ27New3A8yJrbjfxzhKntKcPWvqSh17kXEXDfXWD32Ho7e1yi81AfEDsJKe
BXL2n8G82gcgPyNw3S7PT7OWOdsW0NSWiH1IchRSFTYIoqQmqeVABO3y9oEzdvLMY1IciRKIbG3k
LpvjdxV12EqZBcZgYvwfBMJXUkWxp3G67ZnSBL9QhVVpey+2klzHGjLESjUM8v2xvnOww+kK895B
ULXaVLaoigqppTpNUNA99ysD7W535zCSSmIyysZ/MD+PZTf4JX22FhSHePQPhLtTaUJNWESy992v
Vko8qzHPl0zdDtjKR1Af0R3SrrqP2u4z8FgJMygndPzr++SVMFo+A6fEHRIllaiKFmrvbgBBmO68
xi7+f6skZHd8t01h9pBk1GQTTqPH1vGVef6qiD1AYjm7PR0yV1RfEa+bgKpu3PZ+v7Qo0V6VER0x
yCKrUlVX1uGZ8XnI4p0Ie4aS/M/FkSDCm+z9YMh0Q1rJL9fsNgG0ac6NcapXX/u6CzP/d6KXzgW3
yfvVNApdBANjT3gKM4iC/v9NGscc0NVnJVunVUaAyyTmqtC09y8+eoxssdl2FYVl9fupWgOOVxuD
kicYieP//E+XKK+MIyTGo4Tv8vSsI7OJZcxAFhjMXzZQQFOLao+ym/N9lFTQ0VfbFuZ6+ZPmjQwP
YOacx8QONGL6RAf7Ah7jP24QKUHlEEo3PKso1sgvQc2bZ/hfl0/VVK6XYudTtttUOgMeGFZowRQM
n9tdmMJyTrE8UMSancPdkENUmKpucXNnW4nye2w5vBkJM3z2GgGrcHPtnZ02VIaXKB9/UNRNO3H4
q4LGo4Ha8rt10zRZoG0SXfJWxG8+sdPPmiDUEi9uycJbaM97AE8mhsAd4NFwocTKtAAdYOc0aozE
cNorWFNa203gWFziycACJKNpp51l/Zf9Kr7eKViUZY5n5IjmIt+dDE7BorutSQd2JSZvTS7WdaYr
xuaWrDiIbEdVtxybHzSCAXYpP/GFAyGrO2SsDqgBHf2EVgt4nkRYOwz/oQM5hPw22N4ZFlDs5mUB
jCNDXbJJ+sDLfvCZ1vWcmUf4+HFWq6UeVZfry9eID0KjbsWHnh4T7xsk2SWq/VA0f4QnNJCyooix
nKysqgSAOpoBDatmkJsKUX6MNpVpAO/4nqS0Eey/WNm1UEEObTV3DGG7N1ZOtdZmrSW4/oYPYBTR
qc278TnLyUETd17PzZOe9TR9SDFLdZeSM8gAclE++vu68b6Aq3DDjDqRb+0BieHpbvN3c1x4aeyW
ho/fgFZaH6JUAWWLM+JodhV4AiyV1fWbsGl8gpvtIPSrCJ1vUpGcUhdZ0camO6lPGBhiU5SyAzqb
K4LeM7kXqpl+mdy1LvGYfSFUfMIhQOteoUmTReMJslZ+wSmUI2eefEwuKA2+mL4vM0S57DTJVJtC
44s3t+NpavH1rRg7xGZ+NfvrPwbuRpKC72vWD5oJUtl5Ml4XMS/8DZGY8bpUxDFqNrei2u0CzQHo
cnTjaTmW/nsl97DMabqvx2W8ucgxml2GaQWoyDqytOqxLfnk9y+avAWwe+O4n5AbbdkWi9pilC9q
zsSPOHtpSAOjDN5nI4qbfXJKn7IX+1EYsV2MDpm5B1fog3iA2l7HSTH6Cn1CVpnD4dpslCBTjLdi
Ko+pE1eVYjoTj/JWsGo1GiJqa/yCiJn8xb66YR5lKVmnPWNxvALDuCEZNQYQBiZFq+i/lHpuwvla
v09qxLMzXb/D7BAWiHlpyYJhVwUl3Zso8r/30WTDD8aR3d0IeLVCqx13WmwMqZKSnbmVVqFIc2Lh
F8i7H0543pAeYCcdfJMahIJ7Dgua+fOTr8Ngcy+4WlBiCUWJmfNBHufPAwESaGE1EiAzmgCwF9nw
mN7XRFLtqhk7thY/OCelLHXL3NNG/8z2DtSgNBR5KXQmi/mJjNeTaVeufI12hTnNFw7mGGtWAPj2
WbT4Uummy/Fyx+9pGbAPLYNrkRziArWhDeHPbLcyW0nr9cuAs55kLnXruSp6iv136GZ7qAVXKoMD
Rbv+4iUEbEA5cnMiLd18eGVyrzSpw2jKPMnaSHtws/eECa4DU4MxpbKycYPfOr9CTCWL3ezU/0y3
h1LILKY0Y4GUxD6l9STgcsYJRzAU8R36bzXv93s0cEz+oraY3N1zx4pD4q2B4wSBpth91hECJd6x
k6dM+a7Yj3g1REN/Lyg1zYYKHjIi7LLaSXXjRBpm0ltHKSdPlMJgzOWhsiuhDotqYbnfpciQXuyv
mHHZlKegi+dFAU2JP6oP9Jci/ygYUZg4o/2PxoSszWNigmynAC6uyBBlscjBMIoug9dnDBfD35uR
jeXUKsOHltiFdi9e3OGRCNrxMv6Mm5dimLgRaE1BdMMmljY2ZbISjxhXf4F79InELsvAcEfN3PdM
tEh0XbFez6LDUe5PPI/Ah2CUNuuYEtLPRJmF5xf1AwADC98EGV/bVUmb37E9OhaB2/J2zYrBJEkN
oP3hSfNCNC1UdGKgH9zrQ00vIVSlLbzA2dFTcE+5QL8/UQ32l6FUk564Kd5xLMTyZ/YUKJYEsGCm
AYQeBocWRjxedrunrW3HqY12tnPFALB8ft5QG2rT8O+DFnJGDnu/+jfDrujQNlFQ+w59UUuyZttf
Qy9PRNMzscrMxmhuieZWt65j6T0ueAn8R4J2GS5wc6nueHf3A8diH5UWqY6ND3RfvuqB0IKGPbQT
+9tdLzf9+nENS9Xj6p9ycdpF1ZTH9UD7FWWVpO/MaIggZS8xgBKKDklUDhs09JtPgThkCAUbUYQq
AhXLJLoyb5rrtzb13YnS4N+y9lkYVd+Ts1iT53yMbAYyDdWldxUxhnlzkwal7Gb3CWddIDa6OrdO
A5bnXj+wOcttLT0eW6d0bz7qFy9aXD/YhyUQhRJTIH6/+rPKsat/5WJthkJF4iiCP0nN5yRT9RXg
HeyE3CnkDfQ+yAF9GMLgFjj2sayCLPygCIjfug+fd0/G3fZl9uBdrGmEFl7i38T/2X5OgHlmVjVp
eBjHkyR0bUNE2bG8tLV9dDQcsf4VE/bmzee9MTYLPP6MzDsKrgT9VdF1cNFxDsZnWtLvvYUb62+A
jZOFa5ovKDrPllM0SVYKiHLYIY55BqNKZReLpfAsuhWMnRey1+8JhEQaCV+C5QRh6J1pGPpRqfEj
6/Er3bj1qwNl8t8cGF497bAjl7RcanqwsPb54QmMub941LSI94FJ39CtrvhdCheDQONdEy7d0WLr
Yutrp3aSpO7nxdqJoMzpcfiCQYsoOJqHL3NnbmOY91kUF+Z7uweJhf8kwwOwfgwviF1+LH/ryCdD
DX8GFK4Ufg1UrmXju4jslSOVlbDbAf6+O7RxOJDAJlUwijZizRn3/MjrX/+atgfjQg/cM/RkAYJY
4JQA1i/RyKi1lGqixs83tnZhp3eQ5qUVHvfC4rUrCe1d1RisA4Q0GI9DiqdJoT7irgBJPq4ZrMGs
Ie2nVOJIS+xsez0yLPN9DSDxH4Clyxc4IoYvjLyIo3scU4aVRVInpgqVKEOxDbElzDBzoNr2yX5w
C+TN8rtysEbF6xhXlNrGO9aSCbjziafqCH0oPHNQs8bQSj1aitbbdywmQnpc98pQe8rcaNuxTKnu
AnY0OqjgcUtjC2z3lhYGHEKg2Rvn6fGscJel5CRoPOW/OZS0oFy3194X+jwvoz49oDe+VQuDjrl3
ST4w5Hzw1OXFDKCfnYNu4qX6kX2AF0CqIoEMmm6M/CHylrK9JKduZlFm0SquSrg8VCEULQRT83k1
WnyzpReh1cgJoMpVRGm4mxzSO7/fnZzQ4jgmGdA/KWUXKWq/P5ymvmyin6bOGACFhqdR6SJdJzXN
5zwfQzNPxgXNuCAoUPLS26ZMDea0c899H7JqBQ373BVwGMl/fx/47rpqxH5xO9POYN/R8RtQeBXN
UZYvfjO1lxrjcZLGmrm4m2Jse7IiJU2rrmCPioMjOQstJDN5LsO7JcAQOY3DCVzkQyu5UYdQDPOl
xPk9KI4eekh8mMdqo2XNR9q+DvtBbofT+adra4Bdboc4dZcw+SmU5LhwkWMkPcIzUKKQZDBKS8NR
ok/WXvR7/4fEcTDO8r8wjoCDw4yVZCvN/AE4t3yDcq0q7135T3gTtiqrLywTvn2qJdInQDoyNZ8U
IXafNo9bqWHwTE4amd065qafQljKinODaM06eYdT5RlZLLQiI0FnNujzkSA+nt2Oe5AS1lxVXm3M
8qSLcr0UW4kUDvMTYctdjz9FBLDIKJ5/ssre1rzyyFAZggduarTBxR5BbT9A2o8fpyuz/N3uJAqo
iLjgUz0AEjFWze8NPtp/jat4DIxrxQD860kxddf/FmlUDbRaYAPuO/wer3QVCxxeWxJ/RBpQjvXN
Eib1WfCMYHH0ZjeWm+Y/Hb8NKh/BshLF9pyPndyFoCLoQvbIdsKWFveAczn7TaVt8HZBMiZAY4Y0
BGKtJUp6+Ey6NxaA+ZF1Av1so0QPIhD36GhqaFdO8NOUfCbH1mrUm+ViGi5c5gwGIyrTOxJkMcxJ
STlMypIqCE5diCgYohaWLtlCdnmgDcBdG+EBQrh/RRFgVZ+0CzYQn7X41WPQ8zqBuGbX3PlesK4+
abIT3Kd3LfZYlD4sIL+D3vE92OVEReoSzaMgoi1fi1uN0cIb4uqaZhOAh9TwWpNbgu2tVoubXgck
kX4wG3sNJLnSHrVnvh5UUYOzrIrGgMCeBa01unsNjlfm7iiewyPIHqn1N9Vo7zoQPYV0Em9sqjx5
G9S+PfvDCe0rPv1hODXKBMZwFHNoqFCLuR/ohw6OY/LvsnEk2OipWWj5m/OXd5Y6764UH3Tq7php
sw/NaAoosNN+NXhQ2j7AiQO74WVZG7o7F2dvOAT0G/uJIe77uoicZEasqQmlxzTX0Jbh+tjEl9ck
PqcmCHfXzpbehTvS5NnpM5J2M4mXm0NxLfgzRZcwSUogP8PliYH6A9zDDJgx0nKdNw8m8DMuRExw
y0SXFixCBLStkcu39WE4w8p31EF3K0mo9B8MzPeDPc1wqhgHaOnV9IXsvx6UjLCwrGNpvtAC5Pbz
3t6Ce9qOIRYxlI4GoxmYPb/UrP+Dh5WrlUIGc2pu2SKjfbKRK3lGsFhwi/4GGWXCm+DjlePycMFW
IPsW8UDjqYejSo/VhTv6phBU2zEnG3xCtGyoLdvLz70x+ic+1QAHNLJMrriWeOEtVB8lhGKyakGM
7QvoIhOu6bNG8DyX9Edo7DzAAgVL82tC49LUHMCBGEtVpaqLdofSONzH9K7ZzUOrcUw7jJj5snJv
Hdj6oXx2ktVyOuOfKrWcxWXSffC93c2nzFHIruzaSaEvdDWGXr6jB0uDi2KqIaFyRxZYAHmCjzl1
tBUMy32+MTWGWK5gREVAsv/r3jEnn+JtwXF1AN2hOFUCqCxNIN1WCViVfPnhdfJzsMBoyxr/o5LX
sh5OpynoKhF3ZU8V+L4dcUTPUfoZkxeTnmkTncjURoGEwtJ1S6dalLZjBbRzt4pA8wah8VJxJFF4
lAG9lOgOO1Ii4maZxMIlpGRCop6aQ1ikGSfBJdpVqbWlF7NZHUvGopj2wnMasbby7CeVKp2vvgD1
HnzBIjhTJm17vSB6aY4OE9MvL7KgRaEsQkvKdCuT6kY0OJJ2TEebBFrIr0XKxgomYcvzzwvEuoD0
z9ketdf0EQpkcS82yNDG3riucAiEGh95UvgXVPaR6y18CCwCc/wwzzYgKb9eFf6FYoY+WTzEAMQE
AgrqjMPtFzvzNd6ndnqpIl3vOCXctOdhuYvD1t0lwDZJ+nGcuBdHoftGSgQrNRALyzm8ZfD4VnTT
AiVlvyj/Zbdo7RxsUYsl0jf+jEunK8knC6xOAcgA0chKS9irLidDhV2y4gEU0WPT8vlFvF44B4Gh
EB0dk7daEst6y0xwOUT5UaTvtrTgjiCDFu0DACs+7fVfOG+oOSSLm/J7SJ77RR35+/Vuo1dHz3NA
BG3MHvwa7+qulcQ2y9TTvRAwUJH/ywhN1CJmc4d3JPqFr1JrZZ4HNSF/hFbxfLXoDuST0fhnzM6n
1nuoiNcVRQatDWgYwvvPQgP04WDv5PjIKxCRkib3XaxtHy/NAX/AJohLtSaqjmsrDTrOpFviDMb8
goNK8kUVWxgcY3T5CtjM8Ubfoo1Xe9FxTMbqDRe+tuOO8KY3Ow778HUZT3u4Ou/cLyRzjVP901uq
w4P7x2+51/d9cnGtMvFfn/AwQfCT1dUtNpf3C2hKRux8sOZs33ggrfV6QLeDyQh9MIvXrnW3VICp
FIwGs4Bi611g1m4HyLN33jQbDI0ZnaKQuk4tHALJR3bav08CMV3eJhTBGGQPfkTbQDNb1rLMV58l
6O/cVgmIMGdZKFWbzhUEhYKlbQSzrwX5eDbzZVJhLc8A/Pg7oMjCZpEEo3sm3ZJpJ651TjE6JUFu
n2k+pbMW0Ir/rRAB7q0k5+/IxLzI+heUdPBWikSTySKJ76z6QWsQF6pUel12vE3KcaPvquQZtHTW
WW9Ztuxr18lY0I325znfw4g38HhfCZ5uEtqw0kD3Kit0cTVJcWxacoEsW0TUOyCoiTeIDgSLkD6y
wnKq3rof7mdZWCA37j9GQCFHsosCwhtCt5MqMbpsJ1Z+aO6KZ74JrnECfn+aO0LtKRNbGwaz2aAM
NVj2qrUmUdUxNFBh8r1giuXtJ5jHs0T1/ndCe2HJ00sol4pNgVJ+verD8DeG5zWUSm+bQIX9sMPD
X86nehcJi6IqHKBuxwT/6m98r3mDi7tYvuCWcONDohIa4EYyGsWfxg546/xhy+HR6edgdsiEHLXx
r7ExXhSPyNs5eEuJ6KZIdQX6uHwFJ9kAaex6ABcE7wp7LBZrZFa1qlZ6hF/PIf3U0Cu6E0uCib6s
KX7m3H+1zr4gmQW8t5iGow7lGy+E3TRdaH3LpRpRsXMjuYaTbdcYD4uxwVCP3ojs07jL7ot+F8JS
cHhTlgTfHKP/hf+oZ5kagE2ndEp45e7/CgTT5O941Q/+9aHF+G7gkO2eXDD/3syifQuWLZbXNLs7
jHTNdJrihpl8DAzFFwVgsvTz8qX7PFtU8WgXBYXsatX8pB+i/BLVLuZkWUixPUn6BZgNBZwpnxLL
9cXLrSFxNGyvLiefDEttkpUmKEPA9EuyVeVraWfdxuvBHO7OAXXN9QOiPJEzNZJ2Q1QGybrEHyDa
thUbPyJCuE3LtXxy26rabaN03kPhc8dHkELWDVrN/tb7Fa4aYgHvi270a1o6hleQ+wPfyfYU5lYY
vlzzUzTlt3V/31eBhBVpTIWfXI0xnfXZ+4/bp8IwKP/a5a/vbiZx2JuxAtr0sX0ZGzPPZuFs6+Fi
0iR9ui1SUqWr+ptx3Wxriz02rC0IAb5NUwGRqE2pM/bgmj5ZT8Dz1Sx/HRBxGUFSAKvxpQvPhewP
Mef8wj1odoOYTatMnIFNe/7iGujDQyNMYh2LHWraLbDPfyx8Daxu+03TzvcaAs3BAkDI370lb88Q
DKJBON0hAPaTnd487kKY1MFCprMUcjOdzBw1O8ZorsBkxztgRwGrpFQhTYvQ8ZLo4KNR9WO1pEzY
VcMUrba1V9vQ3uieQuYSp9+tosrCsMwbu10Lai+GRaJesvmcdNigTklVOpf7xhBZJYX7Oref+v2p
qdMLlQ8M5fTNou/1OFleDZJO4IYSrFmdB4CeheD1NQOdR7D+iNDrlQBuVcEZOSFshW2SDIOfIxXh
DJ6sPh5ejXb/s06Y51IhZLd6UrKbUNz7CHA27zQmTTSGl+ymc+10qVj77ZlaKXD5MFJSfL0VSmIf
Zwo80Csyr3D7wp4T/fCEwrwH3gTx4lxHD1WynBWIQ/VdYPth8kLD3JSWRl9io0B9pZ4JZftFELr7
p6iZb9c5+e9ihc3iIYvSm5JIPnw7K7SFybfrjWnkwv0i6WObii3MDwSkyajvjsSFoCea8XPIHbnE
pJTmSxXnjJS3EJjeJ1wWJRH2NQLZZPewBdtpHoywa8qGxGgpf6H8HtdC/GCvKzJyd5IApuXzznTQ
QB0wfBzm0KX/ZLlW11rnQGGiiMCLXLEiI/h1wuOxMFZYo51v+gXfZRrtoElIUxsQV65U2X9iUn6M
Iig2GBNwl8RVTdk8tcnsQZRyHu3fxW/dc28V5Gp2U0pWaGfqDCLEDmpfKnEsWQ+qhM+fKPzxHvJe
2wK2XaAepBwZCl7alp6BhYJtCIHb3L74qEihlboUYzkAZd+u2zxUeU0EClfFrZXBnH0TRT6pQIVa
3PZnrOX9Ig8pqYlaG5HQWefCVvA1B+7A13D8CIpumw72RKE1G2gBo4b4kB7/j8SULFlHaPlURtNI
3kBvp9t+q7qxZ7tIgGLfKe1wUOEEj9i5NQ9hwHE2xYNUTCku2dSI3FO6ZlJohR4HSP1E8sbdnv+i
AUIIsBfvHF01n9G2IKfm88nCO4HtKLXpvYGhL+Y9rzx3kzl8ybQ8dYw1fFnDHZOaMTwbmjXaNih/
B7hNEyBGcFRH0ewmWLsNr8iUrIijanp0f8kHVpCh2n8nXaK7DX7gPUc2LeFzO/nXKt9HbxDOK6M5
LhvJ6MHPrJzlvhnTMwXkEZCMoc7Jyov7kjXGOY4i4r/1LzRlT7NTYTCcPg+noadzAvov356MtC7p
y9Ss6ZIM9WWdg+YyL3kpAFvUgsfMfqcWrRPqZFGCwYcp2TyWfVyPkzA3brKHCU9Cn1J66kS+R3hk
vYSdMLsVix0P2fBRT+v5j1IywRBeA2n6z1ExRyofY9CB0gikWLLxOvm62exzq1QE9y0ykFNPoRgT
Fxd26D5KoD8FCEHWvtmmUBHHO1o25xY3bB42GH/gj9ASQvO4LGgyQ+5CnUDkrx031Z39epdqXO4z
pBvmhw4UWqxJXXXJKjqFSGog6TCpP/r1eFjFty+ehCVNkltFrPrcNC5a11WVlsisxr6ziJOdFy9R
1IVmLa8w+aiq1XNxpBkFxPWMzFMBJnaaUvzj/q/2/tEr6gjei9IbUkvGtGY29YVw6BqqH4VRORIH
uQp41CdYGEm/OHYpx9sTVkU+5Gz80Ql2QOER/61d3aXn02evxU9AytHVbhptmFsERXpOrs8UYMa9
Nf7DUy5hItpb5MvvdYPmJ1Liy1nyZSo3kcY6eXK8KBiMbGTtmScDJoTRyo51b3YJRfB0Gun6Iwv4
eodnfxd1oDOnkXMmXaXGmvyrnsdNhS79sMsv64xNgTTE+/NUohO1nRWXLd4Tgu8yv4UwhaOku0ED
4K58OkJFudOKNtxYScUXQWMTqqxkIU/jm99zGrWNZ5OyWrW4Bfh6eoKTYiTZDOmmA2PT/g74Lyhr
BH92xp6SS6sxp6LW0dI4suOiITHGTnN3z8nV5NRy5UyxHfWv86qMIFL6DBsEM6gk1+JWSMEpzsV6
e79IMsasvuWvy2e/NIxvzo8SeXXJV3PF9JhngHj9KQl7vmROpD/LVVIYo6wBvfXTQ7jXuYC3fph/
uL1uKUKggOPfERWVMogS37BjLVBuE3BuYw+ZCW3juzhhmxxRWIGTeLvnrcYQR4k+xl5eYB3kOqJg
Nwu51iE7gQy6VkzYdim2CDBo862ouXv6y9veTGCwWxmG8Zm2P9EqriyloVzf148BoGZFh3YPe7uU
H3R1vpVVsGZZbw9M8wao3Y4DjxuyGhkW4RMtd3qWwNDN7GeTBw+R3ULdfXQbNjehpcRvkR2MK5oQ
YsnJPvFZ/YpyKgRUulUs9lymLC3w/EgUpLhT6pqJQ/psVYxfm4KpilR6qyeq/EFOqJg+nPefMIQk
DTWuYiu5jM5cdYm+kq9UKaFpJEugF4CyEiU3LRf2OjDIXmjd/sl5nILDIFzG/S8KVhfzYpeKKwrd
wqbB0MeYR2wxCUCIQK8PfwjDjeZ8s5xKupg7ENLEkVrQBCk0pDdYLo0E/7fSCacmRrejupOjn1lr
7KZ5ZrVVscS8CiArG4xI7GAVZmCLWzt0EjZzxJldgVt+FK0jW/nnPd8dfqj0UXEqv8xhiYk5S5M2
uSiiPSVf2vGoKYm+qsJdcrH7nar8N8SgPbbeGeVoHrmlG+ENIlDxWgg5Dt2ByleAUe/+FvzE/9TS
kszswuOo80IxzANHs/OOwtFVEsjg/f3c0ixY2J6JESJDxZBWmHcc779VQqnaoXiXF68nMbs1Dl8V
N62GvqvwNphg20yw+tZXgRwBBL2RX8g/NWV1bBrBz5zYql8HUS9GLaXaGJqQFnWIEHyVhBN2Uywl
LdyDmwZUZ1D/xVBxJ65tpqvr3wlTyJCcEM0ZggCwBgCpqy+V7h3PekMZARR+hui2E7vdhzpcJS1p
AHccIOHZMCRIvem/X4CB4MVs5w0bMOQ0dsFu8S1yiyBj8V0K3lQBqq3zzho621v89NSwixH5xXa4
H/xniqPKUuHphCnVePWOX8qMVQPoV3XAGKPukhuAiHg+NQIFOJJJzNxnfq6hlD/obEOUD6RIDKRn
W097bcIFvuyPBEEGFejdLgfhjgewCDVOZOJyMO041JnHeGZkKbnUKVJEAKXAUS9256YihdCcViFI
NoZsMUT+6qDX2yom7DsZaONRkxYMXag9xWH0KidKP6K0r5YD7zJCjpJO1aCadpuixFUX/oI8hp8/
H2TKrRwn9worgVSnbXxP9weGOcns4tII76W1jnbeNYPTFt5EkbR7v1SzRV5PBjsKZv1zDLrIHIxI
Hz6KOXzdDD+TKmKZsSXKjfIoDcZ6KGLBQrKrEl9D9qi9chnw+2pmjuq3MYduypghVWed2h2g3PjW
mGu5XdMorn4GExW/AGQ2ZeK/WAMQR4OvODUINqeSWYZ/drAYNu4MA3UFN+rhUoF7eRMFW9tFiIEG
OODEoVj8ceEn7zrNEEPKUBOWA1drjEjUVOoh+p2ZrHInH4lnPqP7GbCf55VS5ntPPefDDh7ity3S
Gmxpblt2/dcTYXepJfJmnNvjS49X7qEhMVp0Yg8YzOUccRWha3VanYb6Jr7UEB+wehNFEc8Pk8Sx
6dRn8VoJ3wrppy1RquQQg09zyn2pdktWJTNWH4PZd2qSysSUSfEtJ1KuNxX7SC1hIzl6lJq5qEOP
3/+1XPvBsM7RwJyw/E543JWI5F8ozr5MaE6DUg02b0R5FcvwUWCXxbHz6Zgf4jCrfT8L8Ncfe/yT
0UtXlTeGPjY5yqA5ecEXfxkJUdI0mE4PaW0xZhDlsbk8VSLmLHdVbQDYZ1EBHOXjE7Yq9EFuAS16
IVTpq5qpOJkTG7PGNevGKM7qvOi0zupkH6djPbP3yp7EG22oTAliwCMAvT6lTOKEoFDzhDyFNGWe
/k+b22FK8ym2EVWhapGThuv6r+SifZWyfv7BEiK6u31fJUOVl/65Fv+fYWZtcnLXHB50L1E7pNsF
EZZZv4S0dQE1DRR6awHN4NCmFdc0YNJP/fDILihWGUTTo96vyuGwXykZ3a9NBnUsza5UCggrepcT
QhNRBJm+2EyEKE9A6pRoRgSSniKEqR2x3lvjn8XnqK1IorB887ql7wPOS+bsVZdCZPoiuTtVZ7xk
RKWhsX9XBPz6ncNFUxtEHTcn3TaogE9MCwKU98A4cyn90k7OMdao28oW63vvOEOKKetzYriSEwRu
5G0CNoCHs9lOBKUvrjpGq/5KXClOJE7PV/utUOQv3bSWFfn/2nXlx304z10gxEykKNiXRjIG+YbT
ZSXbwVyw2Yf/zXsIBisi9ktbMBRAfX1FBPOKyFF2UpXTIrT4CNDRUjQZBXD3WkSqE7EsKX7H84ia
BfU72mu+vqdUMqlPC4TCorrRizwo1aI7tKikWiuWxs6uSXAGZrAwgJIhZy+qn4A68yXNbDDnaJHl
AuPM+ElDi4+Dl4F2EwMbpnl+k6W8Byq4Rhm95DF/+gfkNOgirU2BFtOn47feubRHdpsniRO5OLSr
xYOdZG5lV7kHhSZX+irjobn0sK+1XfZKOVx1ZUtWjdmMTQk+2jJoBswyfzt52OG7e0XRGtHvUXWx
NehbJxTkQaXlS7dmh5YtxFBS5Wk+7S5gaCvJXrMYyjnNLgc0vyS9UW0LhEqKWu62MmMjmHnbuhCp
lVUTCXSju71AGJ8Zmw05p9hqUnS5sXsulCHOmKlV7KyRqMPkRw2/R0HcomFCG5kVf4mjvz7QAx/K
EJcsZ8p/SJf0A/HTQkbJlsCWf2UUv5EiRfE3nmBpE2SxhoUcVf7SPBjag3+xWqzkI4PSQEPj0BgI
0pnVRAe9Zps2x4mJ9Gx+rUsurwmFy6ZKqsLtbI5T6aRfkoAQcc4S1T1y8yz+65sQ0eoy1Y8gjiXZ
02tnVpEbyFevcK/c2FGplhijw8scis6K2cumLXu/pM/XdcBV2ItsYk2m/U3/3dnvB1yVFHSOtfU9
27kfQwB/OegfCfeZpyrF6ZpOGje1XhS6ogSBjSOgqjCGBwgG2CIzgJ9P3X2DEQOHBrfJa3c+OACR
lcUU6/d4lEPiQIHr1SwDD8T1ngpnE9fItNanIjqzbUKBXtoGYuQGMTbIS5X6wyhh9KaTQRt5jGSp
33eah+4YE0c+D1pD/UqTpiZ6vBFRLPoi8Dr1tJqBkhlMfT/WX0JgMYS0AxK91ahwSFK/3h0D1F7c
T0T3vMDUxeAM5FvBZag1q73NnLiRlbb9VCry6Yotk9eB1o4hLRuQ/lVR0rLkL2Sbiu4r132Q4zJR
Ad6SptYfxCQopNi0pWWZKTJbJHiAAXyoZdpjjJ4/idNSiYFU+rnMRMXgJpYF8V3ObfgNUveMUERN
obQKprp9kcqTY6+ueRhNQ/ugPa57YthU4HivG8fOaKmzg480D0Mf71cfIMbJ8DpTN6uR3sv+lb7g
nCRRu+3myktyyKNk3dZCezDts2SjxcgfHqKeSQ+D2zHKrG097kVPOpx8bBXLYjVtBpeRFxO/v8tM
rD3LjtbtzmgfBEFTHTzc0SNoPPsLZ93vairy/gAgEvVB+bcHDVCsNO0DCYTaQt7t/IJP+efiRhll
KkRs7fDgcTE0Zdfi4qJyO8k+zIYViCik3hRAiEZsooRJJogUw053E7CmI9gsmF5P83YTAoA3OHyf
9IYBCa1B9IG+21/rLIMnHSRAYfKMr6FiKdiZgchKxt4pu5uY42tw+YhCe/KTnb5Lk+ss6uMshj2y
Nhzcr7hcEc+KWzVxtqhmgiJWhczralQfDB8R2HN8uaX2zfaBKi63j5JAC4gi5LilHjxjuKJFq/Cu
xn8ZDyvf45eWPrguEcOh+JksUx/drD0ZwPaxx/JgjH6lxSHml4L9elR2ikA7s7vMioSSFxCRohSB
Vl931ET7SjUWd5xA86RGMKxdfJD2Lj/dtt0sNmlww+kw8isSgsorzR8FXtyOsJXiwL1W7Uju8/2/
x6iImEohPP5N/gg9D1/xJn3erOIPpOmSSCehXVYzs2koJTt0m09mr8JpmL0QXHEtfPgM741rcFo/
xyM8ODCbmC3txWpKCB1JEbwPSOzhkJblxuGwGbHPDTB5w+txoOz983G+QKg9azYpDAendlHBFuD7
ImhrRdVCITRm/flYM+iQvVbVKkIle6gltDAAIws3AQTd4Ia57yVkNPyd2/J9kLSGZE3LyUrHRwOB
kbj3R+6HtyEhRcWnz92B9VN6UfEPxcn/8ByvNRN4t7FkNMEkWCkV3xUIHtHn4AnF2QWRocGoe2KK
4NGMEN1/4LHrbKgFniwh5lsa9BLc9po51vOU+0ou7KbYbNc6a8bJa8cCf+4/iUxiSX1M/49H+ZMX
KzwlHaH7n/3FXValYrlD88ahTc+frOLMeY/pQXu0DdXjAeHCCIZv1ev37Ke5wu49bvfl59yJDhqA
g15BPAuxB0vUKSUIwZzW/X7SfACrYJMkK/Sb+G5N8kX8iP7mhAw2IAdy5ThYIZC9HIJg1jh0EpTJ
6qUfptzMQYCJiZvP5VbU0Y8KtsyB4bl07I9sZZxbg0xc5OXZ35oc2uLu/nCCY+auEOleqLP/mxKb
CkyKGcBSueeKbzHWVxDHrkXL/e7BK0pQ2Aho3Uw5M6IFEY8o4jnV3ij5ae8xkrM4XlAX2/GdJDZs
L4zTHUsgTJ8MIuXPmwPNq6Ky5VicM1mUQj+FNjk8yHWV9U5AtwKgK16OM0xnKNgbAF2xdv3Xsz31
I1DyqVvQafw8uG6KwH7bFFNiRWq2uw9xsKSftoRxuoCnq33mqidf0H3gRl99jGP9mVf71p4fVrZV
fDstzYvpe33+PFB+uo4kJ0Ezr/E0ZtHwQeQu627YDmNGa5Mk8+imre0c7vp3ztZ/N90BtNROucJC
6Mm1gT7VxxOou3jse32BNpowGa0wiNEUnrotwnAiY/4G32+jrWYa5y3ACqarXw+w/93OESy/nREr
Pborm+9F4V1+xmeT5maTVB91/WlokD38/vxW9Fmq2cl0uEHd60Y2RZDjSb7Pl2KIoA3THFY4NCaN
YkJVx+2tMk/ZsYjpxNfWePpa+lJrPGKbQgeKdkbrMCTnYypULRPXqqoGqmpNlrD+GGs8jKY1Gn8Y
uKa7oY3KogPVdbDgQLbCck7K6GP5AsD+EPG9Om5/UjlvAG3HE3UVM0LjvCLkjxLEKB7OjCpJo6PE
3sjug30dta3G4l+intJsOB/Nu/TBSUwqcDATFZiZBoK0SqfQCqR794orvH8wEGKsKdNkvrUdYvjt
fPPXJSK8q1Z0IAhfm6C4vzkeDBDqrWEqO0pySM8CqGMonTeyrtQnbIwcWNGByWKnsSORJVIyKtPE
WgCcH32ARlBO79wzZ+9TcWFJ2J6EtMa5kUrS3gBhUXJYmIcjOBXmKDnYKAhO2uMb5I/xPrjfGQKK
uKM1SnO8povcErfusxi9WqicwSr6K0ldcaj2BjTKKhL4kTMn07laYlexmQ8f3aNsyvf5HLe8ihZn
RR7ZzYHMMmI7/d5qn2MlqZWu8knVg+jGJuiZ3H9BbpwJ82tj/zu6b4Jt28X+oxsFQCk2x6Srb/dD
i/4KqDn/x0VGROsgHyiBCKlOHlAo3vwH1Pq1kgipz+F6nx6a7FYVsQG9sacGYhG4Q41fSiO1rKGs
liHmNp2anqvIffvCBjNmx+vrstpoLpSLxDHL0vEAm0cywbFOAvYKjeldce3lPCFntLemV+xCtkDS
3JxWfaGRMG9IPJJbIASqECmInPPEI3noZdKfQOXnQJ3OusPob/Li3o58hIqqAtaSZm2D07mA26wk
y4C6mZurEX7adiEhSN/eFnV/Aqo2RV9ZAvkAVV67hFF6cE4ocCn0MTLxwLAqULLQAFnqEkORdvuI
EdYmCWZoYgPZMjjss5OC4SVDvVJIywkJIYWxmrC4KTrMCfPJilB6Qn7T3Tk7SNCHDA+KXgfBVpNw
DGIgncxMU6Wnf135al9T/DQRa1eaZ8qHdPHadjD9XmTdvXsIUXG1Ov7uXY5dR2FiR3LvazEttKgl
Ypn9dTBy/PTuFDzc+6S2eoaugBG+iFg4tbFfw30kKgEMPXiuenyH9gwJnhXpT1gavmXHUfziK+PZ
paZIUMjGMoAh9XQrpmLoPRhpFJ/orwMnF7xzQuZjJODD6m+jp6oEbzvWDNHvnw/4j1Dhog7mi86f
vs9iBL9kdkxKzvAJeNvK5AhD7e6NKoiiM6lfHpatHbyQXQY/eNwL5HkP4OVKTn/V4NidfPmeSQMz
73E9Dkd1n651WANrkzTJJWf19i6oPdz7qBGvaKcmbEcGt6oIlccLKpGm2qyept6w3jiky2MFR1Zh
z0v6AJ3g/In5maJ9bXU0lxlu5OdUmq81B9qOFEEYrpYFUSQ/S5Z6rIt5UQ/pT+h1hzdKy1iffTw5
zQYWjyWrQP6+79mGCDAv+AQBmwFYVwb9We9AwBv6g2XAYktu51pgZAOfeF2Oqo/EWGKv0ltvwNLB
5p2XLzMEpzwO//x0Xc9v6oDAiUMkzimTH8UX4WjNiZwD6ZjisCkmhIXew834j3VbosgNbWMHfmo8
rQLhm2iuCKwhCgXvmOb9hWiuvS3lllWDIvpHSrFBYPvv0l+nEBxFpqYLhNNbw1LxSdHzwEz8DdTy
K+f0/zpa/GqIXijhfek0wYGADLaPXrpm7mDXiY2Popx+kxfwS83zu09c0ckzxonlZ+FddcMFyj1o
X+ljIbncmlK3MHjqTQMtNF0nKaXQ1CcWKsOkfRR/KzN2qTGKxs++92hwGLQH7zTQ2E7xEhzMKqA5
u6IrcZCU4p8jITZe0mJyOl5zENHsENSQmWppwckZygMuoJgAG5a7d6mAdHMruNXksiiGMfclQeG2
lBn54AhM1i94CKJ1lfKQa0bbKZ9jLlvBl9IQqB7J4/YcDLXLL8kflorkRK6toYt/ZzGYZV7OfH52
pLQ8EMo5AeqEXxGMZz5XqMZP4/mZD4WHYmSPWhHlT6ht8jueNUjMnbhdIZuHy11efzjBn19Y/j/+
BXeb8fBPlRjYoriJH+N+gI44vCqRnmHxwrmCbq3engkIg5Sbv1chUzGt5JhcjyCa+5bwe16e0fjY
UVwItfsQ8K3kV9DcL6A/APbG7L/aNFIwKXFVM71US7z/EnhJGHsov2efIoKh0BSn9T+lZqXjv2ga
bsFzXxEoi5ZkNqCHU4hM0PsGWQQcHpvuWfI0WWZ6Fi693B8lJ4waA/SZCtmLWfeS179nytIDi17d
8GxpdNMZLykmJB0E4JOACjtbpFBzFsMWs7AjCrKa4pRc23KL9yb0qN2AL2yNIoflsrUiEuoyPMe1
zJK12FcfdALS57wJqhAOV1UbEvXYY+9QZ2eDPk1OUp0QaBrLJiS9vPeczsI7xlMZLOlP877abad2
9dqUplszVCNPhkKWAf5TX+OVLDI1Ewk1w0I2ezQjXDcwO0QtR1d1fcVaEYf/XgmcCCHG2Kea/7su
wM7a36fGqAinOtq1o92dBMx4mtpCLwojq0nPfmVwYFhQNtp1dtPT2wg/ic1QshgeQfEXMna+JFw9
aCD9BrZvny5c5Wg8hgd/LtP4f5UTXhrlxmNT7H2QUJh2G2c3vXTGgIUHh2zWEJXvvllO+FYwtbTi
XGoTsZNTmgs55WR2btnQo6mQXJ0yFdlTusfmVR1NIOEIhLck/brq52p3Vs0tFgdEjw1UCzsm1vW4
0bmJtvBP4JypezPCNeewvUJrTtW0YddICgCiWKqGmoaqwzWwqCE1LQuNlV6gVcvrnOE3bZipDRnW
d53AyesVZg5sLjBrfGg1aUW2Gr3+s+weYrk+q7/1qOPn3uWeKIHcWpv5/K0GZsxDVNfnNWHA03is
Q0faY+uKbMFlv7D6p8LZaCL4UXYkFrOxA7tL8UhJoRSCRXs4lDRIWeo6+B6i8OmOEEmSeqB3//ob
fWGGxB6JD2RY65kidmJdpKYYPEAjB1jZ6Uz5NcFlxajcPbdXjYjjHlH7YHOruxflsL7DOgdLLg8x
QYpA0KvNULKKOF0ct8I+EI5XZtc6XRsK9PJ7wogzeT4eSbahnAbuXyg+aj2C5LezZ3QhS74emr/D
tOnUD1r8dhQZBa2yxWyZVBbjHM/0IibmsBf2dkInHUroOC71qPcb3cE+uZvKiDqzN7CJtnZLTN4I
1QkgySSP+OLGxLAuVGzQ0RBPeTzJk99lPzQ2VLPOYk61pkUbBoCSH/YlRYzWpgkF2RKtTWnJ3xSG
ZPDKqpw9fwp+inpX0xMz5GYRMWUu9rBxzXXdnvJolZLJ1r40ILZWDwPfN8OHdHdhGP+e8tpngE8a
kwO+LDyzsnaK0yNC6WexU9R4f64rQkRzHul0cPiDpMnWj+q8+84/hxoVr44xbDv7txrz4DslOudM
Lqg/VJrAVFTagTR0qDDjnK9cER7LXgA5I723YVjHN4HjZSBSG4vXeDfxB3xpgVV7Jgu/zqR47irG
Nxs4Gj8Beo4kosz6B9fxYBlYOWEEsMr6fBGw6QmVzJZShUw4SxBMNBuCZel98XpluWxz3Wn6rpiX
zXRnw3X066GvTEf1aYrH4uu67dyMkfF7T9V0Gy6BqsSNffDgbAAkZES6y96B8meLrwNOA+i3qlTL
O7mRcMvgFOATRKi6+8QL0/M8KGPaSclLiBa5U/N7imU1L8ax0bLrGzuDiMA1DgOPWUkyqwE1IR81
y0X9xA3DVxNQ/XBhNgOZeiPDKHW7WW/HXpue415/CZtkcovIMYdQbTTchn9XC9a79ZUlx9LgsDMs
sgQj2fNHZJ/LuFLfmqgQV/g2TdHA8BC3RGAFB7JtzX4lOFsawIjYkaSNNsliKFHvckjxBWwCz2xT
sgVwxctdenYPRcHELs10uEIzFXTCZO0sgbmv+YGguelxG2aE33oW9PLSjQjHmBG9XPqJOqGkFO4N
8OLPqfhROXEjgiKlqkOxIXqU820wkQROWV6u/BAzf0PUuLR/lgUec6MaxI//szceJjJ/bhzO/hoD
+sn1qzp9NOHSASeIFFJy51J/gNiZ20kym0gn4FDQ3Ta7yYVEYDp2cxDbwUIm5v9yXA2wIcjdmwKi
AmT/mnrnegADolnwWsBdPrjAj0AZco1xPNukkyo4azezBBPcIHeP+Zovy7NXNU0JEauLY2NmwkKp
RYJguvx+PnMMrj/zZCslD073gHe3ztNo/EmoAo4tT3ZNFAzyhFe9S9QQ91qg9ZazXsl/2/cdkAHV
WWOym0M5yLT3n3rT86B80/ph8bl2KrwmDsN3swUFkYH2+Gb/1bcVjlcZVy+Xo0l5MVsHN79NCO0T
OvfObVDdwfFKsuxVrSd6NEX9XIs77adSA3awbeHYBM8Lg2aTtDl12epatfivxfrUk1bmHyKZkfgy
ZFiBJYeygIRDzpIkZp7wqI8ebcG86aKJbMnwwdBZ+olrNo2IewVOFD4oQ0k02UkQ1vd+UJAYdl6V
izGORGu8abO0gewjLQ+TTDn4aXdXr6VvJIMRKivNTVEPRM6A6Qg9CwhBLXgxJyr3ff6YkZRiktDN
ijvfrsxjKrORrnITUM+d1RjumWM9a/OZQ0c3lBWzjZ2O7nQ9XuwCgHrJieKlzXslusfb3aZYn4ab
gaJJiqTdVok4wA6lzFFK8Nzb71ekpKei4gau65y6wAEGnA3VB337but2YQL4XuZsuOGuk6oNydO9
xQgHpKiMc2PWsWIjy8W8AMCTvd2V4XjhG70dYyTMd7ACzI8rJU9bRl+tzbVnOv88tvMjTIwOtQcj
F7GKpzo85qt8ogwHlhDHVAu7G1J19GFm+4JKYc90aaLZspuI+szg7jdpSySgbOt2ydcM49wk4KQQ
vsqaKl84qa3zlsjBbAqiyssVbP0stMRlk/+hdzwWn5+y96rKLBIzboRMtj5F9Mxaj/9o7+3O9Qw4
MGXB0gS7hyqos/SGQmLuybcKh6XFHQKs/HYe8/thyzYCdS2nOJTwoGLvtPkzaEBnlg/PrbMvUI2a
Ck6qiaTCRU2GkBFxWZ2fP5rhruMkZywzHj4S5qNnoVdHGWxqnebVdu/EVwTocT83UsqQn5B0R5QL
xYIPkS1FE/EKtbwm+TqRFKjVqvi6o2g7XOtyJZ5ZtZLJqlatwwvQ5LZePwGUlPfRGdY8zRhhwMy+
4M3mZfzp/xlZsP+JJLDlewSOdO8QW8mjOAqJ/VfRNjVVx3R1rrS5qZY2ro89tjgDmWj4i9l6YsbN
JjlAtjKlChWBofw4bHvubnh0wOPwIQln9BKJCTAIThYzQVdeDxV5l/s3h7J13o+QbsCJusHEGcfY
bTqy0AdCXmwns5WGqOqyDNlmllP+Yasw3CtNqr0uY0IvkfNogGbzd7dBRziq8aA1Mv0TGP5FLzu4
O3iEibXNdYjDqXyW4Zz/v1Tq0k7NHuRFiJmRbaJ0djGEEvmYSjZIiEMyb6QZo+KO0dtm+p0TWEge
hXYg9BUQ5g1OQG7U5AooYeTDMniNFIVBvWXjYCjyRMTHjouWqSLS/74f041QDXkvqe5kA9ZkZ6wk
n7sEUdcOv89nZxBI9meFGmlv02+ZPxrMSl2sM84+CDZcW2L1QIzDIgUWBjHDNKLfmFygd3v3jvkW
+6j5ZLYz9eWmdJ3tmcfrGUwusoEfzERpmGjVtwQ1M+zwdE8IvcYMPh9+VhnBJDsUz4i2hQrRt9e7
NhUQbvELhjDdyB5nxAPfTrmOudXFa/56KUgbBshEQdw1sMq/bWEF3SsLzdJooZzTc39iVJ0AXbHD
B4ZPjbg1tZlUVUBr9SOJL37L7vRNyymOywkRSIh0DEDhJUCLkV7Pc6/rj0ofjJtxvkHb7HS7Yw++
iBN4fnN7EMfqjU62th16GwUPzXWBImNDmSfky/QUuhzFcd2mP+rqvKd7ZwIUARp0sm/XB5oz9Msh
gbSZFZ8Ppk93wjmZ1qoxuHAeR40PblAsSoKrkmMzf1NLs1RhbAMAlckTDSrcMpX5Tj8oWAShr7PL
OcXoQAU5LLnzcVFysgJ2/DM1H9JqhfbN7ZALKmuf2i968tbqfHEnJ6LHtjZiZ/z2OTzWuqdfWpyX
Vw63MmzSI3QQb3WaO7zOm6uYrLQji+4zcdLnnatRdkolyXX+IywR6WPineXRFSF8G0IoPU1diWCb
iEbbWNR9bNGCi+0ZCx40tMTPPNemKit6qEIAGMrKqod/Rcn9RI4KMyeT8IguLkBZAK7kQQAkSfWr
m/Lnd51uuTPznzMXhSQMmAS2rvocEnSi9GM0XUl+MKG/1y6viNPLWF9FoKM3w1Ddz9EhMnCoAogz
YWZyxSqHy03Jx9aUvG7q5k8gC9zan8vKn6dGyi1TwQzkrj+dat4BrMyWQMtuXp4E5uAu5vP5zalc
dA2iAaBB2Nr7nEuZLKZuKATQEetGKwbGojjA+lwgcp4nftfEqzSznrq3U6QNL5DFMK1ge1eBAgK2
YgtYmznXOaFLLs8bHTZeHRikkjM67tkuUBX9qQhsWjiTMFiMUaRcqvsXkksFda6ZepruZw3QHz+l
sWnAijZ7CykO1t9OVByKrqFUINN47h5u6c28ZdK4YVBngtwdR6hrhukpr+TNrtBA4fAwakDkN7GO
4l6GfpMu3rDeefSjjoU1HAAMkSd1XNgCNmxo36HNfoeGh8jUK6PijFEv6AnP4K4f0VzwGWFWa9ez
HgI4eIVFvtQrxqhpiygfixrtiel+xMcst45rrzgwdhXB4Np9VK8BT0dm+G6VTdheNFauitn5H71C
S+uowY67ab8aL9Ch9is+l9OHw5wVbaG9jlAes0fzZRVJyaac3smTmx6GN/4NWd7WODbC+jm/m/HQ
IpQpAbG4T7ZJ+pZ+cLCYzRhLpyvVPTxnkfmEgqdkai23vB7aj1NirailIRDQa56dMox4P6K1Z1fs
Msc7xIPV04wRyqYGv72IoFm43VUDz4CVrjNAN4PhdYX2b+05+QnoGOI6eJl0mV1/6t/A9+O7Vufk
V3m1f3+3R9yPfATWXLCiINb3LDbv5LitDBzcpXPCyh6jNaCgICf9wZgBy9X1Gy3aTO/rnP2ma6NL
49/dCadOf0HGLnl/CTeixezGTNZFmYRBx/QeH950ceGxDlqXrCOgWJFYm3mv33sPrIYI0rSlt9K2
kAyapKBGgE9yYO/LAO5TH8187/8iuf5yhIrY7sAOay72POVrS0+HAiJFm0SV1FlmUMpmb1tKtx0S
hwqdqizgcUo/LFjs0yP7blH+jN945/zh4O676P23ykkYs3ynYpE0d3jLGKaUDhBosEzLs6BR4Avl
fqcv249F66J14mqU6YEuVURCQBWymiPeXVCe4SA1buPrVMhBoNB4UyAlti1zn1a+7oNHqoUzu74G
diuTmkbl+c/NUCxw1YY26Lr53nzctDpRwtgi3VQob9Bh7WtbJa1FKcT+i8ZESbtW69kp6/VKNLS3
bgwDKjRx7z3a1exENMKGmoG1WEJEyBLvYfXSzZ0d/5b/jsHcYZc1XwUS9mddMZwG0gNhteiQQIp0
TlIiAKiR+/lZJ9VTRV6A3FYj24ayx1KLZKxISDajPmH+P/23xIhHa+jRw4HqPJSroqPTMuO5Ir0F
gB8aFVFkf3AMZeG/1llwjsxIalbfP/WnKKhuPKVUS5vpmr1UL66VZ970mJNtJ6tEYEIrmKg6pc5j
V06ylN1iQZXzRW6T1AfFh042hMikCFQU+Cq+uxfDNnubzeEXI41zYYtqc31IkKnepYrNfDvyq8zF
QBLBLfjSMQnpywpXr5yvyeNkcExUkHYOV1hgOGLVPW+K0FRzypAem/7BThGOLcklz9gDwHNNi1Ki
lUsgekLxSP1SOGqcrtOS7T5O7GR79OAVc0uXfzh+cGExm8WmoxooQASYBnqUrGoNrysMpT/Dquzn
hU+wkNRk0LjocknoufU5csJTlSRSzwwQ0Oi0n/f4KKvvZdt6SAX4z/EEml2FCM6vJraXmz9ak3tP
QxY1i86oZ45QKRnDAvrNq+2cFlS0i7NADn/YDbHGFGkZRYqTmHMmC7s3xaspY6FUSaN9FyV/3kDk
5XIYd7J9kWr7UYjlB9o8RGGkgVltN/gc7ZcfaUutHe3fXaKzvfOD7to7O0sXMi90lOWZ0Iuou++O
QpztlTjg0NM2bE7qLGqs3tpp+6mXP35p4gVE31pEKBDqi8k7rQeaWvbpY6yylX5k8/3zr3odmeC5
8lnUUlU3t2q3r5IC5E8PgxRNHqeiSK6nOzCS++aTVhU8nLqtThRJFgZZPknpPpFtqiiSpVcBiewc
HHunPy91LdMVZkPeFjnhUn4yf93W2giq1XCqUJP+ag1kzDJ+hJjQJFbFssAv7Cg/xQEWLFNjapU+
zuOqS9S7yTZ5sF69rAOaBaHD+Qctv2ZtGBLFOekehwCFFCkiG7ZOYzZhpZyAymhBy2Vw2Hj60WR9
+P2Zb3CN8hvbMzNuFWfu6VdAyqS1OkptSTpanpJE2G8K89ieV1pnKUoBAIcZDfCuV35iw6RSrW1g
l8lQD9sX1lCRG9YH7o9GGEWSLR2Ph/Cg2pa6jhCKzbf8QHA+k88y1TIogpsqhMq91U3+S8Cjh29/
TYcldTEvB4TAcRXo3X1cYz/UoGXhHcm5rCglrTe4SgEJ5vwQ03BL9s6PAKXMQMkB/XE4EIrI66SL
5epk1+VDxZsQ1F2fuHzi9qgEJz1pPwNHLjV+9fGusgq+cEAlCYh6XxMGzGS2Ot1BnbNjO+tn/O6F
UJ4Gc+ZXfReTLkcyvIoRT+pUvWqUomi3ufCHrKpeqbx0lCcILyErqPV3y6CHB2ebDB6kRvhWK0Sa
5KTLhl4hp5q+slBiJpRLy3XyIdi6SA0/cmBEDDruHrjy7Qt19j4Mi9qg8HKgHeOSfDZ4VlRxO++R
q3tIXtzFBjVdtKIGXbulcvZpfApE6dX6fRn34pXZtHvfN+0bGd2rNgsgthyqHm88vRFBVZlndKXf
dAXDFoC0+H3krht556GKgzrMOwl7K7Pxv8nCZAP1/Z3GYmLrENFpBthxG7ImESl7a86HQXV5iZ7n
QVE1Tmhvr9GzW5tgoi/rFfsDTWfdIjar8sQb6HWMfWTYOG4jp1pSZ5DjUw+RGl3H332GJk1kxZr+
N9mgYyBqmq44CENiB7BbdvNFr5anmElYVZyCQe5uCLEtGb2z11BtqyAhro/W/fJ5EQiDj7NR8m4w
iE+71geWuB32SoSJbljeVHLWfVgo6T7kyNSbjhhEWwdesFO75mXMHT5/gvtsy1CC8T5TxhcpmUr0
JNlRa1U1hM7TQSoaj+gDiXuTTpRSoe/bhhkGHWiHTXLnvfpGlXYTfjrKcsinozx2v752CfQHwubK
c/j8b28/M3A/7PscPJXuH2+mLbBl/uMmc/0mA6ZA3bnn5mxwEFUrS0c9ZqDiLFqGXgZmdO4zosSL
k2JcncY9q/61m1QWNViclyxiT6patzGlAzT0x7KqBkBqkQvyhBLyVvvzqa1LlLOoVQVTwOD7rs/X
W73b/XJ7Zlj9qp2eSkZjEA2H45YAhsGX0BJFfjyoRZTLg3LXS83apUlxLNDaFP/MsW6VaOO6TztC
AW+60I25ooclQRK+gEMYsXnq/xyk7eHcbqWmQcXO97JdFzQX1q9Waf1MmelJFfN4/T5Aoqa84Q2/
VvMuMiXZ9nZhvERn9KVFT2khn2qsH7mOPq3JwBaJDNuQ4fC2uZTVaZJDZcXIPCV/xqfe7Eu+H7TW
+t/IsNok4R4AmT/Ae6xeYzrjRxRN6byjhl0eMKD1aDaR/1ukryeMlRVC5PVhtjDSbtdsy5blpdZN
4ov27nbTcT24B8oIonn7gnpkN3ZoPdkDaQAMO3IAUs772PIpnWQFb8ijHsndBDWr7ywZ/OnBvjXt
CWfIl3lZvtb6reN9c2mMS5VCh1HMPNYs08yj8fDoPvIxifHYr9C3Xc6aFTFK5WJOX5f5+q1u8c1f
NVoFsglvxvrJ72Qk6CmLSlNyzKHyfmBjw2rTnZ9O6IQ7thu0L+Fbjlmbmuc2Im6qwcdrkncQ7AvA
8IvDe1Owi2/M7VgDY3uOCB5oZW7wEaph9MqG7O1RAeaLPvxcsCzSOTyGRtzrDyS7pNJ2fczXCcps
pqS6VZvHu8vmvnaBzIAmoyAfxIF6i2W9ZBe11gLUrqnAvkyERy2bK1pPtV9anLTHdZFCNIDOn2p4
K0f0tTtpxWayCR7fP7vo8433s0uUWcTXM78k8137iRGfQetmoG94fGq8meevDRXQjsZuN6TPkdFb
kco2PjPY7c+tHGAa4Yeydq27iN64o48v0le9D2OMGnhv90fnJEnMmBvb854+3iHjoNmSGzjBlILx
OFMdpOBwwDnGUFVh/jNFfqGe6sR9tByG3zKpO2q5R3dPAWba4eFhaVrvJKavbjSvKSbqpks3PD5B
2IlYTyEUZ2k8Iiua1Vv4be6DhpWmYQQls+GUSuV1GdSb4XcAK/ltLkepWVkpCsw5/xtP10hoTuZt
NzA1bcjmykbvDnCbhRlHC91Bii3knOIonyTWJkgUFDcDY4Sj4ezFjDDeFz8A1F6Cz5MePtMs5QiD
XDB2qkdXY6zWl1XcUGO8ogXMZ4UYH9Jwjbzz/pRaTwh9JF1yHeFTuH73MmvNUqun923v2ymPCznn
e9PyDGR/z+EUqPiAdsTg90ANQr6YCiQ3Wheea1kWFYRDMLEZfwtqnXMjjn33geXYM/7budihvdtT
ng3KKe40SWzDs/xCfNp99EPOgIPmWQKudgeFs2/CW29oCcaZjDocxzv9ZzR958JfP+vwc69YPYBf
7wH8LI9Nlwzx+V3tVIfKQCvTQbBGdsfy8Lro/9utvRJOOyWsmniGjfp4NCkaD7liAYk2ALx5MuRZ
Qh1nqB+tX/lRB9hsBTQRkyRxwjRGNe6V1Fp5lLoQft9nGSCS9cXaexfLwbAdxoh8fU16xNWP4YnN
UJzoBdIdtODJtnsDUAZdi8ICMI6qQNN7FGVrB5ShnX8H7GaJKNemWfoaLnZVHtdhkUsQzIOZyamn
LKfGndGpVLO7QeOSbgePOo4Nuh2q1B2MLpffZ9Ds7YBp9UBKqiYNNSPQICN2xJ3vJln2QrB9q7Rm
NpMDrYOrS/QievdejCe2ITfjRSo76fWIOtrGO/aEigkK38zlO63yFLaEH0Y65pi0LezrmZWtZDdv
9EJe5pzSsli8Dk7BfCDHFKuNAqwPNoOXN1Uh6P2ZZcVuRaRSv8Y2uBRxhPWI/oObua9wV122GP1P
PWHTzCFJX/xZ3wFfBTFtbaYviRas8tKKTZx7ytVaNFAGiYLkyQVLRW7vY2Zmj569FOEKlMTs5a2J
deSSK9mNTO2/JdZZ2PtSZ1SRR2LarQmdpfbWegsYUpvvhLi0+4Z/q8Ysyu+riRP4IekYsQUHpukf
ixiKWX8vi8syd3mOlHzmeJ7rI2TcCzwH7IKp+Lha+GASjGNGrYZtgz9PBRxjF2OifN2wAO3kHxv2
w308rymorUMzAjOd3v0adOE4jg8clR8njA357wWAjopj2/uydD+Y8nd7Hr+G7CLy+uXkyCCg41c1
YUg8G35uXCcuGJAmRi4yvn4XHeaY7sUmnhStR2dPXDm2HlGZYA52pxZn1FoB7v9Im5Jzgydynl3n
RDh7Rhv7Tbu/rziA+RcjL9JBj/7cgcGAxP46SFsadaWzye6drW8WIyCvpBe1p85aJrJALZMPVmf6
6IL6RoXJC1chFI7mMyqTPblZeUs+euXB9yHGatFG1EWtbqTDux4m/fYOaFa9Rr8U6G9zcXwiOcyE
OsmYsqV8OrIudo5WHz5MBAxu33QtTKvVJ4cfHmlZlM9bAEPhCgNDjBhFNU4K7fffnfEU7G4D6lVW
WRbTIjP6SPs4NimG89iyDKanjMk39Ijs4+bLOxTARpmQqlGfDYRVPTgsddexL/qAfJEm/MPGZKIj
UkAXRojCFd1SWlpQm0sSimbMHyAUGTurpSRrnXjkjOrTg/+4TSW97h5Lvf1toafop+9FJ8+23U23
UqvdkuIEn9CdAEEZ0VY9zDGMS97RYO3a+YdVag99Bfkwvs+ZsLdWqdAZnf2qN3hGcc1M4YJ4v5T1
JLEJSeDgfYiAZuSzrob2slDI90y5swSyuygUn62JDBtqKD4Q0+eE05KGcZNR87ezg51KiqW7O267
rgTYXH75PaJf3hBl++ARiY1Yxg8F61nWYRwwKhRbq/z+siJpiPD6ZTm+CYV/l6Wc3u1tJBFjb5sv
u2NWgTv53DjaMM5CSdEPOkCJ/aUEmt6s4vWyRHM0W9vzL+kAbE6TO6gvFB8l9DPAreOuJamsWlle
1swFNiObFtmb8M0k8v+AiNi4O3bqDX5lZf09CiY6RALDqqBupRD7F1nN9ccbEELW9K312IRLxjEg
GtiQsJ+IuzdheOvdDTzM4NbkGUU90xfUipqz4C8dy+Mq2pHdwwXgynGF2qvGMQUOxRKWblxVpOqN
amBdH5tQUE1EgWRVcO6b53ghKmLbKsut0BD00x9oS3WCAuXXjySkSD/Ngrn2Z8rnBEE39TF/d6Rx
7a59kKBn431e6k11eP3pCI7Jt0szb27PsBaiVidMZsogkcqNzdv5/HsYmMcFkxa80aRwHiwZwE76
LYwBxEyhTXjV9begKgbKYwfuVI9FIAbqEcffDxngVNDIrV19nPCCxuiqUsA207X+aWwcXG3tKQ6J
1K+4aw7x+rFCzxjRIFpS0Hd7jn5QVUmInuBbCzWtaXuHUiwq3j9UIwpGLs8QFc1HkCFHBspbSyGv
tZZ1oxplD0Fq+zuA3Uomzo35CfL/jQc3LNyoGM2om9xGAwv0drmpaDVYmgv3mHrI5sHemavi0ymR
ES5pRFOE76Y7B3LfLC+EFfMQ8Kx4NduzCSheC2byMFbaQXHcfh3YwcSvxhv5K4hX1avtB2SGWMeU
OYcbPRchlAce1j/fQj4Xu9VDYBWJG5AbjPiz9ofHwcZnCjJBI7Q5C5lbNez0okN4g1C6g2Z754lj
vCkoK1XM8kgUlEpIyeStgVR+j9bNB4osbHgwFBk56qf0MCZLWu5jRHr8SkcreP180LxyVCn0IbcY
WTXZ34eN09C1PRSTcbpl71V9yOgMagkJ1vL4IaHF3P91+6sII//sCKQBstFh1JXcF0lDXVWYpVLK
9MNKSi3gbzMIGX3cIfXCiLXwYA1QzZZFu7AsLhLsHvVqOsoa/3V6PWdnU2vbbtL80Tux14bAU2Ft
NyWa639sWbOUmItoKDceszq2dWPCowjE9ZrOr9ZroVn3/QEZFOvNv5iqM1ks7k/WXIDfWKy/0kVQ
6yIpQ5C4I9gUWtGIWYDACxIIt64zNJqKoKgGRjUHxDxYrE7FpXBxEl3KubYl+xFluVAGqxNf6bvu
MNIWn9/dPDeU+rAfIb9FdUTpPXW0Uj63GJwdHHcK7n8rWP4h6fyhp1tJzxGcEsmCsFAJG663Yljq
E3ia5VzLNqQdg+LqjAXyuCbNpJaB58C21UpAzEFy8mlHC0qTk994wRb+uFsBLcATWb41skt38VYg
txKNCWqd6H77ftE946/tva5rnjVFHVDUJa/ZDSw4Uh92V11EXwYSd0eVoRPMqVHGomdm4MtXhxAf
l96e1su8h41z0DVtcmlRwWTZKH0CMZzKGIjen+Sw5P5/Wtqj5AlSqdvhDL2eLLSexu9OvjuFuzld
X7FtxmZKjsxxy7OhUMlwmA+4jJ0ojH2/ec8vwoYRvdyp26hkuAmRXcUs0omBdVV9OngPSz10t+c1
5E+ulgkEe4xNeHH9q+XKXka+WZ9+GxEFruMlS7+zXiqvfQ4zej6nnThs16o9gXYfN5B0PzBIAEwn
JgMlfCQmQKfHZ5hW6hvNp5CQ9cGtSPzxWAAWrxW/r1JsT9wwgc1/ExpOj3bsjHBNzCXknv1zn4VT
KXB6hjl1CsaO/s6O6f+SEoWsyaguPtJGALqfVpPuDmL/HygznYK2q+iJH05A9tmkVC3ooCZcxalF
YqeWEO3NnYpUKy98vN1xkTUbnJNJg32Qzqm0Vt/2JomJiSOVWpmMnj11IX8cTBJvwJv4CCrrhFVy
We+IUSefQEMKzOCvCNIqkwMlq/xzkLH6f2eMZLXOf+eHYVAvmuzolGA/dJCjG5sVoLm0rjdX0X4A
cJRAj4rTNTutoBCKNm/ev/MzCKGQdzErImHsSoAa29SE5nA7o9mt2m0fOddBDQQTlXWJOiRNOwHM
VL/YeiJPVO0UWDR5nyUGxGpkCcUAvcs18n9ZzF1D6I+Rr7rsm3uzPmuDdYTttRfEsmPRWp/gqLKG
mOveR293IKaVYyroRb6nQxrROpGhPxB/DFOdMhAwGEKcdr/T96OO+a30IS79w65TZNvHvyhcCEIs
FK/8i7miZJMXlC5Gpbvn4PZ62Tnsl5ZP7+VrfPK8efZ2m4AqFYfH/3yv7j3OkDxVGF9k2d4U6wzT
JaETKhJpFEuDKbtqLYJSKVLJDcQj7cRltNdC8v2d62m1tKYSU5/1/JJ2TYKlE+KVpUYBBU7ji3YP
BuLBOAT6tE5/1mi+xq4b+IpzcFSHVqXmg9ubXKgbI1/jLqD1hEii15y4Y486SYlDJYgIeu61ORkl
dG3epUjztXOwYraSAoWPJeqAkhZI01zs8HcsCpay+AYHaDF+yrF77NhVMB+w6+XZOVxE5bLQo3SH
KiE1A8xL0dSSzlKI19SpebpQNXnpKNvWP8VXG5Yt8hrqtZSh/v7b+ma0AKJUNX+2aO601BWM2/4Q
GIGFnRBal31btASPRDZk7pLBA4gw+odiyWUMYkHT126Nu5bqXvo7rfutpnzZGPSRKZSPHAYU+dNc
wdQYqrmSpoSj8JAQe8ieNGkpL447SlZyQQPKa9kH26X6/kZXWScDIcpdHQDNTXlo5cKH0X9Suad0
PNE5QMEZcMWvqapjLK8d4cMKU/fTQMOlV0JPGaz55pDmvyjX95FtdwuINsGoqvs8KTkj80bhGcFF
dPfZr7wAbNydIEBW4GWRoMKioh5JRTH7xlXTsz1VCL5Lg5cMhBqcPa/qP2VaOX+oIThLl3QuhL8O
iG1/4Oy2/z2/KoPSHl0XVwt8RIjP6fyp9RSpiVulRuVYIxSO8ExKSIuUDV2hFUPJBGevHZS25hNa
Hya1Hm9fYRWH0xxtjYSlykpPEvjPe3hzSJR23RDiEPaA2Gwo/4vn7O9iCpg5LPxWjrJ9xvLTkzGt
Hx+VFaScdvjLnCWYdvSAAj4sxIHOPME3KxMJoqnA1ZUnyo9nRfOv1mykUm2yGsNBV9vBTLXGQAes
JJTpOX5OS7tKFeKIw53yoDEKQmagC3Wcnw6ivAcJqUvZNAl/hxJCIADRFjH6MhE6sWMMpVJQFAt4
El3QZMA2LXCTVK+2PqLRgJgGzlyX1C8iTU35Ej0NFsugosx09XebrqOZ/1bQUnlEYGi8him11ZrZ
J7KEwo0W2wGQG2I9PyW6UDj+X4xtDgn4DhEFAkZGnnj7DPNnd1UNu8ayH3xPYFdFT7wYx8rUVakv
9K0r0WXrreXEhK6+qrQlFSEsD5Y9bdG6haEB2lGBfZCnhbSvLPsJin6OoBzAArZSzIpfXsii2c5w
3g7dxXvLDL76NE+15RBtEZW3ws5VM/XMHdxjdwKW8ygxcIQEz8Y+5W1aI+1QGnnRLQy7araqrl6+
nYcBYRRLyA6a9kZAUSPAJ3Bqh1x7u5Qs4mc4atQLJ2+ybedFu0+do5zFyYJ/5Uy11Is8+Z4EvOsS
6ZGltu9SroxcRbN58veTvoD/5TxCPZLz1TRuynM6AYJ3mFFzDrIqZvE8oPuut9ffrwPvy3TgoveL
w1FRy9JqvChJA9c5elwmEi9W+6j0DSrq6RFx+dSH6gzLdoGpOKfuSEnY2GtpCLzNJUweTPv7D96K
U09lnnYyy/YOW7vgc3KgZMUbB8Id/GqEosHkMYNIgAMLwrLCnxIlt9FkgUFr2HmWLBAcyyjJpcHi
qHMoi5pmHE2ssxnsC6BBXQQF69x6gXp4kF3QYUpSjRWp3ytPEtOWC6YyQjt8E/wpcOjdjyEft5RP
vjdkVs2WXVb9phiM11qAcfJPspMfhKEQ6Axqbr4LGQshtOLaQhdThu7rbNT3N1lJd/3dg6uf+MSz
nxUXQtPN8chhBZTckpBcYJqi7GX/FFRQcLoNZ67iJ5QV5OHTZTkwg5X3jvta9T0Cf5z/+p96EEDJ
vV1qq5pBUuLtejTK5JlaMh/sIUhgoh+Ee25FFAOBmHj5k+PQWSL48oVDdms1zL9EyalteJUXh98x
Lk3jp1WwxDR9kUF5FKSq97amJtTdD/u3wFV6+IzO+9KSN36wzNgSygM0g+HIRDHWaCVe2IA7pXYf
7o4i4b8F4nvvIEfYSJCXSEYo0xb7L6fXAHXUBn8oOylgjQ02A/tDR+mMqP0Go0HCbacj1+96TEyg
UPPWRzuVbDvA+jsfwMQPmn/IscIevpA7NNVv27gy4iuXXYpo0c2ZCv0a0ShEXBDCuvmDmhDkNL7Z
DDJVrCZERALxXqlLtPEPUt1z3T1ZAUQEyDTRPv9c4WyuBzzuJ+RS+Z3DH2g/OmEy/8uPs/b8VvDf
qeWyikOaKxzbcOkDy7fhV+40wbG1Rhji6hfaDfmbsd3idGx3gDkm6uiJA1vTQsWZqlsHqcoEMPbg
xLfMDd1Fs21XOtlg0VPQpkuAikEDndD6MEJRcAhKOKAsNxGUmcGgIwdI2wRQ3cGMWFm+3XCLWP6s
GS6OFv2GA8axnJz6mW56yXuvw5yNNC544Ru6UliEVzztSLWTUrfCWARecr0XV3VN0DpHx4FIqoGc
po/jUgpt81jiE04WVhSal0T1Js5DfoCzUMVDsEbdmFkdf710PM5Oat6cIXaSGQn4gX51TgP4rTFN
60isysQfw5XwqeicWS2m6eYIMKavxrzSmXL8qsK6z5w8tNU7lITBXgahMqsAT3fJB45SeSNaPLSp
QAtRkHmc01BBLDuAX4i4MPGq6EeCFhQUwrj6fstkNybSnTY8V90i7cm86xTuWlGaIsR6Qn5uJijQ
aUuHgQZUO3nrQ+6RjlZ7mlT0JAWF6q5hbKKklYxOF/wIjUWQ8SepUDZtPDX0V4k+/iYouE2b9qaO
W7Cl+truJzXR1iRfcHL8/Vl/cDchb0n7cl26jstds4IqvGv1mU0VjZqxOF9vz9VXxf5Byx6K2M9F
dK3FEBnkpkpJD+2blxxuUGDPLDa4SNoWak7utin9sl7EpabMAe2xVuOD/pdybzbjthz0adrVAdAG
Q13OoP3mS8CH12SWtGAYDWeRNu+0tBp+bb6ALo81boRIEVAl0HO2cnAsx9XVTlxifCpJfFAISkMB
Ow7EnjhyXqbs7XEGTngVAQGrSta8jW7G3tSBMdjW8A/vRTgVQKRs9uFNboV7Y3ZsVwP+ui1h6pfO
VChDVHiYBX7fNNE4nGpuqiKZaLZ6sMfV9DarWMK60QAys1AVUWp89dfMiwb0qvf6JGM6knC2NNMH
4/WVd6PMVhYlLh+w2QcO8VOEObdpPc/TCtuIRcIGGL2nR+jn4GRE9InYMXhYNVfOQQF1oE5DeKH6
iHvSvvvkIVwTjSVJA/35U0RXZPpPhGZcj+LhkBkfGNovn03pjO8d/dPFN6lP11xnt2SQMe7OabGS
tXu7cWEP3LRw0V3ikN7l8IAt5ZwDVVhTOyCT76e8OEfbeuk4pNaz5j1O2gG4XTwfq29XOZJJxtyJ
nRVmRIaTJ7f+Xri4TJeSvDdcjygrTm/mqc7Cp2Iixe3h9fJXA9sZi3C529Ht+T0kUHXdRzKOGZ2I
1EbLITUnVjIycYX09cBikX2hxBw9DWyDomMAaidEBwk7HNRFbOrVTPktpbDjR7U85S2gxBb9r9SC
MLf/kKlFdcVZI5zQTTS8G9xz4oZ+gCjT2HnThcpAFdiWnpj+WbY+0DJ/zccKp0gX34XoTDckg5F4
QaFOmdanvSqii60Ar+gJDVx1lv7mOe2OzbZGR8Kz/z1kS6lhIrrr98z/vH4aWIta/vkUa/228zPl
/NYBM9zHZkpwgDZ69FOoIMEDsjh2c6PUp0LjOFw08ubFgt/e+4hzfxay7LU+7UiR0u7z41BNhqxe
8ie6Egj45j2DMZ+/VkrVmePvwBHFzsDD2bJU99h9VvQy90CdzGnObi/9yMPPbzwtpRWVBTKbdOli
WXeHYu4A0kF3AjnwMboguuY2IhKa/B4vIGFCfETmyxOseq7NysrGzw9sBs2RTuLkkP4qNLCsScnV
iIXEDsVHNad2/wUEWohtZkIYNry5Edu/R+t1W8pQ+OUltJwfWkbwFPfO3Fk464uGJXcsxgRx6ypN
NSNNM+uKvOr9RMI596aJ98riRds0pW+uTP7Q7qQKNoaB+qskz3MJeXIYhx4q+Lb7kTf8OHnvRn7t
rjJMpJe3ksbnCI8+AN+avNmdSmFDFt3ZqhftVCqMjvXzrM48vlk+9oguJvv+ohl5W+uxSdi0Jcdx
7/GDq3UmoRZgOJGbQwFrU3+tI7VJspQprsBIJSBtWgCVHCVQ8+8hCDEvGHuLb7sC8v80Nbtuqe9t
mZ3D+xI+vWFzvqdrjx8QCECmpLMSKf8HmhZYoHcljsxAZva4JyAz35k2qGNSLo2oczWgL5RogHWE
b5i4KyyIbQFT58V3sh7BcJ6K63c5QDYHVbC9GgI15VDJEaLLfUS9a9ziyuLK9MwnzYm2faj5AztZ
vilFCYNeWbGcrrvJeKWJgYEwv1nLZWXYgIHQnHarhjBLj3w5VTignHGR9VoVOCAgk9N9c7182Xp/
7fXeuEnAVixNxRSkGxMxqxnpnpoZp9fj4AbCKt+l/O+8Q9k0Tjil86FGpI/98LeoM6IiNA/ytVrl
FTY0Ua9e5FyMzNkY49vrJwB5j0WHW08uo2T/YFaOrLj9/zJ1dNCemNOBuhJcH+9VJuuAHTWKFc6M
xF86ChXNyZB/oBE0Da9IO3v80LP/85Cjbf2kkp8hFLDsLAAr1fdHRYoeLE90KxtospRWMq8oe+C4
vqefQ0gHV6Dr2GN7TXPZs9Nmo2vXspM9k9QNp7u7jQDG+zVYsxcw+RO7/scMfzd9N/XDhxwZLUhH
v3l0ep9AxcqlVgkCKfXn33itj0yf8chkT3etBYon5PsECSjH922t+gcsuTLluldMLyE/WwnrjARs
vFrX0TSDhAFmduZqt7SwZy4D07Z2Jyci5WCahSs07lfJFOI1okr3edcf6K7v32rR4dRd8RPwRGr5
Obm7Xo5jpLY0FgZwQhRQtTXyvJ3V9QtukPczAfDP0qYAdUcK4nzQnrX42DtxZ61nr2uHAZTidZp/
A/ive/gBrtxMP0xoSXewgWxNr/JlLn/1pABnomVkLAXasqbLXaaOgD6jp7PwHYDrZeyiJrqojJ7M
q8okUKS9rdpwTSX7X5Wx2dkd7v7qEKdlXcoJnnXUl0rPxAyLFv1LymIFgiukck7JR7updbyrnBJx
vHLM0TBG2Q+nuwOzVFDKOpxxDHWlrXQ5uV8Q5d/hUw/1V1tXuz3MbF2c0dchS/KGUdBO9a9dxU3s
9yAs8DQCEh0C8M8ztbqTSF8nSBixEjvFnWIZlJjvCiYBi0rSThuXrMlOQKbsdmSwrLCc0NiPk4bs
d5hxsURBOBMitu1FcdoUXQJNJeCIcyD65G6O3s4pmXgyKOv6NoXOx1Wbd87CZPbugj2uPwDazZE1
aJ7VVxKWd1x2BzMilijLKTwElO8mJGAYtGvzXx6lBEOi6PvwP2AwT08WmFlef17i/n1729IWPgG7
PK6DN9MFCpaDy624VjEsu6MJDicxrFQ+QkbUYUz+0YbTx29gqU9ODzFLcMozgc1OgLqakmJIUmWg
+b//kR89Uo4YgMZUF4tdV2PK5ciusxlH1Fr0xFoY1ML90l2vMgaZFASIiIY80AKxjZXKIafq5Uiq
9OWQIuJ3CSPc1c5VejMxNVu0UrY9kxKkI9vaGTZHN8NH3u0p5u/OKni/ka0JwBC4/ysOYknFG1OY
wlPVVidKMOJzEQSLUIEM3gzj1boHDg9KbtS4MJGO4wdDx/fUR0CgyvDjkXAHGeK9XDZcH/p+xAnd
HwLhg1FwuQ1xGYxsLQp9pJOzg3kMx7X3N5Dx62I+8vc8glXloqUDDEmmLx8DFzTwKiF1XPrB19/K
u7TDcqjBZsOkARcmDAddTF12KuxRIkpvM5qtZnaep/ooLq/xkttu3aVMCSNK9m5dR4kUo3NC6evh
0pDbT5yCKKhIdJCfYh+R1ueYPW1ejSbce0CM2H3fbM828MKDenVNYeZF+k0wCh4iP/Pq28wIwjwh
JdfL24qU4UsPyUzC6WHxu71Q16LZWytx/Q8suAT/d51/1dFZ4Eid0QzyEpIKOORAOn5B6t47jIeb
Tmryxt7npwj3ZS4C20gEHL+O3eMAm7Xwsa/YtEm+MYxy6QS+GBgwEpW2A9FgVsbIyEE8ONQFuGSZ
w1FFerzyNtiFe0dxhoxQwdG01ctD1BmqrpKwoP8yzlEGuHpIQgGTlIhB4vKUJl3hgd0hN6xvcxRo
4BlY88TYEaVIeDkWNlf9g2GDBOkGxqsPXaCuuiqt5b8KSCk15w6gqX9Cm0vSVW/ULnmMVQX/BpUl
g2HuTZYu1ImzDTm9NYh0f7CvIO9xWlyVubGcUD61mlg3PhEehSKk/13+wjBvfsAYF3W6B9TC2rKK
vdPaPEuaSxp+0FEazU6NzhbYKzUDechYDyvv74ICfpnr4k5CfIUr/viwa5Fa4wRQr23ohuRBhELH
641YC9mpzyPKseP1yeWo0Arrm0O+BNQqzBLpUfvaVdgU+KOb67ccQ01j5ZVMuuUUrnJbWRyrIKVQ
wkp/Kz+RikzlLyXQMjBxjBO9pmCrboaOhtSP0KWCBh8bVO9RtHHROSpmydZID8AzzqU4aZAC13mE
7xyUwQesyXUgeBbgVToB4ivJOB+9dFMWBc4Rt1GEQiDibYhSyH6R8JL0zboU6RJyi4YAWirqkhnl
M+koetx5mJRcrIHddtsd1XVHGQQt6NJkRqtTdO7dEU7FM+y89bhRBNwbiUnX3PIft702yOcMtcRo
Sjxd97fLknXmtm7b/srnISTWg6+MKJPOgrW9UhNjwkwutjcqT9lSvI5Vs7h1FYAgCzspmfj5Qy6d
Vg6+2v1fos7FEi7+08D+LW7M/i0rCLnM3GrYOKlqP+hjigT9F95Uau+r+9OVlFnwLlsFsuk1qFbR
sy7WEMsuNY+LrL7xCP57RIrsSBrRxaZe68DdtaxqWY3EOQcfjWpf9KZtKDMPLY6ezYhj8fPLVndJ
SYdL65grv89WNtHn5XcyUCukzyf7gs3k7zUZDBbt+IxlpJmo0/edCWwyzaXZ1j933QPyc6t1ejvg
4Bi8aSFb2Uuhwv1AksPEBbGLa8RoQ1/EG5JXoYuf1jpA03CJ8/T/wZ8Vjo8TLQBsDoAl+/5YhLgo
smSsS+xKtoD+g2KooTteXM+l3xVC8J2I5fuhLLXi2cCHM2cFXJeTj3Dli7/aMmq1X44DMg01PqYk
ZQuCnYovycVK2QLWif5kd8Pqio8HXeLPlyiz1RH1hbqnL5UvT3uAC5GEj3yPLA9xoiyEcDIbNXU8
0yjngW24mTBlEqXQx6q6Ob35uTJg+5Mtu7y1o4y3Ngt7g59s9/JnRdALh0zFSIaKY8kJ/TF7P1Ai
GiAz6CaFzAdzBhqYvN9siFXR9Vkr89YJLkE0rqfatv1gxlGn9kMSn1eKCyGR7dWSAtGRgHnlKpxb
lnh+K8ErCAG26vH0RjITNEfA0j4NBiGvLn2ARvxiOxbNJtuIXQ83PvBqYVw5joYu8bEtUSMvdQEi
7CF2eQu2hPFNw+OqXq5F5Ez3VbX4C0i+huj6NwWjMNCfYgZWnMsjUwt+Un5VEW/GeLrdiPwp1Ydb
p+nnIuKu7EjrXGoOnBh+4KCWVfMiRyCq+E6OhXJV96rwLWWQMFvjtmInk34JGtpgRbRRAqewu2YR
uW+d4unmHIvAOi4uRVFU2WRVb+u85qq0nDXIawsKPJNRI0zBOkpQkDL6VJgWGEKRYjU4897sAeOO
HoKQaPy+yni8wLxlsEBI+eOTt/GeCDiiNqxU9C9GqoB9qbgOwvUujARZe2x5RG3oUWGRomhK1XUc
zUHWl2CFlVZZVo+hbjFS3jtP8stKICvdt1aTw+u+iivEWAkPWqwRm8jJfb6a3wDuCr9N/JoQjFH1
e6iBjDEI6NQYn7c+uTLgZnIr1VBO0cLC6Fdpe4bDB0RuEkFuS5rIqwWiJ0WUmeKBQnlEuLH2Fc98
gXUYAQJ/OJObuXtz3akHpqOu6UCn7CU+rhCVKfBYG5l4Ijo29FAzYNnJwJPicOQ4UtTbTgTZLNr8
BrqzSbpy22qnrvBMnPvcQ/KNXUwFiqF99gUjZw/JES3IwOMpfA2nhHK44ftQmocGOKJzKP7X4QtK
pRbQBYV0aClNjl1tUFAQQsK0XMl5VDex0p3dmUt/VjnVD17H2XyokehByn8urbpTE8EJCXPyQway
OCwQPepc6308bmOCq6kZXsdYe7YVzY7Wqupgdph8lRh62Vhepv3PhiD9JbwVRlbHpKOiQ9wIBFKe
wdAF56kW6/HLpKusKvShHmb1RAFP9nao88o6+alD1/35qwxZiD904iWujZRwrQd61mXx1HqLq+xQ
45O4NNlKtTm/ZoEVzwW7GHxD2EIgSYFs9rIK48XLtvUXvo3Mehjsc3KVtGI4Rz313Kqc/DiHhaHi
onBkg4X/yZAQx7XT7pTMoTOK3mwfDWfs1hHKxxQKgim28qcL0cca0475gVQ95fKcvdUoDU7jTgd3
826dQWkfITbSpTP+PONoPgefGsov8vXuqvmecfxVmHIrY+whtUAkBSeffFhwmpzu11CqaTrgQqjA
c31ReZObqg36UoGMwBZkzw241DTEeToHjac+of7mFLGqqZs9qSsaTyROMtrTcbeksVobnYDO5Vgd
3JTjL2X1XwyxXD0++0qz/khFZXxcJZhcr9NaEm8KO50CoiaP1wDpFi3D4NTPOdvv+gN+H5PXAMnn
gs7gE4D1ZWiYO/UCLWc6b0WL1UMiLTpqYR2ayAAwBj+7wWskROPT2F4tgDHO8mgGadFq+Q/wvZf/
rX0zj/KG8cWJnRkU3lEw/0rbao80Pm96SAW/1WND4vJTmcUGkWaPD2e5DPUTrqcGKaqZ+5cYo4z0
3NmiKXBudnTXiG0dRjdz41wB8IEvkdAE+7iks+Q2RCS1rY6qS/7tMqwCLKmuY7eW2cjwV7jXwZFg
pP3IeCxKjLom3WHkFnqVANKimmE5nr6y5e3KhcISfWf02bwAiNXi/IpyX2QiJGAiLb7IsQkD64uL
PBOAD5CfyoW27y2YT7gp6iUzFet8YMI1mPTIRrYLQM62D1siYIU5/caVSJcLvsluuIuMxNDTWnLf
QQjSdx/w7oXdAV4vlcyy2Y+Y3fkBlPuIeRIy/1O3dSfZHh9V6cpmry7G/xjiTH4ZbT3r+haehLbl
VB19QveyV3cce+SuLft+wfhNqgFYtU6HPeX94XVcgSAexF1qXygvhPhGctWsMzC4z+tZMFzsqBJp
lVq8Jv2219SqnkMRuMVbypFoj7VZ9fVt9eYxDNUfOhcE0ebPMwGxYASfTyv98h3Mmyuy9Vgs1fZB
G9KpAWRAG4vG/Dpkk/fHA4BqT0Bq/BnonW5Er6tCthefvvS98GRgkYiQX9sBsG2fcXFuhwJ+3J3g
1/dZ9tYqOtR67+jhQFJq3Uq2xqDA/NWwusy7vxEOXU/TDa9JjCXJ1USI41Jh2Y2SpyXOzm1w1Aks
4G2Ei/3xYavx7pDJ9OKp4QfmPsThbcd2AL/J3pfeeYQkE6wjPAYUTIPSrZkCLTa1zzMga+CTfOoa
fQBImGcJvU5awPJWDPb7UjKxgvT9uPfSmgcbtwUlBrx5X/0sw06Rt+6Q2g21PS2UKj7YLnkR3kh7
zPWMQ9bC4HSdt+hLKXj0wNqSBZGRXzZR4ChP+xntgilCfb0GOoV6a7cB4wy2aVpDDHmBazKaVARH
a+UTpxq7mvYl2o0jW6mo2a8AwuN53rwywGNvUtNdwm63JDi2H/XuJ5czzIOYZHYhvjMPdIVd+gNy
3YDwUQKZdRYPCgPu+03gf67xmQU0D7uoDk9vjiDb3/Ht1v3Ya2e+ZMwoFu3qS+2PvzNN/v34tr7a
mKV6iuiHw2I76qW1tYL/+M28aBY13Zksl/QY+lZKu4NdWchTDDendGrrr1cJo+PBl9z6hPtsfbjV
0Jlhh34CQyZe2LC/nKo7M+wVcrNv8K/l6+dOttLTgzv+aTE8qPIq6aUv3/aoPGLzY9UfECEds+w8
2AxS7yquDr+MfTio2VaI72IWbD2rdUfdewAKyRnDv0O/r6sD1XxIlrT9xRbEDQfO5O/O7JlVA5gl
z1hlRtHVH/hBKTxHmnwSY1ZshjNmrwfHK2LkAEhypSMLTwP+wLiRpp/NLlj7GoM+ZPRo5HHYVYrU
mz/Htyold0eGbwkhtWquRjvmx/wbzdbljqe7dW/oRX8h9hUNEqVS6wvTHyvcfX7zmywJT8oGE44m
EC1klt1teUUbKOtk/U6+HD+xX1M3cbDg6AYcmviWK0XfMERQNCi8nPftB9kdsuRZ6mGyfY6eOHZk
MqUEhdlqgnv7kBllc4To7Uz8S5tQIrY+Tlg43NLO3t9B64aaG9nSlt171uw+nB7y3/t5yT/l2eNj
hF86msFJlHfOjHTDD/ErHRWse7BP0Q3uRBVTCOZUFudnBls7inwPUYHrjHoZ7nknCbTHH8J1m8ZQ
jw7NjxpqD7oHWq3wYsupzIk+3lABbJ1kC1kRzIAQx0pqNIxE1clIQ71YJwluihQ3MpdM504Pc1/N
xqz7tks2Dscy4anMVN9T8rp7lOCINCYR5gmCzgUBQcEi++F7aUEkhf7lNK1UXwRqntp3fbyMhYJH
SbsjDbmoMXKBctitXuJ61a/XkqpLXSanPbgE8RqZTtpXHCw8ZpIV5NeBBMDk3dsNCcruhT/g+JF3
x7C7ymmiz46y8YSGVKIVQ7s61U+1ca/+6BnFa4ec0WkQ+VJERN0Aajz2lp0ER28p7hYaI/o8z9jn
5lOCuEQ50UEMjX2xOy5qco0rLTXnekxikdXCPetSVAmZLfmGDTM99ifKTNihEZ2RYg8l2YNPnnpZ
TNtiv2DcwGe+jM+csQ/SaUgc/jJYD4P2z/Up7YnaM6QvRREzay2mQVEJTNeQ8AZPHb4Ema6v8TUe
dAM7/0zhpTbSrwz8lblcaT2LWZ4fEQzQzL0Jkaa/U3xcxtrcl2gSsQh70k4IEFaFlMjzqx9g+oxm
ORokGeIHQ7riCHFQLmwU5YCJYQVcuZuzcUilVKZSvOCnEmQIHHUTC5RlCZUCj7znw6K+vrXstWu/
lL8qnSwRhpWK4/ECINqKbL8zsVSHQnncEZnFa2HrSvXSncix55EKy0mDWZKUJlPXQ0acBapR0Y03
y1PtarWZvG9jDI/Ry7u/2ipiUatIkQGIpCLf7Z2eYw2nRZ07q8sGbEklRpPlxoE4uwILoi0YSVvc
9pt5+Nooa2srmcLH4Pxgbhpk55d560xZZDwu/BIpdX6VdzNSozJ1C/Q8+pRvbDMjyCAeocJF6eIk
t5mQ/e1pQTNf61O/wSI+mRTvmtcvq3/a0hLVHbgJfOsrTVYOphclqjgw0eCSx+np3790nRkrHA0/
NTF30reW8MOyKHWAmy6RMXr2cTCQF296+Qc0frod+BdCBM/nxxZ2ccXQMKxERIopbgMiXVj05r61
bAyJ2Rc+NJeRZD2rE8qUniPmgWY7/wyYNs+xV8lQCnjZUz+fcwf8FZ0Xrps4cRrr2GinzrMbT50n
8hXkx3C2roZZlkcw4acjKIZkAhgK3uMuKqGzH94dDZdQOD5gZS5FMVlrY2RgPAx1osGvOmR4L8lE
kjFjVw/PgYG4PjPB9KF6ggndvBGQhVSkJKff7hLkykfZxFaF0hfDZygRLmDMMbE56C62BHiYWDbO
SEmhxp+b7L+UTYgrL9kn3ggZK1xBEmOcwsRkSxPWU/ne61yiCbH62+qNNEw/o7642TR/7kiQqawd
y20OviJNOD8UhRsP940OkPQcGAONVsF7eSHKA1hR2E7iVWLwO/yomao2XH1RTQF6WG4CfeKrE7WI
8nsUa072myQFSCUoN6QjIK//L2y6+A0jKWi5sa1NdEsTyIHWLr2EqVpmA71YPUwUBox59bRt2Cqv
RMKzMjFYWxsHo0+8kw5e54ZSaf6+AiGcV5BtEAqZoLYP5TXjd6pHp8/66wtGiiLQiy7G/dSy8eXE
NfMM8bGlmUh0Ms14wg2JDsa8RmY9VM1w8M34Le2t5KSZlU3bgzwN2pwN/oetjF8FxZTEnFJ+4ifp
ejjntwEQGGCHHXsxpgBlUU3cujD4YllIJYqtqVTsWftmSfwywfkKKISE5MYHikuQCMjTVzD6xSpx
NXnui8wW7MjqoCwZ1EzuquNDFq0Kd5lsgb1t5rhCyY/r8y0hpqWDfhoV2I/2uf8R4bhKX5+OobVD
kcPNnKb1AwsVT5WTXjXkVU0OQ1JTwVTOpfiYf11CC/zK7uFPlZp5Z4dKhAlljYoNQPUYXg53gtmL
HRTi+MZ+wsdAJ4y3zDy7Ywh0EZM/1lcCcAXcxn7NyowTto1+EqqsiR/gwCJCf4BbVIc9SbZT2o3A
cj6J6oEbBs76iONI21fCy1JpNlNzfFOuzJumwvPjKAU8/0mgrVmKWgipb+MTVGSkIMMHuqKE/rTR
RjE6ze3pr8Yz830qCpUfdsSjEXYmef/K/Sd3EkD+t3C9tYsa+DZBTKd7XNBf3dut4BGMRVOPNL1H
HZ0sORH3emeNnBABB/8owJQskQlWricYeA53qP89yRZmgi7+yYNZ+vufO82WgztgdN+3YcJNioS1
8VrYddCCLj4MIw3VWlmZu4P7KGeFc/tnmy8lJQ/oIqGZNwkf3iHOBSHSP8qtfkklurkR9njEB88n
vpEm/jRnB6F2Zui3ewZk7n/sNZnAZ5OskBQuKyFlumWHw5KqIaq4AKTT0rEX8CFaDHCpcj6BEjYQ
x3AVWwLCgxhuA1MDwNnY29xYo9C4jW02QmbmqRTop5NM5MxvvYkbeSQBKRRrmANn4TunvoAsyzK2
s6o/lwbnr5XbpwehrTrEOHXBhWo0RWFEnefQYmtKuNykfkZtxSaGMqcWJrLnrUcbaVwg8B9NkmFm
7pTHUSmwo0zPF6JwfDQUt1+XD+wilnlgqGrR+BqFiBW8/CeLQWYSvVJ3MyfDt2uTSSE135pjl2DD
TvI5+tsAQFlyhbqOiwkiAxhH6/5OUBV5E5AueqaEY90vuFeySjzU/yq4M0TRbCGcIJ0bvGdQ6mto
wbF9GDMFfuFoIbGMtdzbRD5SRoaDRj9JAVhHp8J/2ADi85QgHViEvQxpZZ+SSRgbXPMOvZqm9zgi
Bo1gyF9J1OK81wE/96YMwZBM3lnyBygYSmDlIh35qK0TlmKbhZpPWvslS0YhLHSdxj9Fznh4UYKc
L5GVCuAMon9+dAo0R25oEzee5NkVG06ehYtB7MaSIcXRxyFiKy4ZZAeSXDRBWs2N1DPrFcTuTKbk
ly+5FABpUkGvhdNsHQej47t/F6xSQCpxW9yk2aNsG4QenQ7OzEzgDNiRlCpelvl8wfgijSGw0yZs
5nP5VKMypLr5nXc57rapeYGKDWrGPLqhYT8AHdxu1HCkSaJSBu54k63VdBOm1P5YRbl1UQGBwGW7
3zelgZC1EgM9yspGSpRfAlq5IeuFZ7OsnjurERA5oDUqL1p+Lr1HL+m2ceaOUcx5ur+xVFqn+x2a
xYA39qoxW+4QU885iQcnCXfuzRyF+88WVLc4HsiBdrGOZuK4x05WAm/BYcCDvpUL4TkdzCt9hCfP
4cmahM7NHhi/S7gdpRkQMj4QNjFqyE3G2LFhN0WfbbS+BsdLq+M/DnRHzqPW8Eo1PozsqW+4VqHN
7/c0a+qA0r7lEcpTAYc0BykdwgjrjBDl6eoQKz4vkQaAE6yATSYDyUbhzpE6zs3/eZi7D0pBGQ+L
UNuqRVWKBhgNaJ1vuNQJie2Is7lbDA/PWV//5CP06IZkQzqZblZnReRdUAoYzzJM/jM0f25zvYTu
LYYslugiWc0OyDL/NZQJYVV1Md2F6iixUsSHFjjJ+3pDrBwcGvPSW2kYtikTpSVpbpHoYV5Im1yL
uGqlbaKHslGkG7/7A4jqDpqT4nTAsK/SCP/b3bb6BCYLfGLc+b+DKFQ8MXE5WJjLq/9GmY1EprER
KtzJkUXkieuvSigLdTOd7gRqY7wFoFND6wblc0On9rIXGZyCrAJ9hQf/yL0oGouu01ULvN2+sayp
FyvkjQzQ7LX9O+N3FAnV8Cdxfd4xEkSHk3P7evut5Va1mD4TbNZLVT0jFLGD4V09Yj72p43+YXZR
MT3cnUXAV4jeOyHMfjN2F3UjCYilUeumatMn7c2B+zRA+Vk6ZvwG22VQs3XZ0wNX2D9VvXXmcs/U
ny0gfIuYRb77X7lP6SIl5q3gTj9rHGILW5ET8GTk6a+fVxl+3z9ixtAO+LCJjGOc5mesZ9digIYv
ZyiPOWwEgf/yAa/ilc6hpVsCRlHThW5tSunpn2mTi6ePWs1e/sK2T32M1dRtN69mG2ES8jR4lD4u
lU10t5rVXj08rAscmu1zMAXVv9Y0lhQBYSsr5+UcoutWGsFR9/YtKaqZFitacetu+wfgTma8cM2g
g6DMojvVVoyODi660Mgw+CvFE7GaiqHxVYDSyyose2skJmzgn+MOTfYDeDGBmCKt2u59nz7tWfis
0wV5LSkDivhpnxgemAUoMisLQupoPx3VN94ZQdYmw3KBAKCGuI/EWywWa3mQXrjXO8GcVogGdYG+
KMdJhc6JDgsXuYneBeR0bECl1JdbUfF7dxyLBINojk/62+YIVs9sVccvcdRhvuC2ifjuPmE7tDAy
HSFue0Yud5u2n6NGwUMWyxSiPspnkC3OtF8beyEPCzRYmxp2zem8+iHEHsDNogZ9Fy55RaZMrULE
51sIowdj5VHJ1yCkxgwgyoa4zpKMeT1UifSA27ahrAfeMJlvz8zw0C0qekiVrpXx0+VO++G67cdU
UA9FIHNSobqJ0Jduhz1cJt7y+rBp+ZIfa/ajnYEprvmGEOG4Pyj9ecRw/HtcP6KaXL788dX92bNF
yJuGRTwxLxLxMmgd1ESQ8g7koKpwOQZ9ILbnn/1WlyZbnkWP7t+IYTRpRYXGryhgfceXZkC99Voy
q6g0CbIRm+DGxktBoOqemjDK+PWPv4/SL0ZvGWT3deISkVBmMzIqTYRvEfgUPogBckoYcbhbhw+4
1vXH/8cmUbprnrTfg17eRUSLOMkOtDPSgV9/54SiTiPx5aYyytYDPtUetP2GOClhhuElkZXUGLhv
Cxuvsci9XPQyM21WI0/Cd5648EuF/hC0VCNmLatOfByX4twurOKR1lIVdywzK8iVgzAMxZ4fvnwJ
2eNZ2vux82z+kdwvnVsd0gTBPR+0YTn0qbrXJO7Fk8Sl1oEmd6+J/szqsjUM7kLmuYEEU8uu6ZBl
IUqqbA6q7QvdBAFj8sxTC7dwrwEpsGtvlAocviFT0orLXb1OY/YuyVD3BzQ4H+Lk4HCcTl9BuyOg
ypj2d3bObOxsvj6xqId2PAKhqWlihxEwDDx0WcUaeZUCrQK8qHOLlymrZ2VDFFax9sBRY/x64HYx
7QMvfB4ld8OR/gIrWS/qQBVbn5NM7gjwmEfWS1tVDGqW8dbYwXkPTStzdR6Sy+bR+lJ2x3heYRg3
g4c+0/B62qfPf9mXxrX4r/cFUNHKu8R1GBig9bUhaFXfI/fS+0uXAQ3dp4eH+1z9fGBCI73B/2xZ
pXAhELqthBq5UiqCvGVzk+Zu9gupYuQQEcXUcBFU3HnExSHsHQozcLwk3qcfHJObSO5ZbdsRZxro
UyXefYdo/glTsSHhAg1UxKRHcLpdG0ZAMsDeDrCOe8lhuIAcrOnAn7XQLj/1155ynu/qIc8L27nI
ZqKysma9EGSE80iQ2DRMWCP/oh4vZjrWeTTcNJ2JWkDgSR6UoTEnnEMx2lrWMpn+jePCLVl2iiv+
AkCHsfiinc3ITn5JmXDIk//aWjoJTxDbuit7qqnYThrqmKpxNd1ZCMnA/8jbf12GY9XEwa638c0z
ITz7FWBbFc49xwVQXPrZ3ZULVfmMezd5v+PwIyhMRbvyigNN7DRJzXY3OvlLxQlWY2RmPtsBc8GN
gdsGPmwHbtOh0OFgqf2+4qh4ZeUu3EMpRtn91Pfdw8b5rlsIJUCaTrm3HuBgHemjQWf77AE8vuCd
pxdoVbjOm/ygMXonL6oGNDDRGb/XgQtukwXC48GWwZnDtbngApGMwXij6ybmGCQaPMFD/mHjLxk5
plcBgGP3QzJ4JpXcJpq0WgPXseUA4fuxEIjyPxRl7i5bJw4WrZW/98FOC5X6Z27Vn1zqIzxlw/ma
zNZsIJv9ouBSSQToG0C2C22hfMUlj9VUDabbrhdBFZgU5bHnB68mfel3wXIqP1hzKIK33ji7Zec7
Dz54bssgdZTCPjnUyABPSH3Rhgig2IdNVH1cj29g+kz6gPOb5W6FgsSblJGzw4l5jHZ1neXNpPun
n/PW2R5bzp6z/B24F7YKDIBNdV1D0dneryaYGgi3uPHhYGeQ4m1K0Z+uT4DgLItuH+cv0nJFPQAZ
hUn6omz5nlyUh51aM6O8VoPLSlB9+zCaTbaMrAI3t7MdzN2ObpiOnygO7CCubBfDmrCVhAERKKdA
AlUwOGcRuA6PAc54VVUjQAK6CCk2ojsHUClvqAt7ojKtOSL+F+5hjEFw1BaeFH76h7fRLi4MtjNa
JjmMbGt/BfUq8b8p9+EDCHcM3GG+oMPqItTWhdrIQqxcPHWvReT3r1zShPa/Wd3Z+MYMeSWt05Gf
ClLU3LutrB56krJYR60INjWplVXKxhalqXnic1CPZ0SoxQVSTv8ja/VWw4PNkV9KhvvfPhXVHJU4
c0iRFQwZBgM3+uTcMowBkTravVjnA/ZyMttlahk6hQz0CfVJc78Ycaocd47yBDAtoSIvnAwukV7j
OX9fh2/l1HgiRR/evf9j2r1RvBeCWFiE59xkgeiUD9Zt/7kUlXRRODieHEVbfZN7Bj1cEB68rDOX
sS0hCGQMzyMZvZLG2foTX+kBkcreBpO4bjFNB08ikRt2bUNutjH2tGGbMfk3Fx9fdNK+YRIWr/qO
/4I4vchpYEiKCvlTKyY/PA+Zbpmeot0y4q5w6+qx2Cqo1ROfRx6cPcnDcD87z44uWvG8jr4Ryk/e
LpRzKsP0x2HIrnbmDe1joj762CpehcSac5cZZAJm3f4HkEzzwqZJG2A8QointnGsxrtmwIUzHcwi
vKEwgsiFmA7BWJQiPgu+duoAre6db1iHBzZZtwVOVAQOXM3E8ynhv2ffrNrN6kaCkI1wSSKWL+fK
tBRO51lmOe3mbck2XrQeWZD43lcSD1IMBjgxv+JH5mhDF/sPqpcaQInM/w760qLBbJHIUZ/dSHMk
yIrKeF/E+mg/0jLyWs0Rv+gk1nRNdqpyGJt+nIxIa/6hDpFcdflwXfcSmV04sh5XYzeoJl+rcK//
5sl4ResUe3qSgexR4kYkHjVYSfauacF5nWcT/tcSUGE/L5z1KhCISOVZ/HnO+BjhNhK7dUnHS9JX
lirfYZ73W7GgTyTCXYelMgPzYlc2dp+UgQ8rmUCRjKjZqkiAp8TuEW4spaL49H+cw3iPbraAZ8uR
29tlhObgQOpOGyb/AbqSfi8ctmObwW45yEWABS5loFoz/wRQKg44h5sjzEvrohSbTdRPGCRz7m6U
b28Jr0KYlgvmD9Vt1FU03tBBgm7fMVCSDDONuzS0xO7ZWGTjNfFSPhU/ZD3pcc8JMB4hFOoseCQa
OKDdVaCIv8XDQbcLGdOFRZVPWey6bZJGkt8CAeyZhABhv/3Vt43ewBf2FUFf9iD7eyedJVx24B+q
l3nGOqp7Q1lr4VBHRFUqJmHwei9C6gVVR/0yxPg8MBsay2cnFkYkttxaiR/XWF1Y5bCj3v84d7WV
YsiEXCA8gJq+gcQXAHIAAicQYhlnFWsGwoaMIm5c1ac5a48vbqRqJfx9MVfGcEEGLGqA3aqqz0JX
01JQrcpbnG9UggFuLhZdA/qZuTY276Ta2lcXc4lC3ZkQmVYLTAjqhcNi82YSC79OmZF4ZpZtC58U
9uQvfBmijI2JrrhrDWVSPtVhxgOwfc9WylSv/c+h5EbNq0eJ7AqRsncTsXI5KLaeGGIaF909e0yL
twpz5zN4VBpKvvK8pouNtzqvbO1hB+S0PRJPX3hzdQYalFJaHZRR/6cGErFk3GHs2RcccBupgIzv
+bXfUW8HD2kUI3+xCoKo25Wx1CWBQlInZ5cRMtf3/MIPXu7yxk+rTDzuqyY2NgzrrV0Traf5LugW
Bqh1NY84ddqHp/OUu54RlQrFLyO9e8vrMuFiczOpmGWtfsaLyULwX3RtCBTbiwue80VrVx5fZgDw
U0j+rbob17wfyquAw+oDLG+m+Miutf5Z9rw0fPo3opqvMOMD8TuXaOm87M7orzI9YaplIbmPyLPC
L0jsT7SDwSgvMmMulJuon6wgJuJ8I2h9luUwYaRJbDxiqFWsG/5BqIQ4r1ep2s0lFvtXY+b4jfxG
4bhOj6CnlKOMATlh/itYNrT8gD0IkEMPOu/64391AscpqCx8lS01vaEuZ4uyKl+dR5Z0Xf1XmPsY
yNlx9sw6b6Yqiy8TAiiA8eUkWzVajWGuY5x6a6vjE9JMqf6Cn+U7varF/J3CkuMGqyDCjnMoi3V5
ECQi2+H2lr52jgan4EVaAfjN8mJmKlK6pzK5+1MukysrQ+0dCwkEPYjfcp/lxbAZbAIK1ThHhIuj
qgnsQfd0iU9LQQcs6OR74OwvzLR2K2SUUYuSr7WUZhm4DOFe9kooUspv0nG5abTg4pQEQBc0kizp
ErAoGViMseRG8MvLf8FQl/XXHMbXUGJPxySXRupNj6CyHc3NZBFg6vAUDaJBIIQF7s/OF4T2KV/k
4eH4xgGfBw+mzD8M7IeLmDiuInY0qbNfA26uJwj/leXf31IqMSTDeOUrxwc3ksL34aotVpmoft29
J1SufVgrcF6vmabiBv1lrxLNr5nYAct4yTixjSwShS/m8z1XNY5aDBXa2KVpoL4P1u+WLBGr8GHO
ne8JgIJyd2SwTBctZSEJ4Xbc67vpDhqIIAbdA3/REiw9o9SNO/7q8Srwh0JO+k0rC0dKhCqNWadD
3h8Pk7HIopKd1ydtBQvlRJ8zUNd+SZO+nqjeoZc6BPVk8FIcFfuoSeQsXJfKbwFal2Ir3JAS/jFB
RcBLKSEatp976EoP00RKkwUn6aPgz7zKBUEMIIjichjRsVdNDaPJJE3r1A8kIQZS1pT5rAWdEu0d
S8L+IdkgIUCvNhd5u2SCOng2+69ZuD9tNAAqqPWJIv4BgekeAzFIJr2bEBb5NV1eT2WLwz9tGdCb
uPrH0c7mIH0ywz4xrBjpB8JZxFrrN5xIu80yfBQQVd+w13Jh1VkHAg08g5jNr5c5XZa1hUdccgtC
kudbkMyCiRIpSsrVGCI6hOda8MBMb+iCaCMCaEOvV9jlqG9n3/LURV8IMnW9/lQ6TiRDTEmw2YSI
7RBEQD9OD1cPaIDoYN4cZm9mnFCphhDF7PEZUdtqamMoES1LAJoF1z7raQmj+zDW7nNKj9LPBigM
VwUVbotduWwz5Io2r8nYxsASm6ssyQ0xK9og9YDW2MTkGi0cjSNmNwma+AoEBeNeZznObifF6T+x
bMStvHAY03Jw7o3MfsojuCjwvUiw4aiZbfEqqDBE5YesjF4RATjhnX12r/DUs/sQhCmS7YaTmTI6
4TiE3qe96BGdwk8bdXiJA5DNNWv7PtvLFSFrix0RNpsr3FOiXTb/oIGf0qD5ATP+bqZCHMYMHQvu
O+ACQFmyguqLOB+Hq0Yw00QBI/jyATDfQD9ON0jVzXa3JoNpExLMNxkfh74fmgrPp6FLmNwVm0d6
hzF39EfxWdxJkJi1DVru+ujVP46Tn8PfiGxNILSj4iXvPxl5TGcyZKFMJ0BDvzC0YqIFKCHVAyMn
6CEHNzwRVdU3ZCSf/MdYT3keKKWhp1gOaK0X9JHY1nj2T373rnWQ1QzYqGGqnNluuZ/Y0hblhVbp
+XWa2MdjPA8v7JEFZW8i9/PH8B+5xE24yVHj2zMBHzxG0nS8eMKFyOgUG6HlE2EwNsWxJKV5DkFD
3O/srAsfqYHVWjykp+AXZEax+IXIuiTiYhsvTSQZd3WIhHFkL99guNQzsVEzPHs22u432+MSk4/5
cL61Tyt53MiQkF6JM0oT4SINc6zG/EvYOub1w0aIlOG7teKUb3VMo65P8vTuEZ7QLKfyc/EruOOD
Wo00AGt5uq6WSZjRmW1wz0FWwvrlQ3uEzG3GCUZhJIh04QGDgbhrqMeem5+yH5dhwR6a3/FwEAf9
FdNk0EWsuEAehFrjM+SUlFcWCSzRjzKFPQ0FqhoYoTkLCRUyJSdZ+TI7/wkfRuSnwn1odx/w6NXq
b5SqtLie8Fe23TxEOqLCKgsMhoq9ZoxtkP5UwLzmcmNSyhHWVjQGCVpzB5n2aAmtHHeTxf2yJ4HR
Fie02xlooIYjevgPyKryu0h+bEBKraoIh0aqdlQPzHLnUIedsXJAqZTlTjMDZtOKgIzPIFKOMHPo
RGGHi+qVakK7oKenJuxDEx+QzfFLPHLrZb4dBY3Y7l/z+Xs879cZAHfPR/O0Vpa4a5DC+9F8Pbi4
NF6sBjlhTyDSwUjLZqvtizbL6ePDDWfwxlwAeq0LqB9HKl9uwV88EovX4nMc3hUQ6qdOTgi09O10
22FvEGoV2PMJwW7qfW9BGfYQgnsPmF46VdalBm8x8q1g6xP4TbsMsWHNYubgc6UuU7r4sKJPWDmO
6n/MOirK8FotpTLQ9nvn3+yHbQkamL5lRAfWbdWsOuIrivN8Chl0KbsY4nlbNiy3W1W94uvXyqj4
O9Iwj/2CkPazdmq1KDzS9rAy461xM5GLjrYYMNc1/qvo5iz8y94CPvsT/fG9jJGtQpYP/jyGa2dd
ZMYpxRp33hhDDjYj7xfMD9X14dqBsRGHiYFLxh20IzH/spsxs7LBXXwTG8A7nXhNl2E04slEJ6jk
SbrhAd1LxBop6kbNpJdu3pqzIrotYgvsimTCqUswkjYQIT38vxM93cNywbI0W6VPjZp1iS835Iuo
zWc7ptmCaoyld4RSglzfAF9BSeB0MCrIi4zrkhQOQDCt/CTALvXiEUo9ZrVOxmOEloMGHIEkAPuv
umnzt4+AmfHz8zbk7rqVAoB9ooN2xLo6vjOSXQ2j7HcimCAYhIHcFGeMYHaYtZDgGfOgkqWNELSz
Fq7hwCfatte9PZLUXy+kjor4FITakztlOzvlKvjmITrTPPDyS6gzlWRmjnbStQzmlhzuPJlTLrIV
9S6ZHYrLIb33o/MXTuxof/UHj4upjGIHs1WpipDg9wU9+Hh4lH8BnUvKfmzo5/otJICi/YurCBAN
EZcpxSIVMp5fpG+EWXFxOxQHX0pVjCqTfkCszjMb55aLe92QGPleGRKYlLDny0vxmJdUl6kDe5rT
GP+KEPHhTBBt6I4FFaeOIDQSLsNDDSea2EHwQ6RPmlL+gJK/TOQzXYwHiAUY/wQ2oyxOHZLOtNiy
/RmediUi9HEOmOh3MjHdmhCJ2BeJB/l/dmuH1+QYL2163U0lBx8fbND53und5TQ+ffxU1TnhWala
jq8/o13oCN7lQe9K4DRucASd4VUX2ZSITUz0/pGaugDphm28s2MuuR7f2vbU/5rGUBjDv4iAZBdh
n8Kvj/+EGLca7lN4Lgz5G6MsJ/sulr1ztlUe9vw4iCWWOzHqeDqjWfYJX7AbjgUclzqPpeMk8yCM
3tlnqdmjQ6qJ8aal/SFjBdax6Sz7JGDzbiBhnIEXTceFhYmav1DnMSW89jZkMr3MhoScTj+z4iGe
38RlXtw9zR9Ssr51G0w7y+zk6Q1aMtQnx8G1uMj2bjZQQwuIndbBP1jVSrJ+Xp2NnRedvguKVqo4
lVJDj4sodSeHpi/K1VDryFdPmKIUKEBDhm/jMShotKznYHA0YE/K4ppMuDnXCCHx1HSmviD0iutn
1xJi8pYwhcZRLmfidwPZDOO+EG85zX8ZNdHj27np6cSG/77c5/ED0FHZm9hVaoKV6Ix5XBsqBMdQ
3XYIsJU+7k87aMxBYj79O0UVj1boYCnFmO3CW8pUzk3e4R24GaJF74tVnynTdzjY+I2CE1oENWlx
jwKmuMTjs4JtyhyK1k0wyIu7hBAF8EGPAOMyWuozVzUhygxSqzQKVXk9AGzybac3wv+Cg6xCJwKo
nd6bEciTjGdY07W64uWlUsLTSs/JfnUYyXsrhH0H22o4kPclMlATnkPuZp1w8j/aYWL8tRoAw88D
/bquU84L+ieFU7IhMShljivwoA31CRhiZ/am1Kjrp8IfgfAF9JIWrMeuIXkWuqZYEDF0xYBNLHZn
bhOggmN4e4LmXTCPm5ygTxK53fxrXZmxqLFN6n56p95eK9i4frCidPnuPd9cqHmqY8XBL90LbZvA
6EyIoN5RyJpc7BCiU61jP92FZ1YrEHJgu2I09QsLPzMpMbesvb1LT2e96q2/ra7OydfZaK635Fva
gvnTWseKHrXWoVOxzvOsdta8uFEdd6hT2W2pGdCgvMXppPZbtckKJYxk8aodPj6JT4uzK/59Bhwf
1hptnYNiekunvYXmQuQZJ9B4eRldjVBFie10rpvmsefazXvOLdPkU44qiCXbloF51iSPQBstujUQ
JVsb5cacbA9/EDxQ61pnk7kCZ8P91cSJneG7trPkDGKc2kHiRZOFNRGp0AgBXShBUAc6mCkN0XjZ
QG1IGrMvM7rpPBk1MD2YNPCwlE3tW4EQaCFGkRj6BxR7mtwFz/yR4w8GritWplsDHbQMlRzMnYEC
9NUTv9isk0HpB0F47ZCc+KD10tDD5Q7aYwyr8GF0H2UulBw9X/q7WYRGRqZwrrA6nGf37s190tWi
YRxE3uM5mbG0dBESM/OSjs8kehAoXn7Km7G7SViJ1a8bv+4eFd+RwFHFKnzIWBbBPj3wpvBcshPZ
8dS0laE3vShOKJ4XaU/cO9rjkPTyTP8fJUWwtdQsELV/Bib11WD8Dq/1JKJeStGKwR4zlvT5fYTO
5dCt6YH88FGbhJFxCKu+nEtOYzrSzIiKO7qwwYxJg36NSatB3WBMnJtwoWZw0WOq++lddlhQK2iY
QQD5IVktStfxjmle1Bh4LLUq+VAXa9FSoJbvDPFU7CklxHlkiKQ55CytjYobRkomVBYePJ/smwPk
08Xxqt4426NuaAos02wk0OQt0MA/esUiqo9kFpu254P9eSL4zQNsw3ttKqBkhrdiKD07Xz3B0pFb
O5Fd4JmjAblAt5Jp5Frp7B1VY95yOj59cdlwBxu6rRaUd5mYReJcCd59/AiZ4eBrsDWfDsLYjEoM
18ZhF1aggJi2FYkFKVFFMb0ydXYKvgf0mELFgRYkTzMMoAabvswPXX9Uf8EE4e/RbZQIUWaYBYLw
/aIs4HbWyJE+FOSk55jms1GTSQ4aek5oUI3XW8ttFdZKSVyiV7X7lwgtHqi9dLX0aaL2+HxoPbJI
dsMqL/V2SGJIOgI2dYVzx/R/Io3KmsjrFFGTzYwi2RxU7uhkCHD3iwudSdu5drFyVU8cKoe8VHyr
b5Y7ZlHYGvbscShQSWwrAKm9PqEgyfHReK6MGx62sGhLQ0j7PJnGJBsg2MWSnUZXQyvgULea4P+A
M6oA37xSCxsYIHUAXp/dQkW/ptayXAnEVvFKdmBooD+CcfZCN3BRWCJS+a3470BItr7C+jEJf4cT
taWRl/lDBjBg9O1QuLcVbQg8FAWNlEYp0YzxbLF6hHYiInoH4cI48ev9M5nA2SLUDo7qXkje4OdP
f4FTDwnTYoXPeu4UYpbEC3tyJnXWJrJUPy6fcZKWDhxQ934emynUPP55uregfnbT8Rxb9Yxl/qoi
gBJgb63ToXcMa/yqPBlqNgyuTsijM1SogeS6/wd484YDet/I9nRKI/njyDAFhgcXgGrK7PxIbrAD
b+E8VLabDC/XdtSumx54kSAfDzXkMwZUtN1aXOcRCIee50HIUxa9g2ks9whJyYmhmrxpVQR0Zrf1
wyZO7seIQY2R57jRSAkMCoa4ScSgujYa6aDCNUpMAD37vPNnqReW5acksaxpBNyR3enTnHjX4YpQ
iA9HRqhL/SpBQvl1ZyV3f579ifjwJJ2LRb+rpRucL1jvSDg1NW6Knr6WNBEGVibyBsMhamIx+nRz
7tqcKIstqcteiMe6v1lFx7fl3bgwhHU4Tx3c6h8PoWk/rpuUQ7VEaeWHAFinsFAVX/+jQWdawJx1
iRgnGhhN0ibHrmCWGCZSU2gdYHmqRCWcoMnWxZMSYe1OouRnxdrCEQV9bCj+9xV5fA9CzpIjjdVi
rBViKODyd8ipSa0ZDXNm4Z5jd+pE4IFr9Y5af1uWgOQ8ku4d9Q5apa5b0Ru5IWMVqfBlOC0BDeDh
lfiPFZ/dNRJDAcbtupHGQRy43EAmfVMUDm8i72T8k6/xYY1fF/+V8lAWLX+kU3mSAUJShW6MFIbR
SO5rBrMHCRtPrpVhYmyO6LE5bZ1A3kuLwv0zKsiLIdPXdjxTObCO6+8lgBbEj/b2R/53yZ17njhv
TfVXNFveuR41xGTeww2a3CylG4iKAlZK/xjs2Odwm6gAFc4Vir3bHsNuBCvwWaZ6hL9ZObOfz6VO
xsHatlijB/YgPSH+Pni4g2yGU4msEtWcHVb1Mh/80uOlOksIYjMFkoSa1LnjxZVy2jeGhcJhTHR9
3mYQw3IF6yJjJwm+NYy9YDohnwefvUZdU0gsy/iVGNIfj5kfm3xSkqr7Xbszpzj0hwUwP23wXBIi
6K/zt7INIc0h3k2RIH4qv/z/8ejUkY9pAdxshUpiMrO5SzkP4ztr8AHh3L+yJild12is+n3BaO8e
X+j8JK2wYp4gKBQc3t01r79wTHrGcECRUATP7hMLy6CYxj+Ub65miLPwhb5WTukiZUG3WCJUxJJZ
cmeCzuwe/Fnrf/zBQDYoIWch0fwnGFLRo112rEyhPkwLRJj/MKqMcOg7xqtPhTbTJ6k7IcsP91P/
1VzoO9ZXv/8HX/rvV7SmPaiBN7acwkN3enMyZDdhkY7Y7myi6sLva9E3+tJz7x9Xmgr0VfSSUX2D
7aIuWobcyGUM8wXJ7bd7I5MD9LolTZmhVgwXotLXXmH/cKVuVtw3rrK6ww+GSSWdf4Peo94in3I7
zR8heZAZ/WzmrfyJoFAjFqafaCDvLck5qbE4Am5D20Us2iOINQb/oJ0dfRgFKGbmMcJYgjoxvbjP
3SeTcH1sKTm0MJIfsj0YZWMjqG1DIPd70RIpnp5lMPMLpdyc8LhQEBNzkFTtUzH9hod/HeKu3v9M
1Ox0GS1l5e7yxa5y0sU47fd4EzZ3Ahk07cf1JgstkkmM2DYmbRcScAKk2RnBQekXE1T/NLxf/HUD
vb/t794HHMBXHXSaqgoPTAvDqHVYbc1VT14+k9STi/ye+jHpYYI5/tYnUQ8YQ9C5gFwsskpiCj43
kvXvIwoOPQsU6u1yu14AehLBe1LTgu3OGRICHYN0ryn62LBIRabu/tmeE2RLKAbWQI3Eqhf2vzWs
A274jWOYIb842IsP7HLRtnN/TVyqIXldZY/8GREfgRotxhdqQG9DuGkeKqbwEh7hdWGwQ3RC0Kpy
sStcQjOiNsiz7ViWEHJntRYrCJiNbjF3b4THbsHbvP4T/bFBgrMWh1TT0rMV/avkKT22I/OWQOG6
hRf4S3tAYGdwTw6JbSJMRsOBIShSuBVFT54KDE67zGYaSNLMBRNnQnKmOJ55Y4XFGqf+aAp3rQT+
wTfL2UY5iuzPvLrAvhz574L5djngt9cxGdrZmBhCkrmc4PIw+qfjP7UrIQbKv7id5Q7mY2ksjFpZ
AYq1lNMOFWDpyfP4lkN/xnMOJuW6c0x5VX92uCQHAb6J8RMNr8ZJgTLjmIiDcSkwdK1L/WVzmRRt
dvPZe6pX8A4WLxJIIrIz0jYHqVmwo//yr97bpfsjlGLmp1ZZ7Hy2JLMD5xITnMaNkGl9EIBpKvhy
u3VSdy5mAJzAFxYuuD+a6PlAPshAQ0kO6Rcw14XPy93wgZ/0IAZNgYVjkjBlzmhu6ivDIvua+vVs
ssvTqsFp7kDRFGruDPyMl65DXefY2yxiyxqSFS7kioy4kGIm+d8GQg+NhrcwaEiMS+7UV4H/tEWe
EAOz20uognfajCdyD7oS9s5sDevtS6weZ82/JIVjRTf8ZsMZlhHDB6Ye+tcgofeG0ELwc3i3dAIn
M0xqnJoGa6s5vGHuLbFYDubxutBWFtfwfmODOp8YqCYFMXx3CD+GTbH4vg8ItkoMZk/9czDByqz/
fFTjus1HVP5SDFLEkhymaRQoqLoJ2HRyNxs/ARKO5Z/ygqYucQBv1AaYQPK+Ypd+1x2igRhl4LTW
05HPqT4sgGQwAAztdfTHi+b8AQmf4/LbacEm32x0Skmkarbpb2wvEPD1bz8N2X/CF9qqvMl3B9Sg
u5GgRBTWyAJoYqqAf2kBdDuxAeQofia9lzzFhXVzacpRMhJpeX8VWpjP4it1wnuLbBqu7/mCK7Bx
UEkxJWj5Jy+HvdXytYs1xuNzXzcCUwzi9yyHI2LS4jbeLJ+m9RTUq2k/UbXe4AFAsZvTAEXtaxX/
n3oDEZTnOYEknBOdFpKskKlS6hLJHFjp8xdQwZNfi2IEPDyvKiJeYhMRUNoqRJA9kmP3rcoluXwt
QnNmJf5SfHOYrlUqylo/OQ45E8DLSNrIEx4dgIR+OTWaX5ByQZPWdevaNs5YvcXoQ9uCAE0toUHx
ct86jskPcCa7CO6lrBozOboHr/5qGgyCXnKWmFj8rpUnXT52CqfRQvFoBPiIgdXnWc3Wf9r3Pxjm
edHvHpUrJX0klPFlhWK3KhWHctd0g+8avy/n7/GthT5zJuBPqM/doM0AEZXnqSGVQa+PtQp3YK5y
f2wiYW3yZcGl8ZN3NF/O9/js8TQM3kIMWJp7hlJgDDFGZwKKoL+vLQUvcjUnRfATVwwC/PTceSce
Nt20YBJIaVa4PmJM0F2S2dQMaC9dkpEuHNtJUDXj0PHGv36qPMQMb4L0GHru6CCHm+IJUPof5mne
H8jTXWE0smqGrBWrxKjORK/xNJdjIkGs67Dq2KnB9ASvuszyJGElnEdcritjPhsGJHvDSLgahR0E
pap6MbpwAtcGbM9UFaLtat25T5wwV0foAY4HNGnDDsr26ovJq/f/4TVD4A+YmlgmGt+xTvnE4nhu
BRu4/RHwqNsmqqPWePnEygtugAlDIqTker5XhaaB3ZP0S9Y7FDVW8E6O2tS3gKsVgdlOE8/ZqaoK
/VlObm7AljsQrK+8kJABY0RDSTEkNGVe4lLpXqaDQ5jcYZbfYtFePnacyAxdiwpeDVqWXgC9ysmc
YpIyHXXlk3gopO3h4RAYHNA3k2s/CXqyTT7yUO3ohlRzF5HZ4eVc0nzBPEEv13xtA8rtuO1pjdWT
2r2D5eG5vG3iV9Z7sTk5LKlH52saZpaXCIQXCAFhkF1pPCjWB9OqroeiGRJj57Z+N+Dv/yXsdbW2
yGB67BYX7R/u28Ckl/lzq4EEGLphJr5OKmF93tcKcpprSAwqSOTdloXPfXtMkKX7RRPGY6FWp+4H
u2lJ6YqeOazs888Fs8CsfuPmWFFrKgsAeBQCxsgnkf4VhRc29Y70ZP7Y1GXHMM+Lnzib5Hr9fbPj
a6f7eXwhDu+HFqV8lvdTGXp3A0IX3dj/Lx8D/5wG7IkF9d05TZd+f8vMDIB/tfe/ZCwWCYPPzCA/
aub2FIXaw9Ahgm9rrZ3VYTdpKZUpbILvqZf8asud23uyB7zvcQr+dI8AGYnAZZGVxiOH/cruRMFf
uTHtw6lZ3vOH9OaGsPBKXm3bzwaVpw1nZjkgJZadp3zdrSxw4qsVkVkFKct7yrICbI/oCuwrYh6j
IRx8jnTWX7DxnPb4Atp8CtXGznrcSF33fIt7aT48vJnzqHcGUghC1kzn+T9ISS1rJc7MJdMuASSW
tDvQtjncXVgS06mlqDLknTQd6G3VAqusscSFdJZ4kxZxftXVVj0eC+TIxzSJfoEmCMoMFmiMANOm
SKaM8DlAyTgVBda0RFdozSW34/yM2uNHromdySqB9mIqiXOrSSghDLKxwwnXG5nzCZo/441GYPD5
XC96Q46atm95gcKm1OqJWohF5KypCsNnXWTiSWCp80oJGJ7BXhhA3DRRaUuttqdD3RF4zwkWPdlt
czOKUYU28y312afmBeqW8CJBPWQY8VUNBT/1ftvCWj+4/HLQR1s8J5SEzydybzyIQxU1bc7Rwhbs
eqxiwY9dDeCkU5UOp1rgHctMCa8HeTwPg82ZnPpf8MxvjNnYLWvugHbmFgWm8Jc9IzKISURFERgX
rafVRhEZwDZMrcm80zlIkq57Gfi0gz02RVa7ThbRpcp5gBlaojWtfiDESQDwRj/EX+VjlJYOJP5k
oZVp5LHCPrKR4PkNNZIShwTMA81YLgx0YW2dgs0ZCP9roROijqb/4yfqRNfyADbhmC5cZMmwl/dD
hmr22UDe+45kY5nBluUJuLnAYCL1tVRiegk8dpZ/rJ7ABLzH0K0w/xQYVEn9ntivFZS4K5d9ztji
iCBqefXN3WUS/Hi5dyst/mffhMeVATHHc4uO4ruWmuqa8bIP80CQszAousOyn04nasPMHiuVG50w
rr14IywlKzfXnNm1Nq4NABecjGEf+J9F+Xe+IGs4PjTIByvvg7oTkIGUg38mkXbhjmFNA9VmYdvE
VNxMj8255GBbaoOvARyD2Yf1r1wR5anjaVtHK69+4u4dAijR/Jt5JHHMwy1coUQQ1e+IojHa2HC5
dbs3624Uz3GRJX+xSZBnBkM78tn4qwe3p5sZw7z8ksXaXbHvj73VVQp3lVZpWy7/762+13m4bsil
b1Q0iYHF+5/tvEheYhaOSlUJqb2aW1+iAM6E2l3o7U9E2rUIc6Uh4Igh9FuIbCn7B/3gSo4Hv8Mf
W8O03hMkwjtk0XWfxxwgOJBCneDq7lNS0Au8x03myLFtmZ7ountrQbB++XXa3V7nH0nG87xAGkTo
b2dl53C9uE5RXsFZpO4pGciLMb8VQbjqAbbQeqRLt/ij5HieGU1QlT8xCu4z9Ekyf+uqDQDyIoxs
sA4qq5RtdRiKUic/f1DTMf0w/qkJMC/Us7Qs2bZGxL9AvihS1g9O6F7lmOfyubVDd2p8VM6un10r
pKn5oEqIWWGuR3oX8HpxyOdnYr1g+d+LtuDpT9VSYzZCPCof00Zp6sCxsYamjg9Dxkw8sobMAHE8
gtb7FJAOWJ76T5kAV2p32WCjEIBxQluqhyfVhy/XbsCpv+UGwkwDecBLWLBJYcQU/K7bhVG9oXtr
ruI831UUt3dcOLTolwj5Am6bc8Rz9fkisIylzOkx4hPu/t83ckQcMwu5p/U/JYiQBMLcg5RWXTQy
+AiIB73oJW0RQCEHgpBqvHew7/KqOqEuScS0wj0/rtU6cDL2MXrGQbpod2q/QUOsF+/wfizqQAeF
KCzozX43hQt6eBQhGlrirjAWwvABF9GflkBSCpC4QqqXuvoHqGJ8UrP13LT1LE+1nnHrgMY4DNJG
UR3hYpnkcH6knVzigqsDs5aUs3nw+rp0CG9Zh8L7fVWlynjTH7deTbQ4EWGmvVaQXDaxtH5gc4Uo
CvUFDjPw5r7l1Hv5lDlbWdMq93qWlJkoup7ultSlCiwus76bVRz2fpctvh2bmwxJ11LxZFeWaNZj
aTicLhxwG4KcnsSTi1mILhxxkLUv09GLBfM0zkD+ngKGv1/hECTs1cDHlOJe4kMXoeiM3MR9kYO/
SOtpxk+G7npAr/133RaLaX1SbuWilxHFrX038TyZ0Zra4C3TFt/4ydECOdRGw73apyj0Gm1WLqnD
skQfB3DOpCnbYELgRc+VH/qGdL/Ky6uk5lowrO/xdkyiSGGC0x+Sv77GtmbwM/jeP3438CbzLLe3
MnQDpchAz5cvO8sUjbiJo0ft+auGm7CgPfGEq1pqgAWjflDual+oXuJ5cFNNupY3fM3A2RgC4VOw
/tBK9zZrtx2KArtXbVEU0r2HdLZ9DGfoEiNg6P9rq5l7azJ13fmbXw2DrX8fBEU95e35adno+Emm
EJaBXXBsBOqUM4Ua9Gk7xstzN0HQfYI1KAlhMDwX1q9tE5+0n5kZqFq7lUuKsaJD8r3DFOIWDRXX
TmcQE5p4KIETIur/At6ujgySDnVWHvzDFWAWkgue95rOErRH+RXC8p1c7373M0fBDikiYlRBeQPR
wwIDUwsSlb2j5qY2Yoou2rrcQ4bWvl3soFkWX0EsxL3gGNsiYZwY4IU69s8XtKmLWiKaA71F4kVp
Y33wss+ykIy2tWdufXL9fQJgdzacfiVgCWn1oiUlASFjXqIV5IOWLTrn45XQhA2LTPZHoLXzxltG
fMumXaVapYz/jdTpGn0rK8y8Vd28PPwuheborpE9lt4UepYfevpzVmQ8xcrVTLSqRbTv0ANYKm/9
MF0TqSjMGl6CiTE8IjFhRueKuP6EQo3GoDNqCPEl2qHVDl/9/CTp7A4xrHG8ZoFNnZO7nfdZKyxz
owEJ69reNvsG0VgSOVvYKjws1H1JL523tIwhwDmwd3uWs5bifhMjio0q7ojD4u8aKG1NqDCJLVSF
VLD2S7sTBLIogcFdVfaWp2eHe+JFtM9GksxNXhlxZD8wwf0QjAwuznDgo7ivyrKNcW54iV2W4p1P
B67y4s4N4lk9PSGcG/uk33x9sGtcel06YzlZ2SRh6HC2lE0PSjwEFjj+uBVpix9tmjBrwug6a8qa
MbiMRxINaaT30EAJ7NN24uyNy0GlNfsGoxbe7qCQYyL7AgW+fhHu7XjjX52pMu0jjHYY9fkgwCBD
QNzq07MU7cGlPxBKE9mSLi14sYIZ9LdOzDLl6Kicacr/XJCSSILgdBOzYp0JGN84+QuGrWcDziUz
FPUS0/xUMc1F6NECqd+ZZANW3UpFTji9iGteZWwKkEjoRQgyZDuLiCr7wRGa8jjtnvho0hu2XIWe
05B/+1QJn8tm7zeD8NAW4uLXuTvfjaszc8MwtVAS1zJiI0DbjP2EGSymYnZ2Xjhj3sWU6kaAd2DK
sd9iAGgjIb6ZVpwyP5kXCRta2B1RGZWihmuYr9BTmcL2e0SprtFO47GdBwb91tfTCF2DSk4bvr70
0UMY6bjs/lm7N3lFf9fouoCyLXVZwhWbtopl5mqEOK4Iv2L28x0am5BAcNtX1i+6mrh8In4cWjif
TEzBKLCp16a47Ds6A5HNwP6Ly6epdoKa7GtkVQDjX3AK8Z3oKcPxLnD2440WfORqT9LEtUombsQY
zPMXGAsjSwXriOtwLjY+hSpxDBk8w5Zy63Pzt2giEdYkCGr2c8Ht0vtEjwF139tUgQ6AMI6hoUeN
5LsZ/qp0uHjawBvSxd9WP/G85mGkXYd8xDX2V32+Phvg8++HO8zGHSnWKIDvc+STy/krmf7cjcTl
/hBxzgkAns4lnfkvJ5qaRyXPh8rLVPgew7apg3KOn1TIcn+0u1ynFZjc6rNNXcCzSc7qTCF6BYjB
cAVbYj/rolfhkr0Zkl5ldSZ61jQL4ILpLRKK+ww2jK+1dkYOPwi/k19riQ/8ofQCUFulCohjbMt/
mIiH82ID8B3G3JqTaD/a2IRiiy7M9au6VBZsGQ7eZN/EeV/nerEzJ92H83Ye3hL0jGS0N3O7/4Kw
S/WCPH+9dhpmbDViYu5V6IK0C1zTCaDRAPHM176hYhNtH+4as7SHnsitNaQLaQf/NytUqvCZH8r9
GtSXVH45hl4ncsRytVAsSybP9AISUzd2MrT/HzWzuU0e5qhB03FZDz6SELHtu20ArmPNOB87gYwg
GH0pz2U+Y+B3aYexFAsIaaiBdV+yCn3CPrPsClffTeUFeEgNem+c/MVVKHamCw4zjdgFwZ2Ra03t
1tI4kIfiM5Ff2Qmwj9wnA/eqyx8W8b3FUW2WlHkCsWaOd+L9LFCfZYRJrH9jFKBC+Prm6NYqg78M
/Q1DxfcTleYQuWGsHpGzddmN+tHNIFahk2E2TlGi7RaaFHnglWuDSMb7L1EQdFFliDWeWn2aU9Zf
SygNKOFgrtZj55bC8AUjT5xB4iYrfRf3v15XeqRpTbRwt2frsH3BE9ljX/Et92joY6V8qNbfMzcF
PmTLta/72RsvBfaAzSxQXYASis+n5RQGZJy7wYY53qpN4MIyPbgnBigV16h0Wz512RXg33OV+T9v
3FvXwYdEp8rHe1PKLQdjNDqhOxTfyu+1R4N7PLE8zQXp80ka/+BvqaEimz4PDHjFwe0AJBch06Yt
/HFV+qif1cxvHLg4EoPHYu0ySnFVlXR40lqvaMILGodqpHp7MdNN8rG4Z9/5fMta/Xxi+4zmRLX3
aVVZmKjNRYDjWLsT1taWNi+ipTWziz+S5sX5ZtolRHc/WfflRn3Egoto7n2y8QjiVjouHBn3JCOB
WR6Rot4Ao5a+YtxEKyHQNJK6OcZUcMu45Y9bl8evIxbzqoKNn7FMhgcHFXvS8imiFesp9n34ErDv
9CpxYzyCf1ORkcOS+yyvbd7bN1jpZu6yTgEncCqP/7z2Z3idSMLVRmIUw6mj9JJyHPLoowYqn99q
lTPPtrdf4jP5QndX7QB++AqpDoaLHlXjLw8x91FYj6FK5JVNm+vYkgl8FnpR8UyCL8eIbM7mr6dH
WMDHrgrU7sI3asVj6KSNXQvCjyOUZ1UUYskA8tHnmoco7BWsE+hd/C/Rdi+TGlGSQDhGprm6U39P
0QSJKZFRCk58+utH+CeQCymTdDq2K1fkmHbqYCFXbnDyS6oTLeeNJByLvaHgePrqMkD5CNVlR9TY
Ngsf7J22bAs5veuQJjCMJaKXQr3E+lBaGvkO6+Fggj6jytTTJSeyCuSl+mDOdY0covPMOXdRkc+h
T+UuwpRzVZhFZAWMZMZ7JFAt4jpMDsqB7y1KtfC5VQoybr0rHl5U7WgdXCESsnfIDl/ls5Q1INTF
B2ARrDbMzQfl4ZxTET8S4rW00gSbcmB382lGevJNkmvVgg9WxpVx2Aps6owePqzx6/GEBcTsMfMQ
9GpYgPvQ3CPUHfhOr6WUUM+E3/fprafz6486n183BuMOBSdoeu29mBEGv3mE8leUsEAeii9BYVbR
ovl4/JhJVGiDm8vkwtKrvG9k04EpFEbJF1KBTkSiKq2OPHMg22R6sEJ3fU0Pq42sF8I/zCWYdV30
bA0Ay5H0Iq4BzsewCxMpw+2VJx6JlGqyNdHlsJ/eZFIH2BaLblzYbmrOv6gQm30MTo9q6pG9Vd3h
oGag889ONUtXx3Y/AMU1sqFkAsWRvpOiZitaAfwmsqYvFfdRch4hEmLdOn8ASKRGAhgy17FL3mfB
PPkfpfenCIE1467VOZlwCyrqp4rYdP5KpvQRhodsQ+qpm6nYJGTr0POXJ1QE9jYkfUNahZTPtHWa
7G8VLfX2ofD9EgvlEejWTaAsIdzWkfA/dfXS+J8JzM9/c77K9O91zP/tiKM/bGikxoOnplTkCws2
DD7A2rkCjqNCCDHVjON/z5Rp+uykA5uGCbb3wxREuPq8o0wcOrosRIIn9OW99DbybbKD4P1b4/+d
6Ik8P+2q+bEEqhu/eWRWuijHIyt5EpvjCnWBvd/R9opCGntikoLWKmh4ykIzz+4Lf8Xu9xKSxF6v
JcHxMirL34Ylh+wLL4SeXca7nytyjQyecryDZ2xWgb8Rciu1nFzqQ1mq5LydrMBum7B5ncdUvM91
ADbtZC/1ipVzY6ui5hl0I37nZM51IAruTnh101vbcTyimbJbp2KYhlR91WktO21np3K3FPLruAv+
TK7gtoE+HYFufPVb8OJJsyzHHtl5tZBoWWuts1v0Vlk97ltDRJzd7I1VQxThYdqPPWKRfE07/yrF
XTh4ul8xqUBA/mLbvIquODwhgOvYmTSliRzfLQeo5yOnOYSZmZU+grdXHzaoZwz5DmB5CKUBLUOH
9npGfGpfuwfi/EMjm11GL6jrhorXXgchvcG2SMlnVR8g4vHqvr0Gtghfu/7d3vNJlEKo46HricdJ
tBTdQXhFpR0xeXT0ZBO4adBoNwEe1pulJcqB0RQOrfbEl55qm5IY7gWFD3Ce+s43P1x4Me/YYgJn
bsLnVLnbS6J3QVdLscbXijf++wGnsYfDFGjmSe7bOZRqyi4R6Z3p8Qewo+p+yvme+1L79ZRZ19PM
ePaoxdSqJNSdl/pNjBd/Ifi/LqugWxHFnliK+1zxORvbUzc+A/wppT15j+Dn5bAB1iR7L8NVUyNh
FB7oVXjOHDkjkMrQECMHEoqqxHMfX14dsaNRycTeBM1G1AuHKkrZtzchmfRJvCSfsqCrd/v07iU2
oXC3sVYKqeytrk/pfi/nLgNdsu+uXHz9yRSefm9VFMs1PwAakGXnXEcnzz4mUJtjkeN7pQDmaAe7
MfTYWk6NqPPC7br3GvLTPdnMuFN+fa74D0kTe5wNqyad9uArpsJFldc9k0xBWvtXOqtSYmrjUwyF
QwE/Njs3FS8320oQ0+Q0Q/x5ai/k3/IhGkc7cSV63jJcwGj2o95WT9Di5Ykq/3YbDaybx8mC7qny
6mIw7QLS7gdS+Q/kGfUzYghXAt5SPR5/K19/8KVtxQ2TJh+CKO3NTO2ac3XreVXuKoeaEcKhhJ2G
4jQrwZjqeG1vOhEqi499gJ2Nz37aT4vBTwKcv4n7YxPLjCbnEcbtGO5lRzBFuDB3wwsnVptFt5eN
Dg7V9ZrBj30skRixB8fT4hBlx2zyNiDz+vepiweERHalvxQ5LMDOmNwES7p3HephE2gz+Hz1y+fY
AecMsEmtMSJxhTHaoM3pBnc66y8n2NNBX97Rl7Io6WVnQ7jcHjEiTzWpfgWxXXoh7Byfe3uEgJUU
ZULiQ/oe9US24TY0y7kEg8Xc039CqC68DUThPb05naXGkQFrMhe8jBzbhNTxY9nZ0Op8QKRwvRBf
2BsjyJLHf/FDmqVy+LAy53jnzxHtyFIq22fKczGH9e0D73zaQx7RpS60DghWRjJoc+++JX0tpbQ+
p3psE4cSt5wTPSvMcWS/6t9L8vJqywKMmsEzX2BpuczfN0w5IZzIVE7x5lPOmZLPEi/1d31t7fJS
24mrvFFc47sNjqANWEgF+Wr/ykDrD0p02qoO9nzGp3CsT8+t9inB321zygGGoXGBPyVfpcPbFSO8
7Vm11bSINn9YONRzI57FpMNe6vi7dg3e0XGAPW03EYheqXRFLBuXQR7SZFz6E5/dun7JabO3q3gy
Ly5oOTn6Z2PfXGWgS+Bc+3RYSCl3CIutSa97RJOkzpo4KP+0BdAU2co9SFecJbFoEQgdr61TWf3k
o3YWSwZIIUlbuJNZY1htXECz5KtL+JLJ/bRHbYzO+6YqE6OGcKjXMCfjHcpZho0AeFCxTl4375ct
KA+Gr2bBiT2eb2C0Y7wq8Zfbd2QmlPlHEWlYjWEjy+KIAd9YwWEKCqvRqaQ/oSN4wKeXpvdARFtJ
ucXxiGDqnscpiz/m145cJ+1vfSjspMyx1NYp+zzVZQ2beuLbc2NdGt2/zWrkFTi9OdbvHMQYaI83
l4B6drhCjfsxTIV9DNyCf3bYMLZBGLFERcKYXEsTaib6DM8K9vry1oMrpzbWNLEC2PXjIqFzY6gp
c5k0ccIWi11EbdhzHQo+r97ZM8TMMnUOgJV3dbRH3hlVWkE9opf5NPxESnc0toEqklug3Oh1ly55
0dwe3eEDyvBhK/dqOFJKyBmDFTojl4he4Ozo9WuZZhVJYCSO9T4Cs1c52OG9ET+fZQY/U1rhdgmE
xc/6wV9UtXCXsW/V8mVQIc4ikdsuqZAM2EkvUE6njvw1wd1k8CObPwJ7fDp4xpGJIHcAXlvHhyFM
iQhbjhf9V3GigKadVok0MxBH3ko1nVC5fPWYkJIk6srlgMZc/KXEWX55nSGj8/QF3k8hRgd19N+o
ROIZIE1g1COeSwQa+OlZBR0Wplh7++CO+Aealz3DZXEh709L3+C4hb9RXk6BCNKwJuMIGP0OV9Xw
W+uiCnUynASaKcwNRQDzZRhfzGZ4VbLPISJAAXoGAMsdCc1SIKKxSDc7eqC8t217lyquS/GArgVR
GN4kOGCfARgKeg7o4bPN/SmgqQC7V9cqKWNs4QMm6ySYIV5ofmv/u9u94lsdstu4RqwcVh4LniO9
aHCFWXCvejsEkiWEmEhaDfGm9ghZ/Z/+ROT3K65SMcOukBiNm/+w6sINCVcd569OFuam30dYmZIP
PU3McEmLu1//qmMSS5Ckp1fYKscD48kh1Sl2S83Ip4faHQI2J1KLwGk/h2LeOtCngRDBC3A0BFj6
+FRTYVp+Ub5WHpzbaXdMjSNNP8B7OpiFfj3ppjzU0jl3pgDqcf/MP2AOzN3GURmbpLePApcvLYpJ
Pe1j9JZiMIhr382n9SBpO1ayolVPS8v3jgvNyGibqOCqPIY2QXYe2ygl9/tpw+jxZqvXwC+f1Mwd
6a8L+vMP+M22CZoRFKN0vurzhrJN0EreQTsMMAKsNa2ieY1SlEVxhvMBiZ3SyJgT1UpOeqIuSSe1
wPuE8YvZcJ0ZPcSozIxgb+Q1AzKOoNB06qjS6xVyBXCr7MqJAjzujsNGPWkQs9GMb3+nvwBWSM7v
ALw9LCUXt641xiq3PPi7f33NrJ41xMVUWd/VollGBPIP9QE0a6v448tZRTuZdz7pO5gN+P4AFqdQ
oWPR+w3+nchevq95HY6/2d2EOtk4Czws66MssIujrUE07HtV9RPiC8v9eXBUnR91/skMTtmfN9iS
CEH6K60a2MzwBt2ArUWX1yAFEIYKwvi7QhtWbM6Qmidv3u5iscEOa/sUf8ahj6ie3sYAtHJKSMqF
UDfgdi0smxP9W58CE8MdUBEWpdTrGtpEEx/3lEPAC4fwEye+gyqEMMl39OxiUDo8wkfiS5Ux/ap3
jNE+Fj3aKiZ0wIV6I3U/kbeUvbizc8dwG10xyuxQg39WP0EXNR1SjXOQwEYLS9JGeZLULhOelhqs
tQavIEn7opHfx7DxbSYRuUiVcL6Wqmm64o0pkmm9o872sPEI8dTi+FN6EJrfouaXNrDf92nDt/JS
5FU4EVaMRugIuevzm5AUm4bkSCGNeKgomZ7Yr6Lm6lQOjMkCXN1YmnEAtKx2YS3mJWiB38zNgDB/
d3xXlQIeqGoxAdvmeqbH4Oimel4qX/K5SwHbDWJWbWu/mESxwwekWb1FG806VPBdaRF4VQmXx1x/
ZjPkSkJUdBBW6nj3ZcFsRjV+7266PiXp1RQq2k2FWKvcYSPcigIA1+z4Map8CbjszQ699OCJxc35
JrqOlMnu8loOEioP2IPBbu19AEyn1k2WWOl+PdCoef5uLSS7P3CX7EZ2HUvzZKeh45smuTML6P0+
94m0pb3OOVtKjT9F+Q+JalbP0Vury/bcMSlDOq6OHRdqqXCE9FQYa/lyphn05r5hCPEyKQa+jxPF
/M+3PWrrRnt3lmVSDMme7vKHfz2YzVGnP+Owj831PATguQgyIyePLPdjxVtoIr2ieTy5v42Im8pt
NztSWXrVPVgXr3v9d7RbZDRV+fiwDc6GhLQxge2VcgVKgxzCNpr9Ul/mT1SonQYgkA3wQ4Fx62/V
q9p58xWXmHcJ3n1YfqEQ/HzXPIrlTWOUfS+20/QGXqQbA8x38ALvdbqCQPFTZpx0uiWmfFfsU7Wo
GtAvONpHpO0Kl8XeY5HnyvsrO2t91guRqWHHgxdbB0ZGlp76atT4t7WrRdiTR1lwAQORjy5nAnSH
7Hj6qcVz/17BAr0Y3I6szN4FHAb1rGj1ZHWHIblfYVe62aoUW7dTwKscRsheXrKkSpXhBnWdLb9C
Hu4ScRH7tG8hr7A9IYjyQ3XuN3bRF21m/hKz85t6I7j0osebIveOJmpDuhtq2X3oqjPKjDaUxXyO
VLAia8QsOfOn3fykj+RkU9hJyl7CIQSKWGVGPR/VAMFRmiLTSvOOPh/HjywSdg6EiDck1V0fHxT4
QoPgRQ3i3mjwX1YGynK4h1cq2tNCUgEHDY3ey+FrtpXb8rjTNZ/gzWMMG9O9E87yW3BQk9/XE2Za
fTUdtOumX145eXdXmxj0bm/qnWa934raNZzFCQ4U6q3RTt3jLbNRsLoL8cxP8EsYkRMPq88qw30B
gRw2kEm6g0sq4zBHkXYXLfjiD0MqgeYSm0OUdN+zqpSHb6MWrqsxv8X5fyo4hxouPlAaTPvIa7hi
Rytp7mrGqZqBz3GXQW8R1ftjm987TqRl11/ZrRyoKviRu8LF7qbNGO/To7Y8l80MUkgC79pBkBWT
kaABq2pzdEjVSfAApFi/M39kpEcomL4Uql3KhuxD5IrnpwjtC/XKGMUvaUyNXwkhU2N8mFgPu2oY
O/xlLih8nufucKB9Gawmgj1Ly8vOWrdkPwKwQKNXHPqtTWj4oXwPnBmgrqM45PtvgQgD1WInwyLb
drd0iFoqiSusSmE5oEQwnBnv8Ko2IxxvSsXU4gwCuDoSyUOYheEzPE8h1kIPcVBg3MNZgviNCPnd
mfk7tyXZaokJXLRBKeWc4Wu8elmTEXbb/75aOtyuiydHn98jpzzk3aE8SKOGakHIbyHFdsgnroad
UHqzw2RL0SBb4xq2GeLz8zZBTXO+ZhGWJ1qjd/sUL1w/0UXvAXy5KI8SJvuNSniH0J486PytMxw0
s+SsvMZ589gnTJgHBIw8kcWdhwzbJGNfCRZvQem7UOngJS/CJoumG7ReQXZgfvdEY/6+LYDo/knV
CkpyqQPBSpUjFOM8b395uXT0NSWmENXcWzFa2wZJ12iT0ueG8Nrr7ly+u3MNIPqbek/irT2hqo3E
OW1/cpUiUkIIGF6f14s69cbb/hrJXkoPPYzk4z4kE9qqtER4tcstLW6qLT3ord2T5q2VVVBhZ9Ku
3pitJ+/vNJX/TiYbiYvxmFx9lsTu0AC1F0ChFaRazXoqNutVQaSODDXnXR9ZBFAdDIzpF/VHkAHL
wGg0cmiGqcooNpmGCN4+U1ZtoPE/+S/v6ogjPQw6/XFTXMcwFJ+Jwx4xwyBY6v6RJyXM/uD0gF0M
yXWVS9uflhfbyC5sQJjS30lA8BQkEJHnWHrBzxtLymEKe6wbAeYSCyMpPkDPVwJIF0LNGwyGrGXY
vkxwSzg+5xGsmPTPLKD0R61e11pKGn5jJaHpNgIAlKqprvRQ7DKwmHCLXg/qHOPibZGhYbDYuQUL
BqdCYCLNfwcz0sbxYsVnKRImJKmRupjLtG0lR+iJu3v52zEJ0HpkDfgT+8ZgYa2J1tqvBH1AKE90
EJUTHSDqxUeAxXG26HiFbmJtKjdU3Zq1PGepGIGJlSDted8jw58iEpFUYpjkObr6ZWSf+0ahzDfK
BHu7iEAM6SP2xbIDRLj1lEqCs46mOCmJKfTNLXeR32cIsokpN7k+XRuqdGfQNk3OeddV9kyw4SyB
vLHaMHMdrl/uRKJMBkXriAOC8q9UTgrKEDnE6IEc+ARr38SteEYNQ79I+yd0pBQlh866CaaVT/4o
wvtEUCVmTQjFwGakwJiBDRICAK1eSNlK6QbngRiA+c84QJimz3BNjrM8vixPTJRKkMEvnt4GSTrW
PThLLaePpbBTPEx1d6Hud5wVbMDFlcyfsL/rFt/Iq8w563E/Lbu0+UWxowCUbg/uK1JmW3es9hEa
ZiIqTmXFaguUXEqZHDY8L9byGfwyzgXD8eyZwV0WoBhMeryZm/d970nmRp2hujKn06iVnyrMkQGt
rrZ6cHE6dmiK4lweaHPb0qDSlauWK9tI9zImpKKN7l6WgjrbB7ls7ubfPuvoG2+TG1sftSh4C/43
RYIjXIJ597OG62aQ4CPgCelTi3PDjH/PnlB4O0fdEnpocy9tc2RIqGvgljlgqjSLVmqK+maLF/AL
lDf4khXraeYVE7+Ckp1x03jOzaaEiBMgTZOsaVJCVPe1fDuHSofV2JXWE2M+D0YiB/hvj1VgH+Za
Rp1SeqyWI2UD6ki/Ej87k7jfXmyxpmFDOrpvihlBlAVV8XuZaMUiaSyyMIaHrFhLmjUsoWc4J6VL
eIPUIhNmIutXQX3gU96FmghGQxIrZqbgBPcYhlJfe0KmszpvREtNLmEdEeib/84afe56Ic8fq2Qh
7vJ+N0uNTSfUbsjxOm74z9C/+NAGhRqePT5q5/i9TFMgcsR+TT+WBwNRdVAIrwqNbdTlnZ5DNQKc
tuNpcJmnmwky8qz5ShQoZHGVbHIOV+7w4lqRYH6ggW1Vrdm1LvXDXwkuzv9tsfyofSedSFjDZO8d
mfusYuCz9kScMpo7Tu3dD6zh+iwo9u0QfOdojLchY41YA/7iCNtb3W2li/NiBNX1ezO5XpBRfe7W
7kYWIXfIavc8r99OKSyV75adDW9EJM2SgRSwjVWIfKJ5ji0U/LY1ZALS3iPuXPUdLRSKEmkK69db
QlUnu9xKpmKYPXfGNRIBNPlaR1xXUARJlde24Hm2FcHTYZyAZeEPOiU7mffoKdkZejPUBGkQ5daL
yXBM0PegM+litWv3mIeih5XfgqGJwWoqarpxQtfoglEbOq3iHleCwqgMSq9V+fFPReEyho3jJXwk
FuFMChXE5eZgShux7HAT0Mha+7X4Vu6IaOLdv1nlgQ9ObcYtBnil6/Bbm1Hvcv1fdGokUNr4HKyx
8mgi0opL5Mjf96te1YzUXGpYoMkU5FBs+1JKx7n0ar1I0JxA7wqBJ0BEmTsM7Fz64WltAOv3lyzd
t3vqUOhM9ZfOvs0ZRRriUzvH0v/m7k2aqAoigbYwwCZkGAXWb5qNCz8WcjZAhmjDIfME37KqrhQG
Cdk+eF1yn0iH0bq0KgS1mdbP0rumYTGJvh87+GFzcU5khWU3HmGQtFzfF+daTCd763DVMNZXeGx/
zcJrhfuXzUOHIkjArleINL3z/gFOIibh0kazHgWgf86+xNHTEzMl7zwtLVIpNo07zGrIS7f97p6U
2Mpwz8NvCe5LfqxKGKD/186Xpmtf+HO4tlkXCmRif1sGjxLmuj9pBIcrzBV5Msn7mDFTUC8YdzRy
U9Traauv+YvhQA+Oop+DK1pSkDo+anC4mDFVhQf5/9rngh+seM3ckZ35GnoiaogEBzFzAQ4eWWCS
moQ8X2H8U3afykqzYFHMrqXT3QddHuu7B0IQLMagDTIB/b7f0paJzT8+eS+JHQ/ZZJCvJQh4pmnK
JULYBEf0HVpBfnyrzjFQCVww+hG1qbts8B/UOK/v8bo31j02ouIi5q8mvgC1yjMbKv7NzzjmMp3c
cqMU8mxnezeK7jSrPBNw8alzG6rjqB8sBTslNo2bJDzVwdXE8z2kISl+/gBImGkIm07/b0cPCZx0
Mhzkmu+L+BdXWaXH8uZIC93SW5J5IvvG7oTJF3ss4HK/6m/x1oE9ZecO8NaHUUQLppBhYxjSm10a
so0HYonsTt/4uX9N9DFq6xAFRKYmBqeIvBEaLK8HX8WOf/4E8Fqzl4WLvkajoFZ/EEAonEcEFCOl
USWknxXT0nmf+gyO4b9deOot8TJAnz6th8TGbfPg3aaryiqXHpLGT8ldFdhOXptuv5hqb7fgLjqx
svY0yyfW9ngGo/bjRSB96UlVbwO2rwT5GelP1A9vL6nHn5A/JlK0Bxalw5WijEOR/+w6BywQcIzV
vgbMyD5twjfbvavkcLbhXamGqB0aS7mEtToU1oD9dc0IEN3qK0v2nND+CW5rC1vskd+wWBQk0YrJ
lHkBaxGolW+t2DXBRuOMPesTMcnXk2X/WlahUiIFhRaeZ7GeJwlIHwWvOM9SUTmfsYNaF4Qe+jCn
ya4vUBskbamnd3NO2RMQdLxhGA7lmVV1flCZfbIPhScKHtj/S1wt17UQwzMlBhLaWPlz6YSTr9zp
J92R1JeyAg88b60nOzbdhNpmUje0OiZKAy+5uSB4dZ77Y52gH/sSLR8TRjZY1Kz2FGOoVBLOZ9jS
Gj4b6p28uUG+5gHPxc0d6cUwa9Adr+aWHyi0Pm2HplUsdnPDh2ug1EbPUFEhCE2vaOyE54tOP8Tj
pkdjUi1nxXqiRer99WDGKtNxITBmPle3dLUt01ameKHQ/5VjJXx1ViXqHOswr3Ss7le0mUIPwVVm
nK/U8A8IJCQTFeDT0ZF4YL178xrQ8G9j0BqWNuW3Hy+0uc54o48WthSHa/Tt0pgfTNp9OH5VoylP
BxMt5fFlakP/9s6kVDqctvX2EedPoh3sudYJJiiKitpy4W6a1uSwCahBrWgkIUfuUXp1pU+iGSe6
ebdm6U+L3Eaf3jO2xR1jqTyliS4flIpWnY9OGxt6SmZbZnktLCXgjTDUS1cVOPqm2m4haPc0EG1c
EZebDpz7cCjfTjdRrl5hp9AgA20h4KVAHdX6L6Sla9Bw0MEjw46Nh5BpL4xUsQtnzlGr5tMI6fP5
2eEJWPb9U9TtsZh/O1+SZukrRfEkNhqquuYIGIuGt7AlZZUOfxxCFZhtSbKCuDYLLT/xIfMeSYSh
OgXasLbQz/xUi58bh8SpBz1n6GjT8zY3y9+JKSJye9p9KjvXRvmw+d+BxP8P7D29lgiZ9asN+qEQ
2vZAbFDRepP82CsEHW99w6G13bHxvWlxzVHq4zq514/hzYOBW2U8SEHythDxQddCXPQ8+ja+Iczt
V7+n/N33fZw8DoBy6FTOqk49C0ANzyneqZJ7ShiCsveJwsUApCx1StpjQA1vkZldOIK40UMVt+Fn
YnM/PtjFjrgpk9ITMzFTnIx4q81vzek0aRc5t0+/mVCUoCKpAsRu0Obq9Osgx0yfiKVtZuyBtU82
h8Ft2HoEp71U+5ZZCB5oSSN3qdjmiqUd9rsaIKeDZ53fKasJKt2YnmlFcl/hTlYDGUNtuu3Ds+5d
iCr+/vbmdRIicVkLT1WKAB3prmqF45otG3Z/gn1s9R5yqSh4zjxenqwlucTBmpCXypCOyY+YAl1Q
QRRj3Xnk3nUgMHJq23at53O+Svqdek3D5VmKapNTAhIlFnkyno1Dsvml9YDyGQXV0MWxJww56lSF
gIRsEHvncPieZ1Idmn4xrdbp8KROSq54cR3T/hm03mcJKSk8Ng5F5UQj8MlvYgDIon+I9X8FWJv9
jalrrKRXmcXT4oHfXWOkLgDrVg624eeu3UF1k0zrFBIx7k3dTSaYfMDgvyi0jc7zT6FADgumYwKi
jRxjPTaUe2JDq89mWseGaviDrA1kNyWFIUQXNICSnildoBpGL0gPsxRTdwE6wPqr3iY0gKskzt4G
Kdbc6ITVmwoPWF+1uukfZ5z+b9ameaNv1bPEEKDjS6koZDRFL7GyBZfify/S98sZdd1HFviWfHvi
PefsT4QO6XT6NVRFOA4KmX1A6soqCjyrJLVhaR6xO3JRVHrwaZXdKYg1e2e4EmgYS1BjHuhvP74P
EjN6ON7G4Ny/M19jnhfClpuM+S9ec4XABLH5xQ1SESyeO/HUa2R+9ABvahhhVwTz8UdXLsgevZ36
10w/ru8w005kfADYoUvgJlENTUwEiaIjgb/s+OmbZ0dkfx1V3UZcMw/yQ0qU1owV3aMKXB0goL6n
WKi6z5ResZOHKaMla2+RcKB5KjfrSZVL/d01s4aZdU8+vRe/YKwMxfvEZDFK++bTfgLkaqa1+P2E
5gs229mN6Tpi8PBTMhFUKbGZkOH/UnSSgXRKN3ErdyJW2zQIOZvrESMjnWGtrFB+g2Ufeb/vdIbW
KSHXiNNFBx5qN9vsADBPeSJeH9mI33x/63P0fTK8dkyhtTb0b22PcXMyGScIYfYz5rZAS3oLfLDl
tYyPPtp95kk+48fQaCXQm0JKYw++o6juHWuTdIccdlrJ1oA1YEmPCDsvBOXRpdKO/dPzUbLY9eMm
NJdHQylRA7uiY5oH6k4w2FHiGlfZvPLEK5Dk08Ltz8q/FEdySnGhGS6Kku8j6VnD2xUHevSxd5ei
mjfpdmE2gKXS4/WOHsoyypkZLSXBbRVZMeMkBW71EMDbrfMWjc4lgnx35cf+cLKtGn0tMweOsMvu
yIEvrOdoydul+J6tc4JnNa56WYGZkIJRsBSi9l+Cdu5Cptj87HEsfDzylTscKSMbsezz6CQOVrhn
3/Vv7IsTKNwNLUwB+v2fcW26hTDgDV4Ut9nz2zIyA8iX4SsU+VC9+Ih4T2vuNhKAo79sPRcNZFkH
GIwDkEh06QTlxDmoR2sriQ7q715/CJ4RjYuyD/Nbhf6P3gVrziZum7cYLe69vm/GnXIW08PIM1xc
ChE85BVYztaJYCNaqO6iU9t8YOyMyqsUO/Y/5+0jSa5wnZwE3V3emh75RKTKVPkMYU8tasYOqULL
0ogLdd+AohXBL1ivI6KQiMAjjEgw34JsKjdelEeeJFUOsi8gdvYtdrRGkXb/WpzbPtOYnCMyqAjE
fUyPF1A7bUFaFcib1EkIF5QkVNpHHu6LCwPe5nnVYryN3df1mrmM+WybEGQwZTQtYzJD7VbQIffM
ZknFaS6y9tR8o72GRZSp7l9RdNXPFWYAOVwkklHtqp1ASis9bUhu4hLT5lIdYDDn+DomQ5ZFgSUu
6rI1jB/+8wqk36klwzV8lflEkdn+JHich6H1XUz6ltjfvEUNcigPZHjvsu2/cMn31und5WvTzxJ7
xEb8ktlgkSx7Z0BRzbW2qRVb1bOMa3iL86spxGdaV9Mwtr5LVowyhihYGoqdAjhRtXpgDUmIacRZ
Q25jZ6P4xE7Fms1oM2Rnziyly8Wnv3eOlzqv/ekVsdhNY2l9bXBehc6FejlBKIroioy0d2LssK6B
PUG0ax+hzk7ZjnYpStL4Mg2KM9NXVWpb+Lephrt13HgFmAwI4v2R7Rxgh1SwLbo1gw+lbPTd/Dj+
98cZtQR7qGuO5MxsI7ztXU5HKdOjgCD+p/xC/IpkXW3DHSjCgqbL68HafOJgUbxabw7pjvcGnJwr
OQkbhye/wMi7xcruwKXE3DAGEVuvsfReghgMUTIblZVdcHEgsYu4peuGAYR+iqQ1u4LyJbb20FTX
AY2Eg5qABVxBjkYlcTgkfG+/rwgyuO1BCZIk0nkZn6GuuHUeuhHfd3OLA20nm8fb8BUH1Xwnu60l
Scs79Nclhv3ZYoK6JESeMfkD/Mn6UM2u9NLBWHSFrDZds3feCwPFxcvun/KIV3RpPzUfXZTGrUBl
cZUYqnYk8dadx5lrVrzuD5TDbHcrK/R01m4JclOd4svoaGOmnKU7UFzOHvhA8uPGCIP62o+zOVPQ
vU3mmRNqG2iNsYw4soPuf7CWsfPhiohAYbJp/DBqubCfJcoJEmrSFzqM/yDCkxPNNoYmiR8tSVAS
DP6C/CfvBA5LJxhb9rqi8Sx0DHNTiy/lmvQWdnWyE90uEMLS5rlDddTD7uHbH7F4VpcSo7mWHLZK
XtDaHwapatqfTz+f8N8DkpqnC9sWhzX0cQtX0RsJVmegT7DdLeO7K0CrwhNiHeGg67fd30gBnwY8
tRtQhY7sQ4vFm2XCgJBcqtdjFATppsVSWNYl7I64zY512+yqRkmQR8TtWHpVUFaY0B+f3E9BzLDq
a6WsipRtJ/wvfXMU0FF3OdKa7+dH9BnFCblbnUEXkbn/RY529lGbAvh4mRm7ww/LaMA+zzQ+Ph4N
H5pLsYv6bU0WuZ8rYNAjqOSOZbzRDG5bTyraGli7aFbka86kYDOVqq7Ziyxs4OWQl4z4C95InP9T
9uND0T6ke/Kk9u2Gtiq5iesaWf8sYLcdLEDjUlRRg6kSpUIMxtxzK/+XttKWzAsNUjFPC6ALi0LY
7K2vIcG9WOBmwj5AfI8CLVUv3Wp7M8+WObms9Xu8CUX9gyWSyAnBpIakHAVaf3ozuCCNE44CdPUd
Cw8JnKMjntmHfYViEa4f/dSBUrN2fUo7jlDsEfW6QIh13u32kHlrUgNDrj6djBLlsH0rNE0oz/q3
Dhl/3L5Dw5opsbgZGifYzNlzBTSSYG4TQrg+sHJUmiOldgw5E+dj/jkB/8ek/KqT3BljOU//nJZE
z04oERrH7b0NPGQ2zKXooWZlKADttz+KjR79CNXDftU1VViEH9v9lwbtj/YWd2WMYZVtfLWIlxt8
w3laT6MHn3AFZlV1LzIyknbhbkmKx7DwTduVFoW9mhRYyIDuoJUtPXxDq1A9qjt6nOJIN36lxy5B
UTfAMTvminKwp2DVQZsuKQrQLu4TxWE8ZNX+66CgM2CDrXW9JEE5+MvXrY4wsY/KQGbCYs9XjMMI
PDe87xKz6UWXpf6mxUORSg4HqlWWwDDNCegM8BM0RPf/HW3fxysQHzet03mY+jpQVBclP5PruvF8
MNjawztVAAGpZ03HV8GC+ORAXPqcIbkEko8wMjRzNqO/2M2vOovI/8/aIzoxSc6iajJxHDMVWH03
iLcWi5dWusmGT2ex18poIEFVzyWcvKU330Gx/giSgMpoQUTUch0easHalI5EE3F001BJKyDcUCB8
1Amqoygl8b4BgqzcsAz92QnhPYPprcYunBv0apYOdBZE60kqP9obR5AYtmWoIVIxV6L5mzKbTzQW
Rh32kho/iwJPSd76drzaqHWKegPY7lHvBpDAkTP1PmWrTkXvvcXIe4zzb054/ePByn0RHpwure0f
quJu/xlp/pjAbxH4jcLrtx8N6CbN1FwBBWjnUGntGna+hLIPk8zLYnAb0d2SQfbLLhRP7VBrsyC9
IbjNA0R5Lrt9SRxqJvd9nkgMJKwsc6mFw3U/GtXcoCAkm7/sfaBs3YY8S0dAhvJVj7cYioM1yO/C
6uHhoOvqx47/bNtJncvwjfs+wW7sKq2BFusH9YDR+DNbBW/UUSM9ADTjVyirRfSI0gp3ZIGBHa6l
IFcjKB6jaFXKCkVj0M5o1TLChy1RTSsuhHmRx3/4eu4w2dA16mT6K5aZ36FEUNExAYBb2uQ3wPNx
RkJxkbPWyxT8sLTywbUCKxSMuPEtOdQAnRY+MU3YRhbOfV7NfXd9l1gi0p14+VOSZfW2G+QtRp+o
usCCCsMvB+h5UKxQ+3U1+rX1Irt4NO070z5Vyuqq3djsfG/lyqI4rRo6YN6eMSmAPNax1+Ox+2uE
MHqvA4cBOC1CwWdHb7DhX/X2k1/0Tk4EGCAa8oZlon0MQXz4/oaAodAtFEbJc7JlMhRz+9zn448i
PQ855OYZaG2hy/QTGm/9Ed7gDAU+aMZesnJ8/hjchUcWxZTrhCCfLmiVTnzoHFVp5pIEIrYKIzbF
/NBJo3u49p2Vrs0Kv4i/b3gPFPcB0j4ZLuw2eRDY7nKn+tpzZYiQ6QChXvsop50rF7iUjjMPPB61
x7xxhGu3GT6PGL1U+BXwoOzbiAPhiBzi1jXVRak3TgC+euDUmsNsyBVyZxxsVPn0Fk7VHBkJHkOM
/ommrYLEhWv+F3fI4OJgv0BG3svmTEOdIb41/QlRgy6snJhmhJ9OeFuV8qAdxLFoXLaLGlnNzSNE
riRgYTMn3ienL8CdpQ91gp8jEphovQtOGpK7QJQWXm/F23ZZ4weHHu5SphO/y2MbR3WvtfZjsYX/
jO2ueiZxvZIrRx1Am9SRYqeegvmpOW2E1+lgSJmruaHACJ8dfiqVEFAGyRbdnuys3AeuM4vF5b4R
ZwtRoZ2Myw5LTniIlSyIQlwWL8lSUnEMjNKtw89I79Bn9CElwbp657DziDcQT41cjXF/g2VnQf4H
KKpmlfbHW8Y/y3YzGoE4T0HLMNvkjigjP+u+3TWjYPuf1G+gcCRTF1gfOWiBmm24G2UmHUI+N1w2
fduBU75xVv5kBNyqfp1fgswTe4a1lIrnSTO5wGDL7K+QQtqWQTeIUEmHkVip6A+JWnl/UQnMktAd
NWWyKkI5ZSNBi4Cjmkz2/tsSge/Lv9/vfIPaCaiULPmv5ArbN/HjJn1J+0NFdQDZwsX91eQjSKL6
ozfVJ7uaW+dahcpI43e0OKF5EVwAXvcJpjOiejDT6pj1ygoy6rtJojHlZoiDB1+C3vF++tKPW0zO
g4CRRd2gtQNIuRJqU+3Vw4o+M6OyqEFCd+Zre2pL58VgLVulUid5Dx06pnJHUfsDoFvPiEUZMabs
KZyDLfMjtMNZKsDTtyg7atzngD02RS0Ar6Nj47YjeCXHcBwDP6/aUmu11emoDZdr213RP1iVVGhX
clq4VGUpjWpQZzMTfLSILnXF9GUV5m8lxnUuBHQyzzZxGVwfbLvIIej7/x5sulWgRh2Pj+BxGkOW
IhY43WNFy4lu3TkIXZdUea/1bOpp/pucr4iyJwFUE7JrAu4W1KxUDTXuYpZUKILIfPpC9KFP5hK1
1JPsrRgn+La19abhoS87yibUpS74XoR6BL+VKBWQzNXvm/xiSyLuFl+7QXTa3b2lPCqSUO64OrGO
Fi1Pwv+UBWFtSDkQ+u26DUUC9oaSSs3zjrNFCT7LU5MnV2huD2V4NmFfdxadqshqbW2FodSZEpI4
BMMjMUOk7AuLeo3wWtEd1ErTkYOHd5Cg7fme00faj7vjH5KzGYoYgMQhLkJ15bEgVEuOUPOqDk2d
zkKTb+oiMGNoyJxk1ndygZbozs+jqvsf2KGUFuklRaFruI8y5xz9+JwtIWmwQMTkXZvz+3bFuv3y
i9FiWBEGEjxSeY7Kpv8Roe/Uji0RZ3lEDWrIwA8oHTEAm1+eFx63itgLAhNBATPZltpyCWVsBeC5
2deaOE6NTGVfEX3iZ/TnJ4aT89RNY8QWC4TDTz8fdneqa5g3+6ysvhqjccN1+nNrr/gAbQi3rQPr
bqot7z9h1DlPzptc45l3FzIcbWmMP0PWcmWyXtnS11bXC/FUxXXql+xqXZG9lN0nOcILlESgbhc5
nhT2/36P04lHOsgVos4nAQ379TS5Exm9Rov+WHJ1VCM2d2aIMFN73tyQYskE/pn6HDXrn9Dfl3oY
ZwEVnygefujDTiYl78rZYFssU3lsx9n+Ggpl41p0Ln4JMJ58T6uuSiMHGinxL0iaDopuywx4Cs45
g8eybAiwZPPg4CBHud0R8elDyXT6FLt+hDcoLZhN7A5nedk6s7KaeeUbMzZyxtt14wfZBCZDREar
8CYMiZIci+yjuq84VZ+HgRloRpCzNdd2q/43z+vFFcQUmN8Wcn9qNMqCGrZQmPix1yVd53u3UrkK
hu5B+n0un6zg+PWWhw54IONe9OpvhBLVKwlKVm5yjjp6BBc4F+Ueeh1NP5lEBJ8HgLfDc24nku3t
bDiYZtQ0EI6HbLPzf0x6BMusMaHFBQxX5i4bpOvzkRPxAiy0QC66ZtnaUrnZrZ36FN+9oFD6faj2
yUf7aob1jOB4012ngze18hU9NmPMZTwdwD87eNQcgg37doovmnmLyk5uwtN6uqpB41L2y6iPH4Qc
LtrJASBhRBTnmgK8U/SaUH0pybwsAFF+Y21/xwuqDsnM7+Jq9TDwJYPgtIpB8T4yuW6B/KQ6jdq3
P1sxXIXk8y+IaDHfuz4SDDHo8bSAAT3LPR7qCVone8Odsyy+dXdJyUIiZP/H4YmCyyMHJTumw14S
xZVlOgmo7T4HTR54yZ/XF0BHlfF6N/tEZXFjNz+eWzYS04/2dYBfrm776MhlDfLvlhDKHEEjJtpq
mrUNU2+n0tTdc5Eie5DTEwAtSRXW7vb136YuMqdaa9BeVaLEaVmRxeD88skzRb3EKUIJYr8k/VqT
J8hvnN9YCUXocUJzng5XNvB3Ml7iK4RNaAZRkb90XWw8k574XgdrcLf2TD3b+92Ck8zYbr6kZ7pN
EYEjPTbHW02ybKfkmygCOVrvhjMtiEJuTOG0zaXB8uNNIuQhe6c6LstmL2XVq9w1w7c1B1pdqqyE
RIiES5fIjm3z9eysPXTnnQivyfRbH2+a13+bHb6aKP/R7Hsd2Wp8iM+w/ruP0H5pD7csEdk0k17W
Nix9+cYtyA75m2fuIbWBt/aOP2NEkzrGNl6nj37Eg7NAjTqF91KnMBWXiIhPQvC2u05j2BH23Waf
uBPadR5C1Uy0BHsxxMCx4XZz/O0QbKfYCSzlFShpz7MXhhxk/GFeA0IOK5BxTjq6lisA++bzN4Aq
sGGHNKwuxiXprHccNV7CfKjeZMSjgaGRhPQMXrP7b8eX6tjlf0CIfFlgUPPrj/p3zCi6/Lbc1ZOM
6PEDy5TkPkuFj/jQP5vBSCvPL2pq5RmNfK4BwBkm6FM6h6RYqwmEA2Y+a/1KmYdXlCDbMzsMpL8H
Qs6xDqljkCjupXgyQBTZvgK3PlhA5nhh9ckZVpc/cWOJ8ONB2FPKLVK+Op1aZm/V0MS4KgsSAVzM
U1ur3P/vC5GMVBpeMovvcfJ3ifRNlz+QEUvMc8ik0EJZQlGBh/8+r8TrYvRxJd3XBb338QPlzKNS
/1B/Qb9i083up5jYRQQF+xe90yTgtSbMvAxGfY3QbigYBU8K1S78piYgacZtVmQvHQGK/uumoIfZ
74uR8LJc4NUTd5WBSUY65mIZudRaL0W4KKOY+j3gNctNWwQdpZZ1TqAatZUdxw9v2EwvCn74VQVT
AZ8+UMRHidTHF5nYwVHx5xgdTkFGPzOxhyQYXW340VC9s3Gqq8WdF9KMDnhsEnpy1Cspg15VWvCD
4RztmJuo5E4/YQKnZxkeXwyOnQnISwmZum+0GzImYsl5kLkuybIH1yj8qOIEIjbgSQbGk9bNxVBL
r2hSSixf/DeqTtoAm3x5NZGFnryoXtRkHiRlFxeUPhZMMbnhT1jbUp3jsEqFTvu2/0zC+jQZjmQL
A59Y2qN9hL/XCrcf6ybP5TtupYUT1fFdFcSicksLOWmFyHRQeYRCRbzho4DoYkBFQNFPR4NR9EbN
W8eZWE76H9qtshS0onvdP0VE4UWGoImFmJxV6ZO9BuNJS/XnKuivCt7bwP5rvvxPmOSVl5X3GlZW
lFgRJ/lcXny58GvswMnP/SAdG4ioYrYw17oTNCi0wkb8PkK4+YyaPl8hRI9r+50TvJwK9T/rYPz4
v7XLYGqEpGVHruaaquCZ0pgz6xhZUDkOjMZpGr9b008ZzoNB2hrZ3LPKmapVy4GLptbq4qAgetKv
UAuJ+AWHHqKGNoK6YbLT2ZYjgHh5NlIRDnAifzGINhiaZbv0Y0w5Nz+EGQR7zovj3rxGULyHzqNh
vaLMHnu/X+FRoOjPVHmZQWuMslpIUK69v2jfVo4sgIhyiJSdTF5Ax+nHfeQvAbiYKyntUkn4M+L6
KFmCLpWKIRb/+E4efb3IWcWNUvXwgsp9zXbTKXt8xIj8Xglbgptmwy24gdMNgt8rWWPPRQ8T7WkD
N7Bh7qukqWp6/i9sN0RZNkjxbGMYQrpRjMj5SFmlPltEAVVmfQwQ91nzhcGD0gDCnkolpSOjSPn2
rC5vhanpYs00VN+Eb0ruECbniy2Zk3M9FVmIWwejSPDqhGyy6oYKvY8Y+iJSOEfZkcShSuc4pmf4
Ebkw1rKN66Q7Vo7wuqgBPK/hhtwlZDRIP7PXHzbfg45LjUTZoLtcGwcivQa6aiSQZze9BL6YOGjg
2VsChzf/cpStG7ZzWNT3ldvdT4owDo5vCyYeU5vSDqzYFMMkznJYbWOfdX0BGUE3w15Vh9k1G6i6
v+KSzYIIRfQHcg6dHd5ZzLX+iIHsGO70hZnL7KtSUJcDBigTEdba90R2xJcD8Q04y9Ixhraxpc3o
uGdWLzyo8wc/ElHh1qeBGR93H8x5RZjeSMeUEKws2e93PgfgjIOVk/wp6pTUKYB4F70SQPspEIOw
gjzUNmffsDWpHa2mJKhI8JJyjYRJH3DC7JVw7eUCYcUeWcDjicoElQWIUhtTNROOiZKzNvjlFeG/
rVuPbYaWyQQo8L0WP6KgSNsT/UnMfpFgzkO5lIdMdt3kORUIdhx3LMwYMqNxNL1caI6IvqA5RgVQ
LHBBOfBs80/g40YDpDCDhyBFFraJC1a7Y5GCY22+FZB3vrbEW3+tLSx4CI+SaAT54uwJAOPttRN4
HpXPbpOuckHDrzULtcVVi/F0uDcFqX4KjdQJZ5cYxNh1tkiKmUG99GuYjcEU7XAcP2toNVoNk02j
AF4ZFUKbJRN0RxeecEKAB5w+2JRmhlHZLCScAgnS3oe4ehz3ITbfFzA49fqUr90k35jAL2RdA2xm
+M3J3hfz723HF73SYz7zaXGJlW6uVUcegxroDtl04ktoNasoaaAYvYYlqhOI2vuDt5BMK/RmwYsd
OBQErel3ySZXwehyr/X1MMpMQMe1+hdj5X1TJkfRpSCadXFkHcyQru9ZX8sqWvDpHmuf1ufQBCpL
7dVi0SwLxtEh52qpvZdeXxnN4/FlOdmJCDA9MzE5Csffbd/HVsEaL45dOF/pQhh3QiKubvaOkmmz
CxuHj94WNkI0YBRDfdaAk6wx6ZqwF9BqnjVldBB2ukbTlDnXk+vowvVrEIN45MRj16ncB1HmjDHe
FSC8dduzc6cUZ7p7MtYRVB0FVI/ZqoxQizAFJfKuEljHe4n7T0AcWOILXF0sReSbMjU+IMQma4wj
i5t4BUPIYac6nCrJrSWsyu3MzcgudbcQxYOiaf1BAEROXXrLeeSqn3qc7Vm1Xd9eOptx2Ao7hSy2
/LiBZu97Xvwb37TNqcRDl0orsrpKHX9Ysozzod6nhvwpH90r4F06+ZoCFGF4QGgyRmcqYyzVNx6d
isAcvvtMqVL0+HdJrMKQIlqbn2Zanwy8VDSA8pUsqIH4a3sbigLEA5QykfpoE8NrnyGqw/sOMzZV
nql2I6BL8duh+goSQbsX452Gq2yRzOwiElh5hy4kPr2vqRe7ClpzJ/lweTcoYOrmnEwaS13PmO4t
KNf67BpeKqojyoB2qJgaxiDveLgrSqN1iGLqeI1apP2FrLWGQiaZiPG3lLWoZz3rTkjYA8Pr92vk
LO8uYtPUOQ6vHd8+Vxxqwfdt5v0OpqD22weCGk12ABVFiSpPDSPDCCGsfDbgHzBGdiZw1W9C8hSA
Lt7hDg6N8kzbT80htnmTqg5OsWvVlsWDhTFmjjeJymIR85MdX5vJzZefFJhG3NFSqFo9Ki+Pb4/c
Y9aX0z2A3kwc5lhTYbj4JCcRfj5C5K05yfktH0NdGHAD10iCMVSg2agrnQaz9ltrEPnxR6aR3oRv
/zVfEKYPRq/1lKs84vF1xA/2aOTsMY2HbwnL9YhudMwHi4bGy8Q9cEBSjPaG2UhL9rpR3EymQWp5
oeFw+0i7DTTQmf0Mut8SkJd0lptUeE1pyP/4rNb59MKs/URm00rPmzuSheEvlxumoi4ubJeYwh4F
C/EUuQxiyR6Bna1um6HdxBhS4zmGenpUbxH9IscikhVeyPzZYdgI2B7rOsATK90tbKio6Z/x7anp
SNs4S+6xcZ89a8jb1mW46SgmH8hldbb3PkuKk1qq7dcEpGyCi1loz9WWjAUDILj+Ss2W+uIoX0lk
uWetprgP1Xtb0muGB/pWrAxl7s+CWH1VfXoiWyRELIf45hhNRSyjJAmupdrcES8HDGpg4S8aOkE+
NcT4M6upB1617c02ctr8mHTTG3jtzkH1+t94w0nekVoyb7gHos+DRCHWChK5hplbrIywqNYrY1+k
iSafGzxJLFwYMl/KO5wsi8xBose7m70Fn8lvR1z4ApJ6pKlP/727VXfNZkpQTcwhReMDbvWXt00p
5i6E2TlzWX1UrUAhVAbGhJS4J2BcQwdicVdQP6Up/IySUwjhBcoe55WvOOPPiS2YK9DUxtK83jaY
87qyjWlFgvSpuCxb+u414qGNJPJ9eX1msGO48Y9GfdQ8DQGxzdc8L5vzceLlm1qkPH8pOnMFpK3o
kaCCTo2UhvW+x2EfkttWtgs6WJLpAykVCB/R8Z/ThGgqSiSOPDOddiRQHxfTKf3xEzZaZoPaTlve
pH/IUYhQ3yTd6MqQkm8tOp7MKFcwAsi9EL5mDArtmM9Iyc3SH2XCLzYvi7dVqUrC4l3o4C+mcCti
8l6oEU3pr4PFVs4glq1CtJtCLi1f9eaosUJZ0CzGYwE2NTmHFK840UijDg6EREpoyfsnCPkJHHb/
5/ung9BXT+dtcyvqcbXvMnHQYhy+cmVSDm131MqRQu5Etmm1rmR0HtRXUxy07spOwNaHm7SNI4VZ
Xh0fgdNijzoUEtEaX4VSYQK9SKt/RsrszkaQK4S+8N+9J96fauaHEL/jcCpGPSmANUjlwbCrqi3P
Bc/65TjCclYTItv6opkJLMS++FmO02goymP3d7ZqC+W7BShf1CzSm+3bLURg+Mm4XGwvbdzUvZdq
8Zas+8Ii/jfnIl7uN+0aQVG0+zMm1A8o4w0AQP6Xwrgog9q4a21+HdG3wQAPbCl0Rm5D2m6uBZPX
3EFkBrWY7OyVfkiaZcXNp3jypKUPhzYd8tFS/6PbE3tWI24gS3B7UJzI6m8DyB+SjAsYAl/fClj7
8hG7DUQDo9B9J0wJVzGBH6ThF6W2wKukJFfJSUaBlQoUDZQwyTC41hiaAyMpI9AnLcNDYMyisvk6
xQp+fcVMxXLXcntIXazWHTIADdZoxA/xpDe/SUvxxbArEQvFlF8UonxfjeavPtE69sStoP42XGq/
tovzOe/ROzBo5OXpaJrqc3nFeEqSXqHqyeJVe1dAYHifkkYGUS8t9SK2DKxkbzkQQpUSg4FeRsr4
rb+1XLq9Qoasm7ZyHyI6ivnh9L9Y9YcFFQcfUfiv9x28/4A3Kqz1YwVfwAFsXXo47sV4mIDsZ/+K
8wsYiTmxECnQJc/2XGNst2yR8Ofj2Ls+E/BbSo/D7dWfWrthF72yD/uAbjx3jcNZeoMTaExnQbRk
MPc2LC+79bDMlyxOlroJi6kx2ZE+Hb32ZdKSSx5L0hF9O3RUMrF+n1igT5Si9BoN9e5Qfn9FhMP5
5BbuIIzlTy4W/gMKaTdkRjzJGrXyMbPkzQ5omgeB2TymFFhkV0WFVs6KlJdzpNDOYrfjNajk0/NV
VkRKvJgb/SUlDMjTjXFvlIDzRWYyK/Czn/Pjo11vxHjo5l8d+oQTmmrhpWCuNbDsa/k4qpaFcnNk
Bm2F5uae8f3rLO73q3wRkC+fG9iMNW8CMWm/zEiX74+PTz+2Tb6obvGxPJYxTgY00v8TuKs6XS9c
vEPmcbD+HGf5ZCAd4AubBuChkehhde16vAz55BoT8sT7PqaHXFOZJNSHB7XzpqN4/Q/n18jui0fJ
mTB5gBDf4xpjFdmd/vzEpfPJLouWC7zbXaEIbAxfeU7Ix7BZU+vXOc2u/wHFzrnT6u8ShvP260F7
unCJLE0jNy2MuQmmk6W9d4ZDIqOSmBZ+gIG/SI8TReBIK5hxVCNeZO28Cn7LzZBIU7thHACXhWmo
S1C8FHfpevqz5u8DfMb3hk5xmZ/Apo5CNmohZ1isekf1ftF9T1kgtSbPsIArVNRtRZ4D0cBl/iVh
/fSFzpSjRWbAGiIiWeFhgZQ2MIx+DHdADnFUCQiIpLaFVh7/FwQ2P82chusucDtBk6N0hXKWUxms
HSsNuybbRDWMVWFN82o8u+njh3L16pkAzgFcxW2BbhmVxfSNzAnMJNHJhdisx+bLjZDQKqav0kZB
JkEhCRNtTylm5v7QnLD9O1j9Chd4VyP7tKENz47eOe7ZCvnQfN6URm0dGZAg721K9M36emTqzr1O
ecLZIIPTKU7WDnsOmas04cavvwq2pNJNjDxcEOaJXQxcoQ8pETF+Zw44IpKgKqy1EYX8bRgNvSNS
TrOyDwchWDp8Lxs31FAJKbCafhioZjVrB43rbnV6K+PDniZ6Mpqa+Z/nUpDUdHj92wHF2Ue6fy14
HeantXLpwPJ0VNTmgJ9bMZDlFUZhl1Zlp7fmfQu5QgmV+ghSC8P0C8HZ2ukTai0JZfisTcXn9a8Z
Ql/M5QnlUmPQb3k+8YIkvEuu/sixVVfQJtrjUm+f5ysPYmxP2teGMSAbasjO6LDw2sag446MnVes
B7kwlZlkPK653dbTS2Qt996JggRWEipluyYEbtvmPf6Pnv5Fi+0ghhq/Kg1DKZshgpj1pS+ePb37
nYNlyJyu7nLBHxSN4c8hIxfGYBnzI2DxC275RGP4+ISIKbZTiQ9nIzDgni/B7Yz/e+1Ea1PjhxB0
J/JV2ZKnq2Ym8vfyx/JdtaLOCCGmkCLppe/ilxxu+Q2zjoJJrQ17U/QZFzNCBb4PfS/IeoM1i/wI
+cEht+hVYP3UQB+4TTICWbaZdMCb68ZfmIHREd6EEi9h1FwbFUhypi246B+QPGV9Wyg9phvU5wvv
dL4ys/mj42JzkJ+mi6Tena31+0BzxZEcNXzC9Zqol9bcGTYSOr/v+N/ogleqKRkiTZOMDo06/97g
i16Q9y61xDd9hdcyIrOZ/ESBYWpXfbhDcyj+xus5O3MVigpqeq8MS0ZgHkpgS+N8pmgilRKXQIiR
gEESoNGc+AX0kRBPZnnVy1hQFuQjD1ZgIUd5aY0k4zR3Q0DBW4i2PIvjlX50u25fKMz4G6Wxre8h
CDPzfRH+FcZyPuWv06Q8jQuQ/RqmMofXSO1rKOjYmvX2rUX/RHBoLsS7p4k5ukiQQZgxlJTRG/j/
3AbdS/SyBqtR/d5ODK6O+V3DHGC8bhvTDU6RcDXaLeAA7M3CPOow/9ZLI7MWVJ+oDWIhTlE8X+Y9
JPkNcys0uP6yqE6E1NViH/f2UIGj4bbuuToGOG4+yJwdyx64mvqO3s/9FDyIJxZZIwjbejDDdd4r
K+b1Lrx6cMG2325XPV0FqYIZw++Zy4y4REkI1mC2QKwhJpy3nq1yoDZQQB8Gi2poMXwDSq/gzL31
XUDTkX1tqhW+dDbVQ4JF7HWjsfQOsy55B2yB8MRn+mStuT7XeEjeZYbuH3mJNFaTvBGCUeoeNaqi
YeM7XgdiGV1Scy00uiLs9gtDKSZNUe7W5JrcLo6O+fiD64nutGSK1UBGBd31Ri5mUQOSMntUt/5W
1QZdxIiVp1UuyXuhn+Dc4fbsZfb696IGarRCSMvlRj+/4EB0JryquKI6gHIibmYXGPzrIteeSoHx
7n/3Zj0C8EgjjTqD1b8fLgn07H/L3Noa1DaYfIJSTqK4nM38EltyJFMRI5Nm89AnBzMJrgjzQvx7
9qngTZNGqZcwCXAYBKZ+Er6lMOV89S8+CW+MUDOiJR52fx5EDPqDlwP16apkEEo5tXf333QAsP4h
R0xsvX91PnIY4mJxHurejFya+kaB4NKZkrwRgtz9uYVeihsv7gm7meM79KTSQhmkZ/pxSYkCEovp
tXCaYWBX9oO+88+zEwg5P6/+vUACv6j+7phEVoVtn3CD/K0+E0B4mfP+Bi72zteY72La1NWeMbje
HClsi1ImWJuUUK8eF7x3DX1T0pkMriK/oGCSG/1U8KyJojvqHA0TtYXyUCace9fjwH8e8M9/dXy9
0o3jEefh+xQ0pCsU6zE6hticsw/QlyF0xYI+x0BZTMq94OFsB9BzmcH16aDoauVqyWOAxNZNQq5L
rxo3k+fexeebvigSqaFTEy99VKvWPxD8k8T+/vGncve9XDO0B5/fvC9MkC6geVijPL36yjNvLYGC
mzaMD11x5Ih/AQFdUhhUYur432702vXKLt/WCX1NY+Od2HS6U9qGGVHeWTJBbwi4Cog1qNDhkbVS
ZnItNbORn2BEB7OnYQcB82XU6wHM8MFNO842Gpp2TIve38xqsR0yl7iXpLIBHDwMaZfbV63mZ7rv
WVfjTgV/6nuuFiI/6XqX1b5jBqGEdlLsIrLE/m08gvYkVYWGHDHzbi+GA9KUBejisU+L7U2yB1Rq
u7fU+YV15X0jIToA4E2yXQ4pweY1kTr8Cci1wpZnzkHxzT6E0C2JGj8ZzdkRdJjRVZAZnItS2lLV
VZChSiMi/ZTDpEcLNfrgjg424/PS7AUtk61I10K+D9POfFGabLopdzHkfwXOpNYnyRQ4LlUTxsHu
ksnrlGjwLWUEMG55yD1wqb1QmvK5vPGy5XlBdnwbTSTHsamMlNu5cPyjuG0YMEFcO+oPHyvgBuc1
YMYLZKGkFMuwZ+ZZ+oNFngEjIskboujFTXw2CevIWFN0+kYXVaAYgAA+IALNGxo4Plj6A0QLeibD
ZKark8NdXVtV9cMkZ1TswE8F40Qvzl+jQV5CcBOOy1+nzk8KZuVEQ0FtxS0Hxuc92tyx6nVRPhiM
bE0qweTeFRMhvUhp1v34oqMelJv7Zh44EIq4DlQuiTLM7I1+tzkkBqa8iMxeqcot7JhLtC84/6RI
SgS+GySJLE1RoJxO4QM12Wr35HABh+w7td2S3fXI+Df0h9MJ/kUR6WvNXXUUcMwpJEf3nGnVxvsP
+T9aVHGgBbzLDwt0WAI1PUPZsUPu9DXfBF6J172mUhixoNfiXZXjGPr/Dd7lH62N6Y9ALdF66pNF
pdzlt8eICQlWrjszFVvPmo+ogQIbB6n06iM5uBYyYRWLrHH5Xy8wplzdM3dd4Bv9KaOBRh76HURC
YnwZAXwIB1j0RF9a96kP/3Y6sl4YY4oOgN0ltelvFJjPlFfifHUtvZP+I1YVgnJnTsrPXiL3YKxZ
kNIyY2MHpPCFgc06d/86wtstBDtQBFH0UfUXWuH65z72zWsZER6jGHGHBA8WacL71qJ3QGrVWamO
82FKDi7K5JqozfI5ox8Kru+9Ecr8Ebw5zdaSQyqH7Eh/DjjFHdpnwgjjPA+Rd5RRdkeFpAebT/qL
vffP6BUbKKateVRILsA1vj19Kt1MGni1aR6GPRxwNf2441oJNbCFVSYU9Nx4J6TvX6qnUxk414hj
FniLNqrIE+tJYt2X2Wwn7QzMaDZx5AiCRNwFc0gKEHMkA4LGU9ofJfyUg27Cxaf3SNtWzgdNQDY5
mcosXl5YQkK3WZwg6okq99dgHEcfhskqz/9HYfJroFsjzhBbTyc/Caww+lj5h8DoDt6jQdjtYskA
bkM0tu4GCKm6P+GTBMaaq+b+NVKm29GqJrdJLgONJ1AvQGcP0GQgfW1oRpFC/4G/r3BPvdPu3SIn
NUJiVXccAAG0010paXkYHoyAYVbhwzIBVJmMbSZ0KUHQJgnX1EHRsdIZrAmSMimOxb56dXK/fhhu
oMVrdJOGEwR6zHWJEqeE7czFM7SHKhckwj0vGAg5FA/cyp+g2D55qMzmuqFYBeMTsCPvWDAMomvG
9PBoybBIDdQDunqSkaVsP95/Puf9YMeLE9wEq2YrnoHvh8UVvmglLg1EtQR0r85QWmXOhVOTdszy
GuIMV1Z+yis8fxREq0LexTw3VH3DpwBWExrtMzp/KEsqRYFmsg31McFxgsfkzsIl1osx+jGMaPFT
KgsBDfDFRDS4s2hHx8IrmVfCsyBowyXblO0Vflnn29E+/obPNjCOf+gGOoVVlloTDmwL2vuRwqlW
mfdS9VbaA3L9BxegAPFZrEd4cP6VXX8pxJNXuiL6GVrJYdTo1dnAdgX4nCgwmaFPwAjOzo9Ood8X
XpqIjZLbvMNX5QLAYStGbfb9QGCU1epSExHLGPXzU5P4ixchhHl4GLcAL/1ytq7sK+FI+vkAQVXU
pxjTKZzX5f1/4/GXAmxJ4k/A/cubkCzWAF3TGoNqMdmNdKyL7YhXvDLh0ANhC1+oxB+uufOjIm8z
HTHpyYUGkD94phWuT5NFlJMEqb99jixvMSAo976VbGR/FZqHuXgjTdmeCLGRXI2zpow86016RM0O
r3S7ouMKDMUlX+bCCAyjrPULx96FmLTAD56vjM+nyGVzfEigAZZ183q7WKLYvl1EUHHBLWzzfFEO
wpEzogvpaAOdyuoAt84NuJRaipPQvx7zlweFaIqAVtWVcapstW2KO5TbrHPMmT5kDgiK88YQ8oPO
BzYuf5DHiTveqoX9zzw9LDDrqwN2qkbnfnk3qFT8nhLVfIe/gyKhrAxrvI6CiPVpd+AfMeRAVCJz
nWvrJPMjp8O4VQObZDOs9nROFyLstC6lnkllSZh6csGSZFLlqOTfjvqiYmGFwoq+U8/QPpVEcaAe
hCXC8ucmzwqU1guA4GBp9B5K8rsTS/AtCvwhqxHH5USVYHWa0pIgvFhQ0AUmNf/Id2grQ5Gz5mi+
bb5sKGGuot//UDBK0fDlS1KMQM00jlsKI140QIWlUDD31XJUVzck1YTv65HsQAqrv4pjpcZskWur
5Ja+pW1xNTLoHcFLo4ZchDOhlP5yxpUWQBcbDkJsDr0BkKLBjh8aQ5FBz+hVIw/HKcLV1zfH2f4T
AhBW+I3JsLOWy7775sBLkvpAQZT9XfLkFidiIt2KzlHVVhC3hxuWTQlpbPQOJ/jOJCJp/xe3+qIl
XMHDmNFxrq5XEzEbs3MELSOhNXZfxsllzqZXTzmYxoYEkJjYOTJ7sVzjfD0yoLMX2ak544RxAHGm
8FV6Dxxi+vPz1Lm8UVVS4htJQTeHHiB5yaRSPTXpmL7RIjkbfIy9gqqg0liyLGuPoA0sxyqCDoCZ
g9TW+jGSfph6wKVrJFakZ8gk/r8u1932sPvGxkSxy9H8AABrNVGBv+qrTjjg8OsTSb2eJlHk7f6w
GI7JwlYhNQdAIV8veL3AZUktYSiC7F9/f32NA4equ/ywrfxNrHlOn/elwjVqJo73medOWJmiS9DS
+z5Yhy3JlpzlsgUJp18v3rWGqs4rHRmnCkdjIw3Ac/UJRPoySijBZLM+j1M8gsP12jY7VPB3EzFe
VzbRzkQUpO0pDPFSELLWRK0VP3JWOJrtj/sTR9zSAPmzTYInUYKcE/ImvfWuQfv9qhdQrnpBFSZ0
woeGyJLVM1mZR4i3HlCogAytTYis1W+j0Fvf2Pq/DGTvdg1JzgizwSnd0crGD0XnXE+r17/bDkiC
i9o8eHoMRcBAfXTdqr2/VHjXF+SRGzG2Dtq1hqhLL7qH1jVZVtZC3w4Atd2HJe/OCqVsIa1wkm5p
pWmUnK/hrrIlu7veH0671h8B81ABys75I8QNhh5z7zNmGkUEosCZmWSahrbqlNVMQISIMSEhGICu
qsPcD17gRzJ2XWg1d/UhUBUEHp+i4LXaZSVwBrrlUigh57+WnCt0BiWS+t+qlkA0V8ymmy/6F4su
q/8n4fWtyf+5X0tghos5MWwDFLEzUtr3NmgcC5KkS5IfB1chFNEoMgwbEXbMZeIRlUxn+a2eT9BZ
6hc8td2PiqyYX2MmQa4CQF5DUaHMqB0LfA3dVOAGHIfk8Djl5dZ9NKdqxKQplIJUHOe1Fu41N2nN
LSUiyW99tpxEHtVFRxHR6W5O+eHY85xrUp293KxLz61BbcBt+Y8PvQ4uRoly5Uxcj+FpKeu2jEwG
nyutmwOOQOTwLjGH/jOlUdbi4yP5zSeOF/lAvNNSJquExOgpWUeMl+tCCTlypTSgFbEAAqSnT62/
4H8C5C+AncEXN9bM3cTiV3ofRo25DSaNw7gWRBBdCXOCo7sBPnNi6FTdurhKYr7XjVxz7si8Ln2g
Og6elL7xuxqYD9ia1tnbWwnTKpHKdEr6URUsqu75eZfLsI/KHWnT5jomywGoU7GDYuU0wRk6lzCu
ZOXuoFXLmO2eSCeWfF7Qj1iz/YELyf5oVY5xzdgzVTGPrd6JoSe8PXERejqM5YoGIUfInS550+gx
ZOkkV5BazCCbGxfKyzCYZgBoEExMrv5dqg4h1mt2WouSAnB8sBqcAo/JLoiEJ0msCQfi74gq6mWn
BIWHSRL0ygtlsF58gEEF95nbIAebdJ05uW59BDa08OI7Xuv9Os0qRDbdlXYXxIaLuuSU0gQR1CUc
HT1uqg1TYEZreRlGlhwJ14ZFqqksDa5kq87CBHwIiGsqlklHodnvcgj7Ei2tsFPsIDxeNFp5KD+l
TzYoHMwQhRQWybboGVIR4ElqbixukrhtPpKpBbiijF4vUkd4DVwZ+bad9rEh2I8egSPpzX/S+lMQ
eN78Pd8xST4wo9QAXr98iuv6p9U7Rg3M7fMv7ABh5q/BTeoffpHoRqcoWyWlPt7vn4rhJQwt/ucn
of6kuuQHR23p3Wb0D9QJmJ3kKo0SyMkmwf9PbbBrLex+8qEWBf8UAA0zSIAoXOPzOyE74vlncaUq
8hbJXuc7qVC88nhdUfav7UtsAfDXmgXwTxY6hrf6YH6j743In/8abzp4unmJDeNrEAzawmult/Ym
NwdQm803Q97iXpji5+0+StIbSyri+ttOIqvU/hc+VwcFzrGmJ+6Cw4l3gWlZtMm73uatkZV6D7ch
ox+zjpmy96sF7d9UGsHZxyyPyft/2RVSJcstd3/kiwbq99ylHeyeVXkpctCiRLySWxYSNJVc+Oss
xOYPxPELcrL7mE5qahdzZj7rAo+7yYeB05tHnaFRnIDCrMRdkI9Xn4rhRkszfLjrpYKNCdHNhH5t
XbpsrD5+GoAqXhwTTCluT9nZg0OXM0WDGEQGdOrEYrAUxTR6zJ8bNyiZ5i+alVFSAwnag0x1Qaxf
vKtVYjbzi5Ddh3uMTQoCYIP/BQrpOWpew4AQuqU80pQsfuXA7mKPujliLXE/ZYiadPPstFSe6FXl
d4hod0C0t7ixCRHJYXoaQMPJSUAfPg344LzaNajGZDsA1RVP4nClwi+ijo9Gc3Uf7egKLT0QDb2R
kbD4NuF3yPwE1iWQpCjG5H5wewiskd49AQUNdhr1QF+CAy7WYtXw9prlHVpTTatO0mmmqYnNeqnf
w4JTOemoSMEwxmbojwR4Rbe9BIj2Ugk6I1Sevprzhc8gj0xpiMArfnPhnR9SOiYC8guY2u4vOB97
qDYZ6U0eRG7unp6ObHDQzJAYHI7nZDunlc1qMx4jpgLEscafqqHFpnmo8zJ6tF/ikCBBORxxb2Uo
xSCSN5XtSllsvbIx5e1u6bgSWYRQgCAw+8qW+0w/n2vCBgKevkVUB0C2Ks/nJR89BouiCZz/g6Yk
+euSKaswAemYARytUId0bFQ+a2VxH2C2WFA2vKHXCX7CPyubCODhn8Pj5eOR1mR9QtcK4MeuB786
AliMwX3cl90wB2LAFkL8KYU1WrzvIjTxZoTI3rbHrOM2qAv18FVcLXCdZ7u1dl+RSy5mBX4NQ3+h
vEBvJSe4n1MJE+oxYNiq1NG8ywe+6/oLBFFyICf0E3gX0j7Pc0Br4YMjJTVaC+CaIGH1xkGHr6q/
Z1LiKM3m1HeNrFGLkHiq9q2lTpeoujmHJUK1ml5x+ALJOWZyTnoDQOqcFMruR5SIfdf+hgQyEEVd
+cS8YXxW8QKYrnWzXV3XCEPTPx3+XFlm7jBJNLY6iEq9dsGvmpYRkZ10sOSt143O65rZ6/+JnlDT
RQ8DGKrf5qGLthXRQrK4EQno/J8UwQo3A4G+DscRhP5+LraThUHS7N1nts8rkBVsL4MnNRDZQfjj
TTlQDq6ySoHxYf7gIvzJ8DeXJ74AYJ9nY87ULrn4/lhq0Mw0K8981OjuMRiPl7TUZ8FUNoP1Gy2C
NZuZsDTKCg3zMGBzHY6Am5ppXc7MKieKuAU4NbLhA9jqYgmTO6Ar3ZHLUQatX601KZsBF0JzsUGZ
RD30Reh99DjlQYbZY0gHvDy/8wTjN+obkbF9z1GJU1W5cDhJgie9RTsB5H5DUtIWTUmsHz8bL1Bc
7f3HCdUTcRysTq8jruu8Wp+g3tvIwMALmd4tM4UcxroNZvYV2GNtHPhwy8uElB1Jv8K0bhuc8gaV
YEDL89ORtHJI+js6J0SFzM1+S2U+5hNP3Y5n9Gd54/U3kiQ/oWZ++06NQyXrfDXI7UAf6gisucjh
UJA6r0khWYKfEUEBRO9drRo6/yg7t3Q13KK7g+AKktzAqs0rduwCJ0M44B4B7UcZI08ddTe+0uZM
RvO7hE0MUPGAhMJbnzdtxA3BjP/VLa0h2FYoHTDnVECJwPrHFgAGKUf4PETu3Ao9nagbfQXkzStc
XJqk+l9EgbpVuDas5VKBh4uaclccnu5/wx3u1nlm59/a2RfdrNQqYtk0OOAl4uhRux+5RNmO9455
l6o72etXhbZwvCaBWGxt8HO3w+R5pMuUlCEq9aal0QuvLlYSx7SK9o5L4+WgPkv8AvBU+Pn2y+KD
jP6a4mGXk1syJCIuyg/II4/BAJLSSEUM/O2j8xv01lb+/lK3qw6IN3CHeTJ/1m+6ts5O1eUq9olg
EnYWjRj5ReHlahQpugyAuFFPHQaoZZDmpV0W4jwGMZ3tIsTV0iASGE9E8AOPp256QPaUAWrIYfqS
0/AffVC+FFv7bWQso6l76blrSM+lVkitG/9lhZ5SKbHhi3xQW/Lx2BBytvZd90cGa+FCQBScjL7B
UJG7bPsID4pgWt0eCu8bRIIsCHxVBYY0vztZTNuaMn4+clWYcguG5KpFU0FJ1jC9YiUhHoqBTjd9
i5rKex8LoVHx0oTiq05zuSVA2V0VNfl12YCZFGRPXKKcnlmefMQuelPgX1JXlJw3YvZwu6Ph9LRP
HTzeSe/vcYF7F+L9/2mtG7w+4uGHUYeCd2z0JkI44gCE1ZFJ2nWpdR1U+OsicYYryZVzenKGyxFh
IjIV5zbvxZ/8bpD/+7fIxie6kHRQu0QfrQKbCo5NUvHkK7cZ7IzCyx3NQ2JBBCkTaezP2tHZKqmE
hsBJT4Oe0JXvWwzFssWjmE4gcfJ6BvI5L5a5+m3CVLUFhrUFDm1VbstIaGo2dmAobtJIkvTdishG
8SuqZNkQQDJFTYaZysvwoVVfy11iXiCdpgZAonODfCAJowa1qUVXQfl9vhDg4eaH7eDT7BOHfe2+
FTHZhE/odnBp8zmhxMEvuQD9TrhPh+kkw8YbWXX6IbcK9idl+DsAJmj6F6ahVIacIv6vh+dcQJqo
upUSn91C4zSAKXLQOpECTLNKZ8EKlMgSedK/WYokiUdiM8b1cFAWbyuQoeu9hARhPWmZ/iSXXiUT
XbgpbbB1XB6SNpMdsA3siMWooQcxL5ik7h3O8F0WVUCGGK3AstP5f+MpMQxyIVlhRhFyDuFsL1xh
unKspbq8KEVJVb9OrtArAaobNHekKoMu8DvpGMRiTye8gCkbgQLjOQNjLqWQLuBz7s6D+aw7FXjM
V/eKAtbI0LFFnoLxFjfia+DM9BOJtzfx+7RBqD52l+nc2RC4yTN66JVFimQnVLh7xsCw96zx2IZJ
EFnqt0F99/9rOVvzCIky6hYR2d9AfBGfEse7Xn4wDZT4p8FUCWsC1Mk9rMyjUEgFgKM7IPMfERnj
t5hO9SxtvQEOtsjw58/A8+H2iJjmHrmq8brNB8Kr6OdTfq5EsI4dAl+Pr+f8ux7H74EieqabAuaU
RHotDsbB7fstPahfta0Fb6MX/oMKRDf6C3s4VTFvZ3eo4QP09BzMVAlVnenpbatby6pMU1u9XjeI
kE4nqHAtJNDUbjZL8Qzij5zZ5k1G5tX0V0nmRerPniCGYfgD5EuesC/ApyLbV2U0e9959AwcKjLL
OVigRYSAJG0cRFuosPXITXRzPBUaMVIut3l8TUb/Tsx4NQIB8qtf+K0QnX1ho0cw9IyS6vOehekH
Jrl4CZiqQCW+GAPAZQkoJY2kBBxsmpRf2L56ydsLxnuwfEKwvuf+vmuapVhPwMlQQE3gvuiJp/e+
zckmd3bREDeSVIRqXQlKhKea6uX9zSEvhs7qbq7W+0DmpHD/t+iOjsUFqvsbq/h87K7oPyVK8QyE
HIWK5UyvFdSYiLsWS+yJv0fBLVz7Z+/FO7PRDRa8MN0rgYHRO02iMYhNSCrLJGn77mVjr2xtdVRl
12UyYrB794GREKdLl3ds9bJjdafNxRWBuYefTjNd1HTHbs1LbJntUkSX4XO1H6XMmcaznt/Hevhe
/PKzL1DJTjvwdCIEJFSkrIEwoOfU4NjsHptmSLERe7mZD4gVTHKv+MRQa8cnzFTGpLsWm0YMri6C
+hTB2+BMmogfSYrBtXe8erwGRbbz6uo8Gi1PO0A07BjafH/eSPlGxOobX6bwZem4NfDEr3ewjYBh
9xr9y93LudMXPW1YNDQVfWEQMzUOWoRVwalY+iSdSbRMkJy+hX2OvGVnAIjLycUuwE6EGdIq7vJ/
5sSHnjiFrv2tkjfcGiW54/zfL70/TgtHmxJJN3wDRZ2GXNeofFIlltIvMcppT0plbx3hRW4Fu8OW
Y9+JC9Atdml7JaNSA9+hIo55ZluwRcSIVYUQdo1GXqN7sO2NnQHa6IBfZzMVnvl0aFhrs3Wo8JMx
gB1H9ZcIzPsK0CCCJfn3Xvt8bn3KV9oDk5rMe8WmUM7/N6m5sbdF+ewXrut5iUdQSPt91SuRRhBU
9AB8ay864juTpNUrEwC0XsnAHW0XrG6ZP9L93B1pb2oHvyfZ3PUFdq59JdeDE7+jBgX820V62nws
PZ3OZ7uhLEFC4vbcmRDGR4d3epVr9iGUinS6rNoTWdhANZvxG4V5npvg2YnYuOTRI1fiknz0oReX
gJaFmbJCvkjN7uxEWi3h8hfkkY7Nziq+496o1wnTnJNG2nHVHYS3hJ+/l35PSKOlEtdL0MJe0wkf
lWym1ebnFCa7hH2NTYN0M9wH9CYs7TEph78xWVC1fDWSw6pj0vXrsfr22fI+fj8Yi0OkonCr5BeM
7vPRT3h4vBOKgxVgKKMZtdlrwMstXyXDBEcgC0SDb+6Zjz3mXVSS69BnoB/RDDpzJnLs5/H9KH0m
ETxovx3S6Irk/sm4SrbQAnXsF2mMrzTyUcJUgLiRxJEaRvvEmNZ/jlNfuyXb81rYR4lHtVDkLU7u
cJZPXxY8h0LyLw2xzheKhxDpG3sHUgSjbh3Qb7AQOd9RsQOpXfWIkK/L1gI/m6h4xze5dBqBanch
HGj0VXG7elelPrqm8onPOpplAMI9eudM9HjPfSI31bU8lPFIM86YABZ6+TikTeL3zQ2rJPi6lXKK
EISm/2WGmvNTDW3UlH112bViBjdIrqOkhmLO97zRRfWwd1GZI6ows2bk1x9zLpqdjvoBKlutNMLo
0EnFQE84HArjzxN0VidCjkIfZxjJUAe94f9t8DODBxzZWoSz37kdi0ch7yvCOapUoD1lZtdlxwSu
AmpyyL4PS4NSizNZpTCmlq+TaRT5i/MZOZbdjiURPXMAQfSIGbfF2slZ83BsDaHfwFWSMMuQ8ESq
29J3Mvls3BxO6u4WYS20659lCuWTMU8hqT/PQviYbJvE8475v9wl1xqrlGXtj+hfNgpHfaoXv2/O
ubbV+dlOP0+EEjcX4/MviWk4Tla123oqsWrZPRwexIISZMkbzUl6t/XwOsnSSgQACx/Tia11AkFe
k5963RcATS/nolC5Hl28arUuO4CYBKwr5ik/2HdIzvuFfmuLA7vamUJf7gXGCU+ny97pwLAKjOvw
VQ+TvneJlMH7vG2uaDezvP+csMKbmBVwKRDVkMnzpQAUjOewx7ob/aG4z6IR7o5c6ysDMteR7ioX
+idELDJBni4HLg9gJ8gCd+w2RLXRfgRjnZZ7LJKhuSA5kiftUhz5pO241DRtJe3hvlB+Cs2JUqrs
1O0GlYBHteMPrJJnfHvcECqZlrUcfK+4jBUmxpcWCY+1OBHCk3Isuh/B9QZ1jzmJ8pEJCNXY9Iw1
w3ElOzFV79/Ect3aJo7LC/6NQqU5d6SPNk5ZFN1c4KUYhF69ISi9+J0wOIMDDN9r0g0oRFYPpWQu
veDB0HA70eAGW36k4g1rbH6VZIvD/0MGIiI9RU5KudOhi/I1z+4c/Fnzq3etFW6jRb7CH1j4ALYX
MlKibVBcVaTX85JFeSPLTwF3qRMqrXebr/C+vlPEljiZ6u9lO1r0Z1T+lMlFH9NhVq1U+bFd7KDM
oGNOHy1w1pK7SX4VX8aGTb48WF+WgW7NFUEaa0UjJpQxvr2sxbmvAEz9SrcCOSJjzyVizV7+2oV6
rfFOnu0rbC/Jz/mszf6up4McuUnl7RIiSdvib48bFmx8FFldk1zS5PNHD/9exHdIfR0ZBDhnO6X6
oryG/ZL5r8x2tAZTRq0dD1/U2qDmTu3vvbfEeN+i/7kQNu663UCfoVq6ijtOT+2EJtTN2NPuRK06
6o3qRF40Oep5GZgmaIzpa5bv7XNSL6115kUuzACAghF2pGBH3+eVeRcznwJXd3VTrIopS6LEnYNu
ebAL4UbKI8Tkd56tGvH8QK7BNjN2TyJs+8oOzd3uJbnWafEmXXKTmBRiXAylTrtIrVMTCMkcsZx8
6SaUyaq7/Um24ambK0mZhOaVn7NA6VAMg/OO9sKRvVJzNbJzavhPA6Y9+m5uX6SO98j5kpw8QL/l
vMp6FDyAJ6ejhTmyOs65oD4hyGue2lCOa549/XjtdLZDsSYqNDWRi1fPPL6Pu8uLK3Sqbt0PPWE8
360BdDkYIkavmC7sgqEQAA4tRT3I90Z20/fyqCedolytfWXl8Twixzr7vdTTXLYgGWBv0aQnYPx9
JifIvSihXyUD3xuM7vFOF4vIio8QkEPCVOi/ATbxyIB9gx0gfmpf0ToKReQc2Fnb9/NPZCP1UZg+
c9SYTgQoakH1pP+JgAdztu3LSHKAeqZdniCmXYY8xqVgI7+qdEZ3+R0BDn6tJaI/b8Wj0V2A9hjt
i1RISKXm1eW2slV1TvJEC/fbg90oc3yn6avhff44bEKMG2SBkBVZKk6e8LxlN8R24blY3SOZQZ+q
M9jdGPo+l043WbYvwuc0cRoQg0PRcdQpXNRPgSgqUcy9DtbaA6fPf+Tfh/7zm4JvX/H1uoMv3O6Q
30yBvGLKK6XQGxKkl1etbardhvUIQluD+IWJpqYZrzuuB3NUoXpodQvWXSaJY3qx8JoStRJmBa2t
0uVJ3Fl3rK9sKlHOMcIAF7To5AyB2CDntWA+RRAINgImyBNYyWSWU0/sLGjn5rHhDcbktjG5gKYQ
o3KWChrxDoJk/PRU3oXxCxhWC5RJDJS4vT5aAkwSEfrwwZf/EAjCfDoY9x7qCw93i/pxqWE+mWKO
BHvv2ujVuFdzWDT9vDVeHeA2KpGm+C34QfaaRzDjLFaNhkiS0VlnXe8VBaHjM9SccAMFEX6SOFD/
nJVBXwmVANmjnU0KSw4sJ+Mo1nJdvYlR4jhwrDDXm4PvoqtoEHNTb3TdA02b3j7NuKm0Pk7fjjhK
5ln1vtiJN/BQAB7DpvMVPl2R2tu3TaptN4dM+p027b2HSJedrbVneEyM/41bvM8j3NGMP3QkZimE
L5oZf55jWhmjhFmIOzQ6hirXmXIWTyVxlUNHS1RNQhc9xPc2VeNKbnhirFKU1znytoKIR1+zm88W
CgzMrwv7fNMK/hbu7TaU4O1HaJ5jCONWtgmWJPCNRr6Ryqy9j4tpVua3bjq2c4JeNraylMahcgEk
k4JNOTO/TsnououAlhIU9DLPBFdMgwfGgoLwgthjN5i7D0OW/TMh4Tzl9yOM0wOt9EhcH6qMMc9P
KzO+ddJZsjRUxB8swyETo6E6yewAB5xspRV2dlQPP9g0/HtTfFHWA4rQbyglDbPi/VSqKc0K9/E/
PdVzZZiea8Ln0CjjDweYkoZs072YtoEcIqVNuhKV2UQPCXs2StpIxNCSMQjdcT03r6WjDqCH5vyZ
zqJjCLy6VeG2X+unqeKuQ6KZHtywAdrLcCY78QZ2D+yDWHOxOvr4iV53qNwSCSrz+yw90QqKBXFf
uSylkK3TntaOqGGqSoprwhJnOcA9n/+GOcQBqOKqAAJeZ2RPeY+fTQfEiTn11Nr86yib2Duq18Yd
SVMP41ERxuNMskQaT8kdfN3V5iVvf63LIYJsr6XdbM1JCHhpTrbA+tAOcAFWhUO+zYxRJNjgaaae
ggoavvhS6p3F8jLRM4DSlRR/kYwkTOLkuGYPUjlaNy/iwUaeo3EP97s+/iAFs0MGJFE6wscdXj9o
EAaCIFNSWLCq7xqNrCnqFyXBt07NrfnwNXUyTNeX4A8TAJkpwXYpAN4xtzxkM28ynXmAN5w5X/5A
9ApNnMitPMCs+SG3jZTRH7s7Z7bfGfbEoQz3RykhyNSkU22YRLbJ+NoovhSxjlI7tmYaXnkxChSx
v1NewAfiWBqTp8yAZnKeIQfTs3f71ywA3WmQ6EmzQOhWHPr6epUAjHzhhcxeord+t2d+XHY7867h
F8fCfX1Ow/g3y+1/nDnw9vxgHlUpb+6CiJxPMHtu1iZcnWRyrMKx15ggx8MScxt+TtGqMaXrGTHW
17AkgOI6NVyq3oINTh0JCl3DJC4DuLCsTAYpbFpiIE44X7zUf/Gj+BJMVchvPLMjckoVkjBMnfrt
cLZEF4ViWSHHcUQjcrrz31+2LQLagr4F4EN59SvclF270JOgY4/kXYLEKJr8vYC7Hu75yKYpd2Ph
jsa+T5uEGKR43xqCiiLCkiOl9eu/+OfdtujszZyxS/RquzxeiwCITo160YBIf6DfbIlZ3sJuMaEk
edb1Zqs0f77yO+D38xrpB8v6WYAQCbm6T0IwWaHA8OcAm2aUCCIaEF1/Bqb6QjOTt1ymcVKhmBKW
O5U03VhBlWUza1X8R7GdSjaBXm5eLFRNNTsF/DTeHmVLZ8Yb7nmmFaVO7LXy/djGQMq4YYXnzdUt
T6EoV2S9v0JI2+WvK0+j7e+yFb0MXIknzPZe3tCuV17PRck1yKtIBm4vTlit7ZxlbWjGEGWkRMiN
8+ozsV8Sg4ucp29rB8AlWcw46DJKR5Y5RY5Vl7qGphUx/myhvNO8tLvZVJdmrLupwEf9JN0Ndr53
ehvybY188jaGkPoz/ynWrDqD9QLnR1AHmiegubj++jzOqiwyMhRMJNM77LJvgTnluiqHlGcdcejz
fL9OrF1NC1wmAJ3rYsmzVVse+poxuj5q98+TtQl4Cp+xN2Wa9CAYdyqSCvcz3N33JAzjnIovA2kp
pPYiIf2dOzBJ9BsihRuKZiJwySJTNj9oJzGbE9kMs5xHG9dCe76ULPl/QZYKpHyfizCfbHHl22QJ
kJwdxjdMdj4jAG1WPmsR/iykOhYIUgTEnxrQR9y5xeAspaqAAaun72whGcFa5N1GOKkbFYsKX4Aj
hgRGdTuOoikR879ndnJcqAQLWphqtlHXnH8bYqCce2bmtil3GMoV5+3hUzSnB1VtxX46F3KZ267m
iWSBrmOicFDZm1qOWROw6Sg9WnHJYq9MRRMDhlBq1KmS+cE9G8YUKclL50TMp0gInVW/d7JbzYby
ZKzNYMrap+Bsn6yyqGrkSieGj66itlqJG0LFOn3eeAYBAUvOuwdBU5SEYte91FH74lM8L3yx2Scy
0kqtD0l/fCuqWVqrGSJf15fnV8Oian/ZqPNxdr53TulkpISFfy8tHNYp/nB4CM1V5TfoNt01GGJX
BBnHYyPWFGOCKLyqEq+w4t93UWhI/FvjHn86h+JetBn9QnyrGM4+rbz2rbN1ai+Xg1XlHdeCvLHH
+H+6n+zXWghT0NbJ+UUXp4xqUflFegLmmzr2/11zhQSjzktu/lWT4LpsvULcQxWAXYxfNf/kCNUh
Qn/T94I0ltHNRok52/rA5RpXYpSWvANNHzrabgjhf9UwYaBHK1ok4bG9Alg4ahz7SkrQy4jD6Y2w
QXSk+qL007WUGGd1LqgntLr1/JCCfxnsh2HWuSZUadkMd7osbZMKZ+/5FZfdYMH3A6y76GROjNJh
LON4f1KyqqqwX+n02KDtROjBVqU6zK7hcHv/LqcxFOE0gNxkp5x3iSQ0DfEeq+s90zH4DlZ1cLJU
Cg5LLlS1vDpBokB0LXOO6uEDy2TilCmrAzPAoSSdRpF+0b0RL39Bprr4bRbFXHFsibFiMDuVlU7P
eIm34O1anVTkqMBzGSYlK73yazob5d2lAap9w3htF2/qJfbJ/I4JjWfSGC6lYyiq8E5/W5PyilaK
33oxJfQEIWu5G/u7ZscBeunhTo65rSAQj0Mm4zZUv4ycJJ0IZ04Z6WA65N+kSDCnkfiGMxyk3mTU
Wq7CLeJJqUhz7dJiOZ2wwrROUWX+CkhDPCPLnQoQuijTF3SDReL1LtCs3Y3KRP3FI1CrsIBeuqoN
eJRC23w3aU9T3BRrr2Mo6DlGxi31sElmHqKZoM/J4IXRz9sAuY2LgVGxrjIT7sfqqYUu7K5VCjKY
PIE60qczKdjbmuz8zo4Xks+spmCi7QMipIyefFxgYlG3obvUDR3gOOCBoOuY4AvM7nnemTCH9UW0
W9SHTqAuLEJoZYr5mkVui7zx475KDk9EeTcUwZRqOoX81YwBly38xvI+8v5cX9QTbvVR7SXLtNt/
c7M0+WBxf0N+fYfS67/IxMo3vmPjNc+HLoDhc34YX24xKbDPW55DrRvi1uasbDgQgCLRx0mafh+L
87vCUyiLRFKBlmdrSDZcHobGC6DeUarWWAM483dmajR+QyeYEwWcTfnpvN67a+70+0ixldtjYSVv
jC978h1Zq0pCldU1PBHar/OJIiwCROXyH7PHZC1F5IeUbScbxAcW7kAZRNdy/b4Oq400yQ1+Qib/
90+RSwtw4868OOu8iK50F/cDzGl3R0qMJ0BArGpRIMhIWkP0wkUHBng0msdT14RLllPnv9FzOAEu
xW2xN/l4dn8/KqdGqRUEcAEubSahA8j5JGjq75+Q26A5WbAC1vZrO+ERF2TKFbjlpRlp1dYm4eH+
9akG/sprJU1vCzdl+erTXgEIizoeFcaoFdM2LDr/0qQ7k03NeLSADL6iY+JwSmlg4DYZDrncdYxr
IXsbWjyr/hUYJ+oegQfiPkSGvJY4N1KfeHbNoElmq7ILh2wYYmObPStJtXfj7zoWCd/UmbaNtxrg
SHaMSRvvCm1pK1RyUdoSwq/orjsBxPGunOsiDlCrp0mJFkOBm5anR4wLFk6i7he7QCw03VGBbnpZ
un0zieIC5BBTGT9zdu9Pv+8sVFZgl93VsDPIkaPC8TO+diFyCJKX3zQBoXXJKXPeCdsyNbkxyRaB
Ak4Tl8FdWw39WkhCldRi02DDckbK2+DfrU/iPECGklIzxy+gco/VSJoDylEUe3m7Hg5lyv1EDliH
nqRif+Q4lfAdgXPZ3tSLi0n4kawRydQW19jowgoxjZm/f4CuVne3f1qrakbvf6SkHDZSiDnDxpQ4
1YFJJeBRhcoBMZ6uH5t2RmO2q925NWHE09gO9DRYpgcs+KKDHSGIy07YUSMjNnVDcScBVYtMBl1H
N3sPuZrEezEkYYdI1VLibx4/X+bavn9QvI7MnyQ3MrmaxmKma9Fdk6r+SU4LBD+YYf8esLg+D1Sg
JP6c5VIsGUjZV54Fuz5H1Xtvw/puN8eWBLRLUVPG/859gnp//tg4EYBaQUBF3Km4X4E4uWIETkqr
fFr4zdwy0bva/2ieRq8vAscM2eRtJG4hcjMFQy1IG3RVKAwx0FMVihnlpBRpwdDaQHq39vw47BIV
fiSscMRd3czsMAMBXXXPP+W/7Q5o2RugSwBaREturKvU3INNAGqC6RV6qMtHJyF81lgUKp4qc1//
naH3uLG3u+IaAQJt1npN+I7IOBSFuYLUpAe27XZsD6ko1lG23QsmG0wRKbbR40V576+hrRDMjcvt
WzF7fSYMXaZoX6t9R1KhBsrz93GHDo4FEJs+HTSHAei1PW6dRNMZ0NYv1lElszDo7oK3r6fgbSRk
wPpBTR8RjGJnlCZyZR+l8/F1JP+h4Uoxj4EzP4l3KALIbNnkEM+3dNrSxK2aZqSwT43lHowMSErh
QO3pntQ+wT9WFRn+vPvZWN4PQ+EA1Y2UK0h/czY64rcrRYKO2RuRPmiF8yW6J7xwxA8tW1PeZ5dD
QWd6VrBUy49uAOtN0zMsCNLsOJYLYKcXJfCjiGZ/nkfGDOzQfmzbtGcSiUmMVrIP6nTXSbHIeiM1
Yxfkk78JzhQTYTYfzifnZeicx6BZuWqHtJfNEPOpqycb6CEwe7ex0voR5moAZVoasc2ttjVhrOA0
6ZUUlbjY9ZyVgKjLrXST9nz/6R5sT5hVwEKyfJyE9mYp7cZ/GRPsfTjxhkRIz6tw8gQcnw5JwDPV
B2yiYZESrBPcchWWappapxoDQGiWu6SMj0tTZT9g2SP0R4s5HupGHvr8Dv/of5unzWE17XCrHhZV
5bApsv9AczLtEWZGXB/BKtom/f0MUGZKRj3wtOFQ+b/ZLySg2rfQT7aA7TArqtfMnuTocHbFoJ2b
mNXnFPCcYS/5p7x+g+2PJzC1mbbAkGRVB741SV40ioYV8c79KUIi21IbPOWmnlJy9W9PorxZX3w5
EQjsxCZadG1U76HHh9lDlaoDrx6E9VY749+ixrEmQrNmGelCsBL+Y1/ePBHVmFm6Nvt7XXK+Y1oo
3oRxeLfA3AL5gnYpDhgVvKOrR++9tr0wrnwD66kcu0xfyXyW+vg6IMjejB3+CR9if6s2F/sc/5wg
p4bDQjJYkcdKkJtDOQv48mBDRLRgFB5BUlPxJR2ldNiDQx4w/CjJTEc+fSOnQRzEZGvdI8/CzOvr
YZY7sH+gjkBV5ezeCnISj9InImDzroGhQCf5DPd8TrSozEmBPuiemeojmFWQR5eA9gmHKNOW2Oo/
Hr9f90snCO9yFsr/pV7QBy/BSkiAr5sk98IWon28eDQZqsyII3z6igVfn7nvo43GzfBD/wU8229N
kKIuf5GR2G7DXWVYiBeQscr6C3525iBXFw/+38cmgtL1WHDdqisbXW+V8kevaZldztL87BybTZbJ
HvXNP0SOIFP67mM7feXAjjOZbp06X7jCeedxE03KIm78Z2KCSYthP3HcAe9PgWduWOUmuUoHbHTj
8nexHBzd4JwBk/1DfpsAr3MBwapJ7NDlXmmWuYg71s3D6o4T4qKo2eSncnlfC4eh4UEudO3yQ6iN
FHLZs0dzc/wo1ssOj20zYNU3qP4pDaLdj5vrXBm9huC3Gvj5rrmbyqmNJqqS6Zt7fULd79FmwumH
hgHxfIIBU0jSQ7w5+cFPNHGMsdCDCgi6XUsFg7NzQlHslv02N1OvLmdNCOLF+pPz6GKHmOLSLcLd
ch8itkOpnOT3o5LAjoW/+mzvA0Btz/+prTHVz5V8Qty3mrfBymU9IJOO2WVofZARflUOtAWZx+xt
c0PtRt1XsVjDbxn6W8p9ZMbpJbCKc108WhXm7NUtgP6OJldKVZxk9DOCOFhX1fyzv6buZQ0gBRnq
h2bHjzqD26aCXJBkJmn5oSYsnIk/6R6RQUaw+QZ+GVDDN8O2mD9dO2tfmRZ9Xq/hMhehX0mE4rE8
b2Ot7KEllkPu5T/tyKMM0e8E2rA7fOnaOmkpCzCe+qW/6rRCpPRR0iCJvZpHpq/KHLiFoXmNnLNa
ayD3yfOwWQ6faHTQSpKOMCe1mE2djWNZGLNsah/cvsFwl2vQ9DbqE/84fsHvr3BFRMKOruncVzfX
SFAbil5qLIDFbhz/iopnFdQeIuwJ/cxuwxE1xf6zpHICSpuP7RsasltDNB/Wc9PufCtDLXenljmp
yAFLVMM9JXivadQNRcnLd363WEVjdSrQ123/q1SFmX5g96581TPwaZDnUtfTj0SKSfFKMkczNY96
kYsqJCtb69TjMR51WDGZzZ2G91lqviYi7VqwnmsP5rjOa+BHAUQhgyKBEoiXZVLZBHWrRJC2oFD+
gRNm9khjcg4aV8jvNkK9GvMkEx8Sl5GLFMR+Alfk+9x/5y3TaS/vaHRy2wMv3uH0TPgcHpwUbXLq
yLCJpnHq71ykHWsRV/INmUA+hU8IFXmMx7MD1vsUtJ9161uyCDB+fHP7R6NLL5QqbEBtoUH9kxZn
1HAgqsjP0qeJjV1eSIV1C4FWM1NFoHU9y2y4wyjG6o5VxKmMuP5CpNxTdVc8WejDOhcx6j4KQtYQ
9+3NGIxQX8IAZVjJgI/63Tn4RucyIirx4fixXTuR2kbYgiGa/GVhB04NUYWLxl7fQofFckDnAdK2
tYQxiMr+THmzY0Gbgv0QElQo2hWPyeYc55ND9eSadEvZUoRTzs2ot0qXzKCpCqsVMiDRZqQy4zHI
PkhjG/hB2lsZOyh2zl4Te1dUgOs70MX3r4SOSuWndQFWIG81KYH6t26KBjOzTuVcQjkoJFJB5Pcc
sadMy1TIiJqcb/MAKbWhqF+OgnuxM4OF8jlmIzdz5bF62On3xosrJtstqNu8AujyhZs51k5lV1Xo
n/UCMsFzbPikKnihvGgKCFM/IhnhIR0xt+2w92V4T3MBcP4AEt2VpuxlR5tyhtqelTdaTuHhqJ86
GB/+hl8NDyKUGevKIoqJU50dWT/u48duj6vWgfVfq1+7ODqVHoVnx/x83zmckrSZFr0n5H5y1SgX
0DgKjrQLFRT7B+u7hmbXUB+UF1qoHXzLmxKSOUMgyT5XuAp3mhc//oxfpdzWihn6aSL24S/1t04/
JMn7Taos/PDb8g3qMkS0om7UtagNLCqlhRah6+Nc7Sc6yz2xKoYK6OQVN61CEREk0cGt1R/y2zZ7
KI9++WEVCFjc/vNg+E7/bsnQ+YF10t3gFFdPIIn4LP+BKmp2wihBAUa9zEOyRHXz4pkwWObWT1F7
HfeUXG1sQwnPblcyy3wS+SqK2M9JX/HkhaMlsJ8w+QrATcwFLFoxkgLRTQP+LnP9yXnjhZBpZKZw
g081JgespjztEzNO/3CajDSRRIgNeRjR0lkBaRRQGs7Udqur8SKC85kySTafTHAPKEKipcbx7wAO
j5DOlLi1+ZVSbOvu81WcuaYfK5xR7KaWpVqfCwkWYQRiRDZnXOHl6LjEzr8/aj9Yb8aUBOQuKjGy
bZtQQ0PowKxnKfu6cbefjWex5ZnHbMBijOUku6fD9zAOXXcm7FzDPZmF/bWwKGAMnHf8rh7Fsvtt
QAS8oclunuXEYtJK9nrH221A9Mp+ZSQotj4lhoJQ5Uo5YpmEYJomi/jUGzwLowJdVDOP+ihTdxYE
e5mRA1sRttuoO1xPhZPTApy6YrdcJcany9rRJrns2zSVQTyClKobBK7L3n1M4YshGIGsKNhd6wYG
/NFhlOofs9uGlCBThdz7TNdCVgo2rNi67ZJE7cP24r0MieTm2KcEqLxxEdbs4y+3x3mu4umNtBsr
nlEWCuz9i95lTntIaHKmHLtQVR2op9TtqswIYia5I1R9vmenG2xvYrG50PUAEj9URb1PVEWw/q5/
e9q2hMHFwK7aGHMYQ7iv9wNre8Hv1s0TVM2CdOY3eO0IguFd+xv16PCYaFLz8eQuAhvJUNwsILaX
n/bm+iKsjsyEaFFew5mBDEK7nlNncew8dQ+Fta8DshIFmwZkkm2cJCZ5QqYm9fg4sEla+OkSdsFK
PYc/uSuRJwgS20gz1HNJM97vEy31gfGaTJwVKSAzvqsXWhRnguE4IPMUK2DRwoFAxYRdubkKCVtm
e1cdldYWPOQOeyNKCf2Ql+THYHfKdbJcOOrjFJcpQu0352RPJd4QCRd3SnC74V+Kmtg3VCEGTCch
yANjNq6IUJhPJgARq9V5FSADOMiiNRXDiaugNJWdec2MaeCJoxfhNkI0QQfZmEj1vkRyFNQtFG+f
DcJPHFHytGbLNwpIMUIb2AbuMI9YeOSzm+c0qVmMRgXhAE8q0BE4hOpr7O3tyn23rn3+8HdImAej
KCvm9pxr7CMaoK11uyWY38l11i0+7ZvTRcaDcwaN4b2nVAbjt7sHhyPIeKJ2QsPVyQUIoPB03PdD
PPdFWyYKi839jVUJGImbTfabSTQx9ZItzo2Rf+/Vb9i3OM3W1uq2fqKtzdX7SNKYPl5AdQ9pN6Jc
0J5dfjFnIhcMfFrt6Igz2S5oFwm/EnvxpnAugukTtbsILX6PSsmOlG3ZEVNty9JElu6m8+cqzEWJ
c4vlMWE3q5KXE3TmQJ9HFYvFm9JjVpIdGoaKhnYXdcHoSAptG/zpQ2RVTuJa3VYKtsLqLdDoZ/+m
KCCnwT1R2+xdw1ElbIGDNzMLYwkwDM1pkNslIRRFazakttRMppTbhP3zJkqfccOxvIkNMw9NE9Yu
b385brucZXc2YRNtB7Xj4awxJg4dULT/7XSDI+2ZSz0zE91FLjAuYlJ4Aat5hFBQrLximTemUn8b
LwUkbMPuZsRiE2YLAWMSSxXg2sSuA/vAE+JHtNFtA08q5mraZFkAEp5XksieWYz4eWyTI5htK93U
4prmv8XxcjiySdpbpagyybrOAt4odKGdflA/d+6/w3cLheGYfpaFpff5JyyG8V0GVSebs+wv84w2
2B1h8xeLBiBF3txNWiy7+1isEQLsc2J7vActVMPxOnvKsvuK8bRrK62cFWhQu6/e3Pt6j9ySAX/P
iF15Ep0QkQdFtxvGLowv9esOgepTG5vU4TAhjDy3qk/XEYBAvA0JY8DbTcFXdZ/bXz0U36pUqPed
t5pfbuk931TNEzysoFBMoQeckH6r+N57MZGXuDfhDmc9H1Y0h0FBP8T/tNuWzyD2KFa6kL5k3zJ/
DXXZFFPMiKcbbKjHCNE4KGr4n/GkOXB34zJN2Z227FeJ+rKPd9DcjoeLHPXOK/UyE0qq+51ZxAin
0L/xfIrK9uDelRg9dctYSvpC19tPhD1tCIV317GdwvFKYOixdEcay0GHu3ostf9/KGNwxo6ztpD9
SWplxiqU9qiWr7YCykjBUqNnpsOAADOFn0vJLNcaOeEdsvm2aI73xXC2eYI6txdDn2wDRUy3IiFO
EfTuqm/WM1LrW1HORusv1kKDjGdzoZGY0Ym7MwHL/q6yaMRNi64OrlCCrR0rtIorzRJKDbaQOmTR
S2/dTVYfDgUYWmraT9uW1xYLFTN3ni1/Bv4pAwqpsHB3aXagOZYJB5DXPUC1kq22S3ZmWNgATa3G
RHevl1Y88MijNgweQ8+5XSsWWVkTtP8Eb4KRYi72Nr363cBa0nBLtZ/BXKrlQ+5ZO2BsJxy9ky1K
ZdpAdXnX9ip1JJal+d+w6zksKFTzEuTqDRHNrB5d016vo6yDr22WmJUOgtNuNZtSXY5diwNMGlks
L2yFgnrB8oVFZ4SJaXl9Xhh42uAvpHqFuj2t6nexXeG+HzpDp/XlppKXs+kPxJTf3UojU5MNssqW
1fQuzYiq+hWb/y4St4vCv5vDvUJlWA/+Z6EaHo9FGWrm3HQaPnnwAIGVEE2C3dxwbGdD2GxNwK6c
Ij0eH6zlj3k4FN7PIhBfbaviHPB8wipv0DoD7dL2dWblMkDbu4L0bObLaYSUuIoQ6uS7CaRcYqEe
ZcKTeO94eXrd05dz2WZA15Ecn8GIMJe2Dzybiu61i9K2AOtXqNyGd6CQBHMveMawVhqMQvYtmgN/
gRJP9+Tqa9vVmUKdLMSfPZ4UG9Mt2SVof9AfribRMLlWtuM0pHorz1mXbStSqQ14UkBxe7KNWCE1
y1Rxa4VMptic3RBzkWF8Tha4oXswR86sXQ3Nh+IbiVqe728CcCnSL5kfe8Cd1Sf05++tHFQmVdir
mWoTWoWBsEfi/rJqeFOZ4kh4yPDzy0qgquhyGFreUSV1xKwDXEF2ZPBtrKAynnbAXYwvp1fu09bv
V+/DrMifI21616mRM1p76eO8kBVjKMebRaXj03vhWpTRzY8dRnYF7aYG1k0xJ62fJKlUCpAdvfvj
K+ULyd3fwPTggt5IxKh2MO/kfxLsYcgsZDRsH8MzT7vr2oKe5vul6jYWs4JDs+tbM3xxxQrE4d3w
OOfhQfPoMWwb+ZGNS1iApSQobR5239cTsrWP+q54939fI6Cb9QduYmvRrEy2eTkNSpWEr/1jbd6x
UpVazHHnXDHYM9md+BEfyPvk+SorYRvElo2tbSXmTIITysq15DgA2WCuQoZX0CMO5AYqzi8maSpn
AK5hQzienePj04FmPoJSlubUI31B/V2cyByxuSXVNSEFbFxj9TMNV7gJlgBZNtDpwbEeYi3L5Lmm
1DyWeG5/2XU642Ui9HVy5cTID+YEYlT9IfFsRrbj1NIqwJpm/1SF5a6E9bIYq0jKBewr5m9R3Rep
YJZhDCc/AI1V9BaS69UV+8RTOXsIzh2eL8K5c98td009Zjm5KpwINa3wxdbFZtP59QTIu48uy0e/
Gx9O897q1Pb4Yh4DK3A4RiTuw+0zhS1YXWzuLhNIsiT5z8xvvI2ufNaywJyUZrckG+2Uap9AQj5W
tPr2vrnAgA4rV3CH88OlWPIDTRGVQyvylqDiwqtD0esQuJbZUZpHeFHCfnT7wcrDsgNdCuJafdII
IQb6FxClQnXfJOgs+vkYjOPQbB6E2ssXKXnu8+qpAruP/K45XP/nV29gWedFZWLriHJbuLkKDgOd
Hqpnkr/jwlEhR23bAnRGTM1k/AtEK97yICEsjUmGxRd7eGcMHcf5/IkM89b2lWQ5xCNCPRM4Jami
OvR2yGg042edC7maATBAAb29TGjtM9EqlvM2iUn8yKHK0BHy6FErDqSiXuclacS55wY/8ke1fFTJ
6mziPRPmZ0DX30kQ5Q4TyYdgqxNGGu+Yo2Y88Khx+Z095oDp6jMfuyR5BpV/9vRpuKDJX072xuSy
gC8DqxG9y4g+ukuKDDkawJU/gA6BOepK5yB0PbKfMQW7GlBqP5WSZ4r1pll7bA3o2vLnV2xe4ALp
sBwpjVEwf9/vNcHZlRWGAn6AJw0aZ4jIhkRhMS2nQ+T6zkBxU0U9g45GCHH6PYi5POfL6MCDMpzD
hafS4LZik66IKO0OKsrk+6b9Ty1fbYyi1H0aWfA9CZ/XrMXl8qMtJIPOfuwb9R5qIFDtvs5fsKSo
wpdYL2uIbK1MpaeptZEj40FNC6IjR1JeQQqmXP6iG8TIFPPFW9V5DATA+DaZ0cjkrlKCx2prx3nj
5ONJY0Lsx8S/Y9eDTetBkb0oScKToxJf2sZLi8f1eyg0X+tHaSejF2t+JzeVxAwZXhzkwbnsZ1Gi
pQpcNDuXn6OfXGpM6pSc1zan6vJhFHnoWP4OnYmCKfD2zJBJV21RoTydVAiVbnz/0xXkWfviY2G4
g1HDrTP8yzpn3pBRo3m0ajrx1RhlNioTjpKQsflDMBYyHKOmwjP5tuA6prOEZWCyaIeyo1+QSnvs
U2KriGRERssomSm5qt1CW40Uv1+zH2pQgNyYhRpYtSXv47Wbb0tUhl0/WGFiSL8Lc6P60Ga7Vxt4
sm4XihHWudCQA9rvzPsSJqf4ffvb+p29PtF+8jauFpQoMHQKgsoQh/x7KkwZuFexNIZpMhi7A6DP
x3Hht+J4qBD8hXpKOp/gjexWcUfCawwTzmLDFZ/TbACsGD/joNDXCJyXZwyoSwMX90/BmkloTFvD
NX9IKoU22NQtyoGDkGYW7mM66hWmH6+ZExWjgDQMHNKDxfE0UPBMt75GLU+cJNnbzS5uGMg6p3iB
PSbGBHHnOedJklaUmyUlo04JEmZTkNejav7HRgJiHvu+aTXOFSXO90rrbejMDsEys6nSmUxW4l5j
zw9Y5eKrVq2rw2I/kDpENDWCSySPNK+XMZ1xI70Y+X8vVI7GsCivS9axm+SGP6Teftn1a42HV1S7
NdOuLhXMp/f91RtrK+fh/RbHD1kGuPxGptQysbA1hgQuZKqg9S1eojzSAQ2CnEUKdZjK9MzkE655
bjh85VCoihulQSBHeMOoBZAJDh1RNDCGcdY7tfO2NtiQkbCkPV1D5jZIZNw7BpwaF7OYxj4s5Lqm
HRSLKlsH1vg5xizp+f6q2lOwIdxB7mgBOGJ0HE6Q1YF+cuGqHb1AgQbeMvvKwTH8Xoo18YJwH6pj
47L/9QO446CF7CpQs8vnJUVnOjOuWU/hFeqeIR+bvYelBFqxFHCckyMg1DoUK+a8MVc+NFrh+VVp
WdkILKdQXx65+dqk64+oKCoQhDKiqsAuDjE8bpCJXC1CU9RIZkLJqYlafpoZIlhzOZDp2k2MTp09
VYVgg6S0IkJgTcxOZjkKddopibbe68Ky+zQsOAuPh8K1uJjb55+7Flv42gunwyun63Ul4vJLuBSc
0PEaM7nvAe+C3Mt7Kco6e6dijICv+4RNywDR8dBehX8OIWgeWKvPy2pTo/UjVjr/aVb9IES3nPEG
44Q96qFqcgP2p1ThAFYBIv8Q8Skn2yKs/4dxcaSsXLk3zJoQABONtCA0WoFSWKcxiwBWbzCJ47p9
dhZTzxzu0mOcJJGZsS/HBEf/G9dFnqzjc7PoqCwiGzPEDlzJd+U7wUJPw2L+GP2KJR65Li3mCGm/
1uQNx0lNcwpsqtohp1mq0Geb7qH5eDk4Nvharb9cBa40vGzuaTOtkuWoty+n/0dEBJ2x+gi4HZMj
Ug7OiZyfbtQZMOv6LbqsswOsubAGWKnIpdQtUyZypUrw96r9E9be8VK/0i25RLB1EZq4iamj4sI0
xiWQa+LSlBWTKmwaTzjAgal/NzZQ+FsqEeI+o/H6fy+WwJCYD2ioUSLEsDgCW0sKxH02xdDYCrJz
+lYZBgkvhPj84X3iuojtCgnerMBqzFowPkiU4zD9pZ3bwBzbId460wHrjT2MMRpc1OlYPjsTGTr+
6pN2nTSqAt9YWcd/S26UvSe30OtFVNReZ1v9s8f8HSYdFKWXkerqzPQlufMWzDkdCuQ2+kPlZQpF
3Ef1XEYeROYLCRi4l1h+5mwFvsW0VQIGm/jVXs9E6bbbr6cXG1/W2WSmUBNT4iCMdQTnxPsqNI4P
2xybbELJL8bleoAt3Yu8YBt2xRFhVlHcYrl6Mb2h4dZZMmsXRH5ksHFwQejoauYJT72BnEBjTVOD
SNg0nvmVgzMmHrvaQvbBBv39oMj4CuEiDv9LxRBxsAF53MVBUbzOp2HmzIfh5sq5/IFWuDRDNvap
OLqQOyFaEy434gaEoat6Wa0zai5w5gKOJJLCu44XTnTY3V1TarYxp+nVhT7LtWNSLKEmW9nRdsGC
9R1SU+qns7EjAywHeOJDl+Gyxl90cC6FMKEkozcOSCXmH/9ifK0PfVQebxuNBzTAedLVBX3GtNgc
8OC7WeuepxAofNxslRZndcrkcxblR7ipjVGQRe5I+P1C36vnnYZrfU49vzLc7Jvb3qh1MebTdmT9
C0DVIXdKm2nUdm/APAE+2XBD/JS/3eDISsPhgmVCddS9g2XLK1vebUN3lcziN/vDHwrxDuwDdp7z
55+VzYlkcDdoO2cwCpw6CiA4iV9RD9bCLlpvPZjG0re4Px/4gNpVv58O+JMnj2BpG++8g9ohkY9n
ikygHmWJ65oZ5ezfHVnDytWB7U7gZuy5MP1ZtgO296lzE0ciFguuasvANZ6JQ9qfdxy4clpyc7Cg
g/MMZhji4OzRs/IhBs0PP0dxm/6WoMvm3EmBIX4i/hMVsbIJKQl6SFdL7E+cSKOIN7XuFQ88sXFB
6p5Df3SMyMc/cHslkqqDPxyxIe2xyZHSuwxaI+k2f8jrQgZKsdn9mG5Yc08EYkg1CyABJ3x6zc1n
NxnEMEs6Ma4Z7Mhdwq8lPLrpFucy8McSixV6ciNkJF6xM6lJJ9KTpoe3iGGQHH2Ipan58K5mLyYc
VtotqR1ugJ5EQ9xLscVqM7jf/cSkvij/yl5Npmf2ONNlYzlUN9FYQyyPmVwIaG5c4FR0B0WN0Odf
60C3j3ae5iMgLpmlouxWNS03j5JVqulpofGjWdPplbvQdqKlG+kakBk01SClEF7O/JT1Cx8OZRqW
uw/d9tPqNx43IW/dECEqCVdV766Gop4vXnof9ZeAA1i5K5qo/Dwu1AZtE9yRJOFG6kiRyuvWCD5J
Gg4zUbdRQF9/rx5JoXUnH1PsMkNz2MpXKi3rT1KEChR59tXzZK1M/o7OjRixqsUysTUWNs/qVm+X
szYJ0b0pHVUjZM6ifwCPLaAHAuVKw8bOlhAsBvOm36fds91RDi5ft4LDN2UastDnibCgb31mWdML
AFTGtgFv/PvPNr8DuZQWGwz5r6tyh/YrmrKjC3+QEDD0cqzs2jtMvlJ0D+r+LMJJ01+DhA/OsRSq
JZ/UYENO8UhlYNXbkHpS79ebmDF5dtiHEuLKkn19mSKcz5gjbBIBz5MUN2scMnMEgoFxHR8fl0Nd
i02H6fumRGVD6G6xRZajw5cthV5xSU/oREqn4rStyKLu/QSiq/r69OBWjnKUoOipOdVW1pjsXvDz
gGblYlbcz7LG7LQI7y20QQ+bQS/1GgRmTC3poZNlY28euyvm0E/8rQsRQedITzrZV8s5E/boNk8C
CkfzWqJMnU8FmVbPnLm8z5CD+kwrlIV31bx08YogNQFHCWwN4IyYjQ5ZMq0NUppFSZXgV+qp52TV
RMzWW9ZxuZlL19Ea+9NPvuu47d0pOTIUiZz6MLkXyjgTlchgRNI/8Ys1XeQRRRIjdgxxQlpyjaPN
nV3p7JCGctH0cnx/k7LxBQObAG1Kmky2BgYweJtxb4ipfhJn1cIOJGiUzh5bu6UUctJ9FxZxfYJY
BcAgnzMUk36Sr11duXblZnDdh06/j0hou3mFvl+49Hi+h5TSAthHjzPumFuplFxBnhus4+h5NcQ5
PQSPenOVWJpAu+w9wI5sJbc1kO970reAPZxF2Os4g3s2aWvr+BNX7wjmfmHNvVek/mLWKaVtI40W
bmzytM1q+AChoOd1ev0DvN6KDi6wAu2PegiGMjvoAl1QeMTPzZ84laKYhnEli0IU7pNdljfY4f7y
kSy4qE+0ZrzrXNk3TkQt50/Zldm0eVdY3Z29FklFcWWw3r2ez/ErPt/f7KpEHvKaOWU4+6Uhd1/8
h5X3ESEL4YEBkDmkXjbK1NOTFoLRiJUFt73BMCirZDcfbXURZilJmPFold75l9rf40dHYBysjJsL
+GU0NxstGUDjHGgfbkLKT5eCquV21F5H1b2cxkrthSXuJUcwAMk1BxLUXlx9kErZBICXjkd+WPn1
haxz7Pt6oMycO7jnRpeqvu8qGpw9i7Y3mkfLur1lBnGNON04xJODpC6UMp4fg3qq9spoCkonAUqP
XsOGVCw3hNmov46Llwxoz4a9EuG/AmAqOyFR3GLTwgm1ls4JrIKoqBrjRpQc0RwSQPqcNhpeXq3m
Ki86KvrUveWRII/1Iiilmge1AdChctbWwVhmq+g+WEf1t0Y3u7i6mLK4Ko3UEGrcQjcFpb14sEBH
n2qfP/wwbD+BwAoI8OkkBOtnP86/g+9qS4l0AbbbHMVn2yYn0dCs2JEYcS2dRpiOaJxIAJZ4FJIJ
qMlvUyKO6Qjj2FvspkPSt+DK4I7qIDz2PcapE6MoyoKOXPuCv/FAkm+HS8vm7s15A/iB1zP2LrpF
uVnxfkcp8hEFuPsrHylu0vjDppmETUr1FyPSRLGgfsdqmz4ICL2ohZYgNAr22fvgWBj4etNJyAC+
mjMRV/C/nZUcCA5hhh3VS14ABagbA8m6OyOqFiwA3FqVmVIIUr9cCLk6rOwyj5kTZBVZ+KgRhttz
hywdoRp3SCKH93j2rxBNXFW+bKtkpKz4MzvnN8Fn6JdVMzN2RppfoPkj6N8/NwtGVRya2myQznm3
LGj+USHhnmSAxJjOVp5n4c2AvNBeNNFXGxzRy9wxmJRtpgNi42K1tdUp2EG6O27biisZpLLVBc2b
IAmnnsY4NgTjqGSN4JN3iS4+kC6DfgdY9phCdy13b1yA64LbQLtUmTw/NhLR6uE42QgxVXC8zMir
MMp7O4CetEWDWPA7/AWHmrjQVG5fTzL+pYZicHHWABgcCt79pv5Q+XIpIiWSarY7bFi3KyT9z4m2
2rW1sPrBVdlmXglwGeZa4q8k1rqrQLcpBGXW0xncEMc61iYmTi8Hi66y9RjbPl4r+DXPd/5Qrbw1
VzKrIBAGX1iDhiplotFfIy3DkhC24RMTG1a24vWwOmglggD3dGfoa6E7k242cKDGH+el6UB+8JsW
7OalgP2kEGQeinOVXjXtnoyc4ZdMGw2Bl7/2Hu4IWk/MXKDVm38okCfu8vr+PfP5sMPoMWmCQmgt
EDbUxDBU4XzugiKsvAEuDVUvYONWr5IO23QWG6+yHnHeARN/PRAYltplh6hWF2YrXTEQ5mqpnUAQ
7BcaviQwA7WAdL/wgjYNWkgnspXGQ/b9GL1Pkz8Or4lIZgZ5jyLVudvynKlHp075tiT5VsJ2MrJJ
o2nNpEAWzkdfTlSAIfLudVJKp4O64b1kqqwrqUBgU8Sf3FbwX9RGUOBEHWesin5s6RxiQhjSlh3w
gcm3oRN2KUdDS3Mn43PNL3+h/GJIY6IWK+w8nMPRwKdYjZ6DxKaScUy1izrYqZMouAo5PQlLCnMc
/c2DmEPq0FiiJWYHbg54anLoyn279KDFiWdOMY+kS5FrLkkh5YxBkqw1VikIz2m+sdolavjip5AG
RFHl3AkptCzhkR2d4wTZwxQwZYz6sbeUxAzgG+qmZsbhOOc0N+GG8gk3a9svW82mJ1Wtf6pRCMsH
jwDKdPwlDsVUCsW+H937OFUMVERDmo8i/dPUp374/clI5QWyoyfN1qZ/7Af8FB32Ql8EmPjAJvJi
ig/L/iHNFVRp7RPcLqmUSG5YZg6M1QEjhgOeCjIeAAxtTXUupplRhhQCqm98miZ0VehEVjfD1cng
KOxRoaXB9u30ldXYrp8VmSW97KdDXmC+7GwwNlDcryo+m6nFGumHwmVNq+Z5aBF/Edc3cJW1YYh6
6p28c+nxlfB0DGnXC3L1Ree3LhmpcTzKNWVdHrz9QYrGTjiimeFKGGy4JHKWoYZ2FLCUV7pLdf+o
VKGwBjZmusjjxF56ISFmtopDzNzxLqK+PWdCU8HRvcPOsk6d3lKtnzQveodh/GapiqPoH7NI2pZ1
DaIQjUiYUM45jUKmI36IID87frGOkgG4KFzPwV3wyrhEuvoVj542V3IDJ97g2e/09kcEcRUJAggn
Y/hqT6Vyrc1yCoI9hJML9A2cGyUyivOC6niHEaFNll3hAjsCgdfoY8roj9X972XwKRYLGMBen8Vp
n/VP9X32mw7NBeyCAzEqZV/gS+GIYvr2PnBu2jO7AGK5pjTXi/I8ZLJANwuW/Woevuclbr2Tvnnv
uLuJqaTwRB2e6k97rXSwBedpqi+DvSiy8/Jakuhu0ogh3S1m343y5BkCzfUs1T+puu2nqfgjNDNP
oDpYzb5XmUodgVcesIBUTNZZ9EJMLnNvzr7HQoFyEN4h7fa5T/OquyVXql3vio4KXSvhEiQPIBT1
CsTx1J3VUtT8p0T6dqSrAi4qsmE0/iKU6okdh636QdHK0EJX2jQ+toQ9XXIPCGfFkgeJ1YGxUiGw
ZYDvdC/xM/0XUTUhcJFXnt5ZIuoCqr1IOasRVKCHBIKqDX3kV84wElV4RV3lgckpTQzOgpJxMSzE
EmOsCjOl738tYsd8X+SkMQNTvjQT3lfDY2FS/HeC6vVoUPSdCKZcLkR5x31PdWLN0KwJ8FJslLa1
qEI4OFLUIeU8yjNNvGliO0MY3Q0oPqOMzgpKWelAG8f1dR0H8NcVEJrYGG4/Rxk1GRKrW5bAjXZz
AtRxHWXSm3qJY1nIsRMkdpsQEc53txi2wsHLhvyDvQ/2WMuTOnkdo26QlSUVs10+S0hByEwFwfuo
sLNKxCBaqcH83rCee25Bw6AOCUh70CwbFNQ+rKjH35cTDlef3HjxTd087cp62mKH1bsmYFvTcdBy
JByu4Qi2b9IC0m18XncN7qV8QEQcdHO9NIz2d+xC90USXzZcAzG4NBYEYqV7aECc3bdZjY43ztTA
Rg1gtX6TPMdbIwaeGD/4vUfwHH8t7QspYpZze89ARpYK2tzrkcF9IKKF4CVHV/qU7oGdHs4slSdW
QScQ28ANbWFrf1zj+ivRLiDpzeGF5otPHPLHdhkFIwIw//Zo+/igi2qOp5OCux66v61ab4jpvVye
Rf/GHMjoATQDRH6dNDAUwom3ZJt1D2JFg2avQBlVHqNeZRhdp1GTmeUUMTa4Yg24YtyponoTxGY8
19nxfEgT2lAmQ94B/5jAo9rcLdlu9GX8+VoWy2HF6GzXDYopJONqfun+jnKW5zu2KitbMvbv7phm
ZlTKP8DXeHgYS7YTALc4e5D3zgzaYGREJGLHrwffc4ZmbY/RXu28TNgeESMfPIKbUBZnaeoqbGw4
9jRbw0SLA3UB1d8hJQpgNrwh+kkynmFV5x1+qwEhCswnflKsY3JqZyEoQ+ON1Np6esfZCsMHSBdt
qoZ8dniva2+YxAKb/3nbebBqTAWw+Pq2avftLXOSQktuaOP5mAnWIdFDXixInCsXjkz/9LGOVY/W
nUFSOs2a2bFglDZnRlMAgq2Tf4L70yojVuNTfivefFBtW8wmE+99kIqUFzN+zWayXPKN7qBu7qpm
ATCiLtdafzXLzPgHHnuowE5D8a3OFfLdRKdWrWsLu79/Nho4M8+3tKetDJlbD6OozeItfA498F7v
NLgVULoBXuc8XORsuTUbTtYDpylEyBnK7NAj8pXUBHdjQSziB1IsHhf0YILIdWpgH+fTM2qkHYD8
nti3R8cEpqf97xgugvMDaYs1zqUhbGkx7Q/YvJwvaL3brQu9hCB8Ww65Mqt7sVFoSqsLZSw52Ns3
niv7mGm8kOvufqqjgWobpVDtsYcgZvfjdYuo8uOADJ+Eup37GK5MCylHZh83RVQNmGenn95JBI87
LWVbSbVFeZLrZv9b1980hcpUoTXmHmtYQxsiimrdpRnR3viWPDIal+Wa5HCCxtlsgYQE0Kd6O3St
B2GCQoy4OE1tIUeJDyrkmRyZyHiDrZ1D4zsq/UCslpc4R4CUz0SbydXHbkH4iA0B5xthHvl9xzx+
a7zTdCCUjrAIMQ9SzjzoDYjcIZXdXQe9pIHyiFgmV8uOwgyViQ8BE4qQ8jBJQPDlPQ5gT6C3zn6+
pHwo8PqEAX0w6iFso4U0/JcWTmOJUuxH0eLTsN4+4fGbyZw2d2tlv/yKCO62lMI2yLlUGf1rNef1
I7fyIjkoc+oNbJDNrlZoejv1GKggHjJs09nxBtE7QxcxxzvJJ1GG8sC4xMca5fM9pXl7v1ZXY4JB
4loST9RUA5n0ibmQOmfX0Dwixow+BaMGOkDN19QaL2wr0Qd6GWoTKvXlVsHpJzjJHjh8vwHuZrlq
/dOe3IsP7+8mApv7p+hfF6/IXDDXVd2OfeCQUPiXNawv1D6qNMQdqYQotxbAgoVRKwrbF0WFhb11
E1GrEd5GZpVF3M0rze9xNVLOdVmdoptKaXHbYthlQ5RzsZCUDXue1YHJTh5Sz+FlaRqiVJ5tp5Yt
FdEgUqofOPPt5jzSmsT6+XEg0SN+FBp1w9l4tEuvOFlEY0G/f15pD40gvsQWjlUHKgvZcmiyRd6O
UYhEMbnIMuI9qCSyrkx6FEwt1yD8D46lxpYIxqcPSVRs5i4nq6Xztbw5a1XRo9mvufNaqkwpp3nM
qQ6iZEX8OeV9PXgtPd/66tbI38oXYbwipOWpXkBGdDag+IQH8v3M0bgLfCCMbWiS/Tw9ISkajhBq
lBZ4BYbpqhxMtJhAGP4JQ77iGKxKNc6olihG82SX/p36A0UM+RIxVwbSVae4ZihNadmEkH/mm9u/
rPOY5cV8useveObmkAAY2tgzEEwhEHFXa9Vai5SUJrQY4NQcqwZLOJwj5UP9wfTyH+0WhiEJLDv+
j9gamRGZ5dIvH4fHXNHmd1kAqaqMHttfm92XI+vQeT5jHBaTuwmT9mWzaurAxYvUD/AXac0l04iC
3aRuKV2FSswbhbgSgu+po7AeZaYoH/domjZQCv1oDFMzeqvPGjEkKL0KE2rrOrGd8SHQc5GKQ2xv
1mWG9rPvGxzH/+sdaZ1KQBDo3PoQNNIbuhCyJn1fek7WDjs4t4X0JW9x9hDarAiqInQDLa1FebBe
niVoRHFsHbclyNsDXHN+nI93gJ2hOj1Ru9eh8PBSq9sAdi8MB8/f7qxuJHc0PDDDDm57psgQdMis
1XDrFRZ/HqY243zHX7MfO68TaoZhZbpeDtVuw0XaTpNc33YIbuzCK2maWyumK8aqic7EHCQmjuCj
nkc1idPuJybQlwsWfetfa5ckPq399iNKihNV8dkBtZ570zpODCEwTFChoLIdF6ZKGINyc0oKOhsD
Axxz+tOeIqQ6S8IwMc9bM7PWU7iOXFahkZs64/gQEuPWQEwXzr9IdpgpsgzlzntbqdLWl/VZHEpl
iIGHwXxVET3eItvqXYX4ydXqxGHFxvQT23sxG63U9Eq7YVXFCoNuxB6l3YcpPmXkulnJsuDHJoa/
lskwFitQNK1oY+YsZFG2ZtmkdWAwpBOn2Hr5MMA4ZlBVhRia7xjVr0QUBjhkuiFM6QG1bXdO+7Zb
3IakwjaWXXDBeMWeXKaTbt+yGYKabt81udwh8MW8zt5rjFAAyv/c3/lompgbzq20aS0GR+5D6cO+
Apw0Je/qMeu4Fgc7CIzHnMu7YJ3gnijl0u1cvlbJOZ8C/HLrxff19EAbgjNAAeIFJB07p0cFFd6q
Od0iD2Q1NjyAhMLFxYc6xTcXS5EXp/DRCZEqEu9TrZFCPGrvBTx517ebPCr+NAr7LLy1b0t1lcq5
BvO+ou6zh1MrxMAHWpgQcaUDsWuKh5idS+9SvIQzQ17K6VR4UwdKp2mWVLBsG0Hd57B2aDv+RGdt
c+llla4yyAO8oGs5FuHDxguKBaOg34AbPRYLZ87BpkLK17EibKcMGMFWPm5kCVs9473NMoTGZ3KH
DX6OlbrHh9ccPyuryPgiIEBR4DfZlsABYNp3lo90BNb/yl0Q2xKhgMv8AQh7FJmIXqWy3ITAMCgC
TsIaUPJyb0ZeMPS0duGz//553ai7+Adk/r40za+xlgMckibTk47sFKNI+po+JXRo0IzO9AKeUNWI
i3WoNblVehSpFvGqn836jvQnesrHI4h2+SpzC7yKzN56k+3cAf7Tm1rr7mbbmeiXFUt6ldGo2NeO
mhNYJv5f5BRvNz/m+/UH25py/scWPriRVkU3Mbk6vgqVreDKb4ymPPbZ55MFwR4kPrOMtANWV24d
bnWVpgUcHL3lKs0z9AzATUNnf8nda2GQZOE1l24SfB8WR/sQ5YpRCseLuGgCEedX2Rm+LxWDut1k
eL3sg0oh7nHq435uBS2f0Omt6b1bqrpNqacW7GpsItTYhBeaBsUnjOFXpkrHxn3iw/DOwXn76MAS
IjXGTIv/WgE+GrRQttZ30lac6J50DQhXIi1mzyLC0A3f+ENGrmhlVl46+W2fvm/09GpDeHhvOUjo
UkPBoU7LuST4bPSQrSW7Wg++71srLWRdGNhuAynvHLOSv1EZ4ZX/jx935LL8RTj2V5SFtneVElKi
H6W4nrpHZZ7txJKI1uJNQhqr4GsQwi0uUV2K7eR4w249A2c36PaROTZkmityAkbUG/pyEp4+xupS
VtYhibDYx4cqrIX6rQf1/0X5fDKadCABvcBdrtr45N5PmrLY2B7ElNCW2Dj0kfckUbfjY7WlYSW9
APO/SzUgFthyx1Jsh/MWp+Dt7ME+7UzPPv46c0OeYbOuQbFhqtx5PhsivKJUhmNai3Z1u1nYWBTO
c6nQ5mlu5PyXYsL8TILGJotP850HotewDT47dIhWgI3NeCBKyKF2iynM6jfOTy7SxoHLKXrIxQB9
auweJodJNcv/peARhnl/Oo4+g0JPbrAAes0ZbKRWpNR450nJv/OvZ9E0lkTYAEffe/Ytmd2NiGm0
Z5OAVJI7p98WxrS7Z+OHsEkPpmZpN3ExoUQUpLkK38GQASeGeRM1vQJGBVCBPsz857tOibeocuBd
hdJXP4pgbrRM24xqstm4jkXLdPfm/Z6gbLKuPnpWXusvpeUxZK/Li5rzn8zIfpmNcpYV1Y8CfFU+
G7WBD0+LnWGLZbXhWHX6lW8m6rw+Hlzp1sxxMmPK0giAZzHJu79/0tTgHpsKUSgIC02oGLwn3K9i
Pqhqhh9ocSa8fPjCTXIAQ7ssaKT8xFKbVCHvboU28jfNSEgLp89eL+6TIa9n00PLza9NQcVg0u0J
ezFAIiD2HuP/d9IMTryzgai/NLize9Ytow9uWKIuocdG5YDFMqlKslQ4sBLHdfpMyFT5Vm18Wyq7
AAu5BqBburX3IleHUH0UDF1q+pfSLLUDJWPRwUSO9eujUuso/ZBwZLbSadz0t0+h5Bd/lg1gymVT
Lj2EMgjCaTCSSh1wOO+3zDEUhVxTmLhCaB/V94CAi2+ITzHnNKBSBUsfgGFSEXkLaVXlfDHXQzbV
wGiMzODHLoJmT3YOM9XJw90z/u1E9DUEXzBrrjwgxT+7EPgKIlBrOIRzjTlTxeSQnwHIW+xctJ4w
0dMrBzwk5/Dwofx5nT7T22QzopODwXerK9H8NgOIi76+D3FBJXv4onwtqVwbwNZV86dvIYDTvekW
CVqFBUXRsjom47O62IVsb5NNW9ng6t8qxYfFSAYZaY5WWyRe5NohZjR47YgbMlW/i04nXlpQ7anC
Rjokv/uAiKICgHq1IiMCPbP8vMcnZ6Ilf0ZW+SEYQmW79X64Qg/CLYZdsOGtmfDdRvWoN+PbK11p
PC2vE9vkwN29mEEc9A+g7VSEObVnRxsCEt7R+YtBmObAdbmFC+bUAj6lYafDmZ4DcGwbc3bZRa9K
Syz4nr66UQIrkyrqE0fh9ZwsPlHu3ZPcjTPxIJheRDWahYCMOOmECOjnlHXSsid+cDMfwA86xyXs
ZeOPdFmFL5aomXdXQ6IAI5V+h0/5tAglnwKuPZEiCpK0s4OJ4NXAXIr7P6PX2TUN3LFn92R6akYN
kfiSUb8+vT9O2+pPntiI3F6hpJc+JAN1YQT8n55GIreffafdPuS0VXxgSwYTWIh0etL6mzNLkWkb
AYcyGNBpRYgJfAa6qA/3swizXD17H0NHVFualEYLkdDWhM+49sULqibbfluoHEjtUe46e+1m2TdR
0QzDazoMuSXNQ5UCdq9ph4vasFgEVjPbPYLr1fxPCs2lWcvXHjoejJdgQWK2kc8vC8kd8ALYQowO
2JX4Vpjwv++dyWVCHnbn8o++FwjsBiLO9tg1cbanCcLcU2gqOAkMglOteBTPHbs1MyOjXMUB121d
XrnBgefRdWCbGYXamth9iUiVlZLPaG4C+JjGVrTXujUeUs0h/2fqdnhA0dlRVu+/5BDEUT23RzM2
1vByNpXB4ZLl+/5D3QyFdfyuwrRpzkChNYH7VDZbWzQ7DnmFkNfSaE60bSWLBNyu28sijCxdliux
+3q/rgfEE+MqkjVwhPZP/PGRkDTfJpqfUkLRSdq9Fp2RmCTJGORsPOxhFOBTQxAZVvMkBs2ap3b9
c7rqEhY8mYrIt4ZPCoAtlcr5ISdABdnYwZBo34RGT8Z6ZBCRMqMEr36gpza5S6qV8tCu96wrDQVS
93gIO5WY989fbjvK2jGGPxxBn7LVET5P1zeL/vH3S/Oy9hrhpGRIlZx9R8EZuJSbsW4QH/FT2Rks
gpbcMyROWV5KW5UfyOU7OCQY0ExNXQ0oswYnI2/hs1taMNM+fLF9UIZV2H+IrXwDv7RwMuYvG11w
n1m/Bf6IaFdezaV/3D456dBVOJitUsLbgbDhN2M0yNEg2SRrl3eQ2Q8r5rx2OXWCuHt1Bn6CiJtW
ESsFGNGmCi808JJmaMv9VP7sqWblGKdBKvv9qKbpsGukQCgz1f+DY7IMsbhGLh5Ypn6QJ04v7XB2
zT2R5KfmeFlWKljqfG/JUxoeAy45vbgPeSiU0awo3x4WeSxp6Llwu1h9Owk2IhipTxTsb/SrvQuB
lq3Viq3K76u6ACLdNuj5Uik80empSReH7Loiuyw1DBuJWkHDFjDFSZJuepFdnRqqz3NuFCRHByZy
i58B4An+AF7BQgCqHuDjyVUJzBV9hFC6O5gP96I0tds+FsAdDCUDepkV0U0q5ToLFiR3qqt/lsil
ONgI7UN67vrB6lCHBFPPWAHODjEf9apGXm+dG45sm7HKxDvKGfxf0QBmWmAQrd7bFKfO5LLFCJsD
2IGY8JsuEY/V2GVPumPiI+rSbLhaus3ziSEZ7SVhrto8ZvTGR0QQid1ED6ILW3KuaDOXpe5CsB29
OIc+i9BHcRqyEcheZlF+3pmD1GjjQgunvElzVP+DviAZcA33U3m8EJn2tVUHf9+B1t0j2AF/cUWp
2G01UIFqyCuIFCIqP4DC+qYou+YYdUDporIUY3WgeY/B46D8kmpd4LP94lEy0Xp2Bkxwqro4TamL
pdrEEPF4oC222EBkgyemxEFamMZo8QgdTlzRiuXTsArrLP0gAPjYqwVvffE4brmr8D8iEE18+8Mh
4/bVx9dwjHIFEvbIi2PDNb8D9ValYRcsj5uQQCfqga7gzIGp9aLbijfMfAfmbX7EoFVfAXDfYyFa
Dd7yKSgh/L852krP5Ty3WUM7Rkbr2eEwrin/4Ek1tfN5UV6BRhsD0xgIDJ+MV+tqjWpiNISKzA3q
Hm8CvKHAhxijEQNZzVx8pd8CyfRsMuGhxq3LcoZJAn6llgkGBbxGUe7qxbPoTMDfJqfY2OUs29Q4
wy7Xx08W8z6gPYKtGEi1ZeWzo1ejXOUNdjLWi4wT56qocIROQOkeyxksMD/+Wg+oJCL6TXwUcwM9
Ge+MNMYuE1CXRwr4pqUim0FhFKZqH8Qv5hH49Iu5NWh227vkfvhVDj0sHFF1Yhz3xV2yKb4ELe7G
Om7HwFIAIDLWgHdlyXp2VXOtY9Je2qeqnq29Ep7s+PVQCY9ia9iRU0jVibpfZGhGTEcJHipDNR9u
bqEDvlIwUutcnfh2hNwL/Jgzg3u121fJDsgcrlMsfJ40h5YZw58Ojm/dxGdWKdXLU0M4U23M3k0p
V5KmfY2jB/T/Hac+Ompe+1OWyDzQX/SnCwS6WZekVYjBtE3EpbYiEFxQ9nOhNaKgKiDtra0aUeDy
oh9oe7T/PQ2DXkyqqHAmlHXNFH+wXPJn3o8LkHbDXmJa5IXR1ExG6S+wzSqoqI2Qkae/RNYkbEQq
mlDedjWRowRozm8EjmXzPDeKkhTM2JwmOT2XuEBg/XdKvOUvNHsNtXgY7f0RbnBWxPPDIhIKzS8i
hP6FXijFZOGAs9uwYKCauesg7MoBxcHdL+mHhPqbSYb7Ek0kcDY+MkQkxppfa15nMCIApUiRvpg2
M8SnXZc18htwhl88NLnGRsHF4lBgB33tNIiC8JfZzFfRrceQarp+7Z74pHOB+NbWAAhXKJhWe4Le
K/swsKtC8sz2Yl4Zl42i6YYdD5OASDOgXye8ePsb5eq41/KuTpQt3PM6+W/15gzw3/QxwUyHNlQP
71vj/PkOEMElSB37KgmmwUNVqD9Mttxkrqd6g/q/BT2SsAmusL423vwOlP20rBkfJdn/YTqeaViu
VswKVofDuEU4UBxKhyUZJT/u6HaYnq+Szcf1FrYG9CeBXa/Coel6GrEBnksJtg9w1L11lzrKiAmW
EhcbZ+sm8/R45i/cBslUN5FroQJIEZUAgQGZ6o0qOrtgYra3vQkiFIr3XAXvEMdBd8Jg/mh1BKCB
34nq3T+06jSAx0bo37GLuV+DNYjfRfkGUstBegrVSdrYGesoB+ud94/sdjLxpDbxm+ktfj369lt+
UEDkV3X6RFJz1lpZoGjduywH2b650Y25ujqxiMm68KFmc30/FnoVtwkDZK4minWgxTyoCz80/Cz+
NadTasHnuC/g2YbhDHf5bwCyHbzbTr6Az02zv8eVcjmxkb6LOny1UXBVjHUSza66ZwEYTOy4aHAL
ikftDnuodzjYuEbCWeHC6qri7UOlqKfo893rd7QvjXnBduz6fe+s8tmLWHm2XLE/w+1JDF5o2t97
EmDEG4QulWdQVIUToPZaejlb0pMhQpawEQqZqnbakJO9jZvROJKorX2BTKER8rggc/nZJy/MOnRC
kafyuvB6o66nVU4E3G+bgdOZ9Fr2Qs3SHFN6QOwTKPBoEp3IwDAUlut4GgzR7ebJCiRWzj2qd0sY
TlbAdQYwMK+eBU7mPusmLdwMQgMfXhngA3ikwh/1xM+0nbiXl1OSkUygWeGGm581sfXb4XK1941L
JID+k9zJr2qf+fel5s/abuccaRDQP3Mej8K08LyVzmpSH2UUERVzru67RtedxHimc5ABXleVdBqh
/fTcnPtim1diWH45hCz0qcZOXI+M/vppDEcxMii67a682ay8FBCp0q8B+iM0bUiXwg1wiW2nawA0
aEm2lXpoq1DOET7/aZKtDhpGTuiiso/nDGqD7mC1z0s7ZmcpZOD0VObLXzOfnIaBuvZIqVqyJjzM
nvpDw2LR4AD7ozLm3wmou850B7oODf/nCw80DAVGw6WtGFhNwUJtWZvTGkK37o62igNQBGtoLtz6
TYgfuxQ9wTJJcXqHZQ7P9nHErh3aFO/c4djqaeDFXGJhK0LQNVXWuleCYyMluhIenoYTJH5jILs0
RUgy+VGbcvYXAMjvCpvL7NW7wTJGKT4oTFRS0pZMZcN8MENJLq/4Ifmp1A0oloQ6CQnWgjTfCMtv
jWscqUIJNvTbPmuHWaScCvChL6s9E+KYTcEISmBeMaid4iKsD70ZqMHpE37LhzfSuMR7DIra4J5q
WC0o0w+s7wiLdqnxOhbZYCNX6/oHv0Ax3CmrO8YvEsmwt245vYStjSZPLPMciXJr+LIMRCajzBes
8T31KimbZUSOYbCATU4QTIj0L03Wx/n7goyXX2FmLf4Bsp6xuFGOV0uz1fTxP+uBAojzbm3rHy/n
5jsJ+wFrTMVaQ94xbMdge3+dmFIqXugL0jydMqROh0YWfLarh3OslJqpx8Z1DlmutyWZZhEs63Hy
php281OkLc8+wjujAYY9sonnj8Jn6PKnZ2BSYWhacAi6UPsC4JOp5RiKSZto+W6y2eEkvcQ3a7Fb
OV3nN8hBqCzpKjYbRln5+h5bcy1eG4wVN/ECc5swgEx3O0QF0/MnfPyTsSVUb9oAOVXZUWyPrjsE
22vc8T92PVlF3NxWLV25d5sDVxDB+s1O6e0Br5vLpDMhWNrtqZ5/FbR/Xcd+EpJlh04/cnC4O243
yOWelFPalmXnoJC2ZsmnI6e+TRWYso1cUzO6QhlH1o/kndOIuUX3cPnCpDOmMyzjf7WbcEiXpf4d
j4v6HvKnIRdplYMtpwhWyICN8RM9CnX60PYdEdsWGAT1kxduQxRhJG+jvDvhVaqGvlvsvgn59mcx
aYepZybyjah3PbWgHaWt+EYjBitZb7FSQVa+Sm6SkaMypQsQB1Za3g6JSRL3dh1XCz8j/pSaLXBA
1B63mLhhNmlAzZntVfy/rPGm8q/G2a/2NaEwrI0+zivpvzEDhfV1VsKdxe7LbguhE7Cxah45d5+U
0NnbMcgHOIfwE6cwRrg2qTNhyielcEZHr2E1rYESQVrxsf07SJfvhcpMSB2dQZr8a7V7llL9lwL9
JrIWWyRz5Uq748KcuWw5Wyt00qudXuUJZG7FdtHozqGPOpad5cu7RGptJSGqTRa0FPZ992M+WA4w
yHNDNN9QagOwgHDPeKH+RLf5dx+ONdJXixt0m/SO/EA7z9TrB3M401ra6O2XT2+4t81b/YB6z0+K
U84gEKEuuXashhINQYAFWr7FTV1faorBbrIL5+u2fas/KryAsankpIxbFE3iK8MpR7p43pz91CKn
3AWHVtxQ3XYieX42i6RpU5y5VAOT9ll+7v8GVa3+DO5trCGvluS0M5kBapvTleY7ZEAs9bRy9wbe
/u/PrfC1K3aBHtnv9O9ltEjDAf1gw+XsG44YnEqVWcdSyE7pe0OQyfnbgNap8dN1dmHg/nzNtax8
1kCRlMjJhPlngQkHk9956MfmmOXbvVZ4Vs0XiiJgG0i8VzPUjYFRAQwYudFOWcg8/NW1iv8sSFxt
8NPjFgL67thdT4Wkn5W2Z8zx8zLujiIDuWQvFnKt9yaDIdyxktnr/FcxGAjOc4BaWAkmM6CoWe3Z
NNLUCzRlzjHdroaW4X6uzVmQVNe1Ovl8N69lqoxNdlUWAevtIPdgbNcKbGtkLPkeL1tnKslmLRMf
41pl+e2H3JQCpzOQS+0S8KjRG084iF/gFJ0t3TEOb/QUStrYc1V3H0RhbahbbTCcNnd8tiyOcuP+
+rA/XqrqKuhSGklOpTiEEajWnuzyYvGu+3u2iJ5+jYG4DpLeCC9JKBvtFzM3D2bQcq1BEoOyIJm3
GmiE7kBkeynBJ83bc3Z0KjLre5AKBtkyobC5kkpblPOp19pSF+izmSVKlk+eC3ndQE+/GWp4b+Ye
2Ht8J+KeSKDDE6zHUBOxzNeRkzqYtL35CxrDmOOIbONTGxN7oN039oTPLkme0T+Y1tLwGtmapqWF
9YkuOBcm7aVQLj0eS23n03A6EhEhb/6if2G74Esm3kldmTFqcdrPHOqfwfjNqdtVW1mBXMLkFjS4
4pgd1r1C3gh6pJHfFTF0owDFOmNwnUJtUVYHXTCCy8N4u55ViAhlewQN43JfB9NMlv8sSXXZuHPJ
UwaXOYJbGCm9NLfe1GgI2KPkki/wnu2Ipcmbylfiv9EYbwRo/rfm4f/O9YSzNwcEhgvlpUJmWwDq
WSsPrrwSD2PZdqaEKHEiBhSfQN+08899f/7HrcryzNXZvRhtXrBMQVspY5iuqJ17WH7+gt2dgJKJ
Q8emNbizYfcj6eMvpJ6g2mgMnw6okOODtsU++K7xqS/elvmhLd+C6iQELrQN03rctWQYtN2N53ys
oRwkuLw2G9OftJRdezmUN4DzSdvl1ABQ++uC3c2JSHrweorFimZZ8yjnpMLWUNtuRK6o5E/TTpJ+
B+t1byg8ch25YFlcYGaSf/FBSz+3v30oxa1R/4IgvP8s2YZtX7B7XO0txK25uOS12MxnUcIjY+zU
1G7wX91KM7WLvIT0U/3pn/6BCndYqP1HAm6PWCIh0lwSEf8HC0QazK2iE3IhIi+cokqDo7MZMQWk
X/BG8aUNhtmcaQPAGJTtffT/mefb3rGgsR1BVjw0Pvf3/WzStkYAVWvFSicMabNyFnQFuZ+mZpgN
xcARF6tEKLKYk4ZdkMAUc7z9GYpRxwCfRcfbMwhpNyTHTKAAOCF3enb/JqWjM2q7TkRGW6zic63p
F3mN6LyUZKvotrz8XR3j1SLAJ4msk284u8WG/GF2lUIS3RhP/+xrel2WOrSn9FA8osLkldfEY+zS
nLIyThQA+Nort8FkvOZHR/R/MbM00/XLtiRn72g4PK1HyI7N4l2x4h4Tq4WOoFnMadeAjPT9YSCM
qQJor11/fVQ+T8XVDmI48m/DXc726gVAFpMgjOnRGkBiUo0nJJUkHB2KIQJQMKrdDV4H+QbNwsFR
8BUPOwkTDONCcJjjDrn+eFQyc3jqSkFH8F1H90WJltF/qHfCZfcaqaH6UNiDL8qRzh0tWrLuBaaC
WpYxX8lEJztzp7uFR1VBjtFYolSvA9sySzQDDrv8aVo3l1UGl3qcxcXvri6DMpG5Z8E6WkJ3Vqpe
QpCuuXoh56AiGA5tCGeP5sb+pEg2g4uERKIF1Y+yJ/3L26U1cJ8YU3Z9jz33OjLjJIE/UN2LLa8Y
ldZ2dU+hCO5QqNtAlYoI5Xg6wSLKwq/CpbZRn84c7lGwTLksCg7UzK+5CJcTgaIv/vgOvrE+Wid2
alk701plmyGuUEnU64ZOcAjBk12TZ0qstjkRM4jNnw1HGqtoJXBOZkmwXJR4SJbADjSC4SfJlObz
OXcJdXaoH5N3V2lt2tRVHOVlE9oQ8yR+it33FG4rLN3o4o+2BeJobXgzgxuux0Q3WNdgvDl7clOQ
WgCoN3rGTH673+lTeqgnmXgBDQnWyjITigTuIu68evvHGDCJmcZdaEpqEqLCrD3ABLzsEYofCrbX
E5q9TOudbW9XRcZERhudEleDVdrH68AKAX2NjVTRWDVb7wqoDZNJvNtaA5FdI9sxiJ9SlpfgoIVF
1cbY/qfOrnTfO9pwBLtUNRO681XG2gtvPx1ZJz0j8GOhtgatenKgbe8fnVt0Ul+fdk6xB6OMjUJg
G/VrsjfoBPZW5n/7qXn9PH925L2AoExcOgeajddg5ClILc2FE+v41Rc6NFbm8ipe8KJ+Lgxig3I9
6C4xwdC52dvRoQO5rqtApTysTA/QZiwBuIS/GyipqYUNmqusvu/POeuJbVUIypuEIcDHGdpTvMRg
vKBs4bI+27QVqzA8jOedZYVCDwjmrF7sAmzkxLX77PUjiXw2dY10gd4G+K1GYpAhEixhsGbi1N3H
UrNQO4rOiydGhZ9XsnJBPbA2uAHglVcduieQir9rB4JNP0XKDp9uoeEYDyBbG4/OnafNVyGx5S//
1U8ZBvb3pSvG/bLGmZ5LMJRoZO4Uq5QmfVV3cpfpDWTCSwXgf81JrkAXQUaY+xQMCpJTVmAD7yuk
AduAG61+9rvQOik20MbsiBheg0uJ6eAcxaMzBLnYkctGGfaGO3BBXs7cAWgfujoEXrMXO5bG8wpO
s/XA4Ac+wF6yFdF5Ku1kW0qoixRCA9S/7TaTbyr7cjpPH6AbYitGb49dUfLIXN37hhLMJEBpXtdL
WKUdCYL1azNO781cX8rAp9TvDn2rEENAOldHrb7R9Yng+CPXJqoaT1rk5ls3m5qU5dPBntknsGvS
hq0SsnDlV1RXJb2IlV5iX2NCf+MFnHhGK7f1j4CfyGJWWYW4hy3Hi53MFlXUa06Izy1h3cSFs57s
k3JSVcXIyxdOOsPSZlFWrsfMNYfUzhSXw+MUavGQb7JAvwvWWiIJ5HZKUBsSyDdghqG3Pk84goWC
faWhPjrSTG/lfEXnMsyPhI8tnnif9YOqWpcvVWl+dtNvwNIPjw5vwNizCv+i6YnLZTTuvn29TGKk
KSAhg3qinD/WORlwt1BHNvqA85Yj6gJxaDbKYlrlGY8C4f6ordFTBWZvhJgJyBT6gBvkx2UTzmlN
8tnEPuCWG7Vb+4EBG7dZ8JAU0cksvP6bRMo68NErpzOAyUnFimtdiX7gqlnBXejxvfqKpIizr+mR
ndFtNCApCQAYVh2UngGJujpbT8pUC7/Kvqw96MblOUwFaOmxZTFDCqI1OIIvb3QQEp4+NwqyOdU2
gE7rgmr3Odb6lNmZk4oMmkGpWKR0qM8Jx4eS/3TqIiGj6RifvyOGKY3X7l2WJib4gjqUBZBtodv5
tHM6K8WHBF+q2I+w6C1dPzpAmJmIm9uAD3KeBV6jQTMHN9l6K7K4irP4DYuyoZA2dk7Ja7cSNSTI
9ZMI1E742wuLPJdVJvC9lZFIrpxk7S3Nhaz4d9WeHBl0ReYsCAu+Hj2sNU8/PecPZzbu6XbEqjPP
5jYJ4naa7mfySCHP+0uIxqTBZIDDLdiK2b5DwMD6Jcy0H29BR78o41sB/cuEGcMoSK61Ua3mx5jz
StC51qDnOHm+Km9NroJZFIo5KJ36GtDbeADV6sVocerRdK1ejWc+DyVrPHhcHTqOnP3QYmnQ7/Bd
iPMXM//WupK3UD7oDkHxuti2dQgc+zjh1FJLchVICEd3pRkvXbRQ2Xzzzhpw0hxOEnFf/8jI15AI
fg4NqoP2dwYx3WLT9Ffd+f0X8qSaeHG88+CCCB+fT6D2/pJVKYTGk7OkSNbuYl9zAvFwULBosdQI
pQDuEDniDG6nWoyi74fOmgD1jRweGGPYM6eKWghL0+pRJN7CUa4j+q5+JovINAWTj7uX8GF3Slmk
QFhXDLMvXy4n4yb6lsWmFrwgZhLCysgUymaReIY7LL/jKlqT56M/XVWw7ygLRtT2sz47O9P7VtN6
YTKSDGv5gFAEH1nrnANq22xL214R62/nSb94zLF8dKhiWcpEnUfGxCI1u5Q1h35DAT3xWHMoKE4p
ptd6LvInbKq7LDMq9fjMYAFOVyynDih6CyEwzyV/OuW1IyTIHTM0I3E2gX0SYF8M/OQAq88aepEo
5nEtyjHr98HIpfx2IMFejdi586jrYvQpwhcsNUBL+zenpElsZnn/wJTV51zZBtnMd5qX9+Xa+eVy
0/wMComwQoFiObCw3KgkVVtMfciFLLp8E4g6RKmKccVt/64+k/fswJ8F6A8UbBUapGC6avDaZEUX
33jL3yKzOOwU5uNmE0OHP0j2iqBwd5/yYHh5wjbsgXWREMoGsyOaoXkO0wWUVuBdtRIFURpnN12W
BGQB0BMgKGjjagGyp0rdezkExIw17k41zodrRcuvRczf5W3YS4oJWdDoiREqbTiqOWX3CWYQmJAO
Wh31WHooOwy/eo+NuUvevIXtqBoCpka0pUjQ9OI0hGV8LK0Tje3iI3zYbfvmob5mCEyZn73BVZbK
S1Le1itbdhvFaTAZImMFyBh3yinFbIW9DfbzOPwzCL8598lw5Alic0yv+8nlwq1D31ruiXZDCA37
ri1LAfi3dcbfjGsUJaN8b8zMLyoq7m8UF+WTRJKE6KCoeXa0uO1kGoF3ExjPRX5u0GG0iDCC0TQB
dVYYDoYTb7NZaXHuGFq4QY81MRT5/j6K0UN2573+P8EEeSyia/TNo+qrR4cijfIr9KtmdkZ2KkyN
NJHSbflXgaMwTWmCBDM967AbkaLuaoYzpIUzF4ZqmMEOhhfHHXbn4zOtJQLYxUnTUEl3OCwp4iUt
qXb7tFO2VtIhz7tIkJdHteSirxCKS3Bwcxhf93vLsEV5ix2ydxRwHM8ls8DBs4nVvWt0EBnshKwL
gvI89J5kjQKW2psmot8j2aSdlamEANf+Pg2uiZ4gU1FaGuVhqubNnEPGTJSwKjfItTLBIQjHTpoK
F3yJggerVIPnsWhovKAx016kcBnxKte5NmdGP7NpGJGRjM4Z4MQGziUgdFgUPN7MbbNtQgBg3q/l
XIYlJE5ZgMzcOkABhWP5HHVApDEGYlSmtjE4yi6mzgyM+NzWJ1yXJd5vFibsesT9efEqcYJRtyyU
G+fNkeJad5Urnem7iq234JF1YmcQMy8he7DGCLwZok7W2bV+i7uysKGwJa/TCdIl394i4wteP7HQ
Rk/rXgclhMJC4m+QY/L+FVyf0N4FNG0YIVkYpq/weul6wOaB7nEChZU8X0c77mrAnLLdzzA/lWWZ
8SPJU+wZZVfM3/3f1zPoG+grhB5kmQW/19IheG3kcErny/SNR47/ggcbhdOnTNrsZZlegPlmJ/WS
fBQtqIrs5d8KWpeZPqyFiW1O2axaT7xD+Gveo9QOxznzaexS3nNX/6mzGeXZAXHnIL5r3mwQs1KS
SpGxYguzp2v3HotJsoEEpe4bCw8ddzQxTLT6x9nrUfzhboICiGrzSydKyaI/wp67vfkaHrNL07La
qZoywW1OVKM8G/Cji6KrypRMuZL9nc7rdTjusEfWoAgp1A9Rr1z3bgrl1zg5Wnc42DoFs4hF5f83
deIGgkY/jhqoC+khCsUoEQYhvaDZ9sWxvBpmUuWhSXUo00keWnknvj6yL+BwTZG9oqlOhkdzKWnD
3EETnsw5L7kXcolbpbrqbX3mhGTkNoJB59eOoIwM3WvQSnAO22s4Es6toBmOWcYY8uJnnmdAq2iR
m8NZYyIl5yTi03FU/Co1QfXZ3zy0ERFU1KwUYmxNDDBIoHjRIQ3J2613lvStLvK1fo3sNwEaTWBC
DqzMeg+tYt1C5Inh/SgeS4El+KIHivZ8i0bzRO4jRZDWH8SzANPZIr2jn1imGzrTeIpTx9uj/YFp
+KEqft2ACcIJZj4im5mZn4ImzSt9Q6gY2TXz+bBh0U5phNlREVAtm6fJCWxcu6nINkOJQS0jkr5s
mpp3VVH1X21J2XHTFz5ipfkJw5bGuiu2Im04cJ/Q/x/Nx5jvtNwS8Q7cJBG+1XXG0cJA7ckVTMUT
m9/2E8qnxUzdA8idZO5+BlojCwkan6rHEzcqUtvAYsd0g8lk+V8nHp/xaqa4JyEUKMOnU3uo7M4a
0BJNcdi3Z1sNlIFTUoYr8Kc3hvhX/33ZQ5KKWXzw6TgaXrk9Vn/F4Mb2Vx9Al4QLaegdw/rg7K3t
6JydMea5k/anAXeujt8MGxvOHxmmis2o1ZC3ZZcINxlwC5yZEcrJPkCfdz4PwRaN1DLNe6Jsy7yF
RskF9ltASj1ratmRtpqu6QqzTDstxjmvv9JBNKKnId9/ZqtsI5QDc4MvqcAdN0qOEnP3ipXtT3yk
KoxNtAFWTbAMjTp6CPDAgaOCocx10jjnj5HnBfakOE/k8oszwJKSDuvyrgpJMTr6tGPovzA5zcnS
AWMMlHV9Y6Vhb7TMmdnO69TbKIijMWLC2DKfVQkDuQBTtQueHScESnWlutYhQ+9fY+KqsvMisXlQ
WbS7W5fsCU2+xKK5o06QGdbRUtZnavd1obDluFmBYYfIldpO4yzoPalu8ljiskeb/yF3wINQmyTn
rdNSQMi4BcjewD3nZkaAZryet/NSmsB4jgv4ZdTol3aAYxP09TvjD7srurCRejX8d4npcZGvBXQR
KfEzgOPGR67GmhEIs1WZ23lAK8qvMngREsTgt9aQcxOYG4ywiAHcZa7qiUTUoH940LwHT/D8Qov3
relz/VU2cORY7gKdWpTmLKuy9cZh/Ot+DEsDYj4qxPYVPGwQafIkycpTDKFJUBZ5Li+4Abn8VjwO
dZ7OYTn8fZCT5lLQe7w0i8RQdmmYxot1XR6ZvHPL7iopNAdL3Syh0OI6cYDd80j5iNBvjVexO0re
gR/Eks8mMMErKJYQPqHRMbBk7noO8A/GzlEyGD0C5vlhEk15X55zjMVmFrJ3f4Y842+4PgmINCap
rBHNq584rdL/dJSfD7SNc4RyI1EiCP3YmgQnlqBdrOONstcndImqRVBYIxXm1uRqQgeZ05GJAxn7
K3kTMQ5slyL7465tbnDIhwVzQNc5jYyRTgZzm+3fr+kh3E3gy8HLI3WKI24qDRqcnftkJwDr5QcK
MQLBjZHhOTsCCDk49iHV79QtUbPOwry7hzVCgZ5tjSsek9kRBL2WGd0BhvZHfaCrbislmThFZ+x/
3beuPMOhug7Vg3DOqneUbchGNuHIQX2/2YSy2h5HdblnwczBM+TXGszgFUtCXgnYXGHJCouK8vbR
8OIJidl/XCqK3ig9G2jEz0G3Owns7UvfFj66XES1vwlP4hnGmy3y0/WO9uzcctB2VPhz+xbJRIJu
0lSdQQmeYkJZKNkKpfwPr8SdHZFQ409S2PQ/nxlt/Q3hiCyHv9xQ6p90SDXB496rhHvXRmmlIhoq
xq+osUicEezCTeJbUOkc6yHze04HrxhaeyEaE8Xolkii1JdS0eKSpFo+ZlVkc/d+rSU3V1AU7yY9
FeoheH5Wm7yUgziGM1WY7M69MyQnw6XAwP8XS7CSGgQrSdMuFtpwc1NJBCvsK0KTK/0X03OGywiO
4k87ilGUb0QcQi6E0cB+F2V51BedCSkYZVlUliJDtliOAey14maPmm7mQaKRAYe81jYCjiMKu/sL
3m9ILjES5khy7aoWwM6oEi9pTxr0AD9EiHC2QETtls2PEhhcRBmzqWeTzi43mA4TJvfK7gEC33Gr
xX0QFGgyH7fOxJea4CBjZB8S/V2a51LB2H++dQTNGLKoP79ElcBSLfrMhmmIolvDd8nA0YWfUbuc
kbFexPlRQFhOBHPOrxYeQXACCh6KkLdcv/8XU5cjcE9+UZfzodHiYSsrmniftBlKuIVHBmlf8LeQ
adiRYCOomwe+Olejp9Lof/uZM/UPmpvZ9zk1FubemTD1XmBZ6BV1cbMncFpQ9by5FNSb7EcK9StV
6c01+wrfQiii1+BWJ7Y1h+ADyeviBj4vZMlBE0dpZrO84tA+7mJpqMBe05LapjDDZRzK7zL6uWXL
q45W7VneglxHAOIR/1d5uKI4r/6EzdY/ZkLdkWWqLgcpimySPGV/vPFxfM0cwOzmopbnKam/WCX8
0/qVa7Hu68H+CvWF6JMGePVmX02Kihj5aTXg+DKN6qubLAGN+tHd/LM+9kvURxykCoGVMxS5V48u
4KMY7fMOQ+LH/J0l06G6GVl7gxSnGIUbXWD4mr0meBpkhrbz30Ldh69SoqPhHNjon3Y4iYbaQc+9
i4Jfpx14RKrX4rMfKEdBUkcg+xAZBUlVzr8/WcKHWk13qkEGVijKJcT90+12PoFZsJW05/yQwQRJ
V/9RidvCxzZO1WYxxxjM503DlpmqhOyyr/bPC2WaykYjcsC25z8ZWO/rXtaIklwGJKUeuYILYpYO
/zFIuPCf5Po4GkGVZxnh8JzFuUW0dCZ0pc3Zk/j6soSlsvs88RrTcYLONEkOd6+aEAK8lS5a/JPA
DL0iAmef3bYl4LMdbRQN+2boNbNPpmxGJ8ZrU4Wvv18nIkmd9AiR6F5uA933pdfTCbVScJbX3TMY
z8iO1WNRzeposFbDOMyR+rE2p1ZRNrT9qLupP4bYlYL3f28LtxnP3k8PE5cR8WymCk0nu1kCSxFe
ffU6Z59EGvgI5p6/KhXkkhtzt/NO142KfcwlNb3JZIs6lv4TETHxN6gccuvmqTiuClmKttwD42YM
LSHWJxb60sm4LgCqPNsl1Z/ObUe2GEIfrHmI1Hcl6z1rEPNw3okLiphn6YIX2saQnwlASoDq+az1
igq2pPvR9e/wz5f5Zh+d5WP5f9QETRuYWfj3m5pA3n4YBr+VdC1YrVsdy6QjVIY/3WCW8IebdaA9
GxDA3+x+SyoDZIjR4dNhSOp87y5inCU+t3EcD95B3dx78PJyeKW+0V0As5CM7hsvdK4rHC7fpvJl
ORU+vC6DXZfmt5N2f/lOIgf3qeNXGG05qtABjng22WmaIZjSpBARASzx9treMQTzalYLEe5wV261
z4ZpP77MK2NO8B0PCoUHQivBv9qcKuiEfAR0YP3BwvJ5q2WSzTQwaJ1XmfuJ5b/1eTEOLxEY7uRU
K7BZ7Smkb/YSVjMbxDVtaZ87COkiXaCS84f0vub4zMiPCPZiz0+ZPSzDbhD5CytFXFS9sn5IphiE
3P1F/Mls9eP8J7waRg81wGMubvynQiva3sM6TbOVdKPfRQ/LsG1p/W+OCmaG/pBm+onS/DPYlMWy
ngbnFQbfj9AJ2CFuBE4VSunq4R05TcoysFtN9XRqEy6SctTU3T+k7E5tqWdnW3GmHV89xQk+8+aL
5ng/0Q/rS7+nn4woCDeUCKBWczIKKJg37jVFXAizuj3Iv7iM4EATizWlgv/KabnVUr/O+c0ldNU8
TV6ckVREeU6SmI5pt+lRzMfzohIDfT0SgGK3YBm9LnxL4HaDUB0+tgsxd2BUssoPBvH5fqKAIi8T
yJtvtLSNljXDuaytePzLJFQPf8v4rGXCtlWmu2oZRVzm0KudeyBz3YoN9YCL5RVPS0U5vPuulZX6
6LQcEBBfu1XryU/iel/Kki3v1J6A4qclRgjKMR+dJxfWOtEXG5azI0NscQfXVW3QbWVBbh1j9471
1OEud1vFDTnsqLVrOxTMZav8BJNZCoLO7HBUrAsQIFGY4VjjFUvAEHA30ycWsH5JSeNYSKNFe+nI
Zczm0AAl0Rutzt7YSv0zFheLSuMtcp/eROUK95+KN9gN2dsJlQeIvp14heT7Bnw43g7laNt/k1x/
2jpULx3cv+iU1SjpPogIreJKxDJ/uv34VGYSwgr6p8zj6/5AUarPVKk4HSZABmtYK3VVwK+Wh7UD
sEL6lmeX9HMOUvDA8uI2NbD0w+xO1X0zw8ialp5oFhAGSMQym0k07j/ynkHCRSViIraYibUXV7tq
0sxqOM1mdJL9QOYKlJEPe+j4inXZrTdWPtWwEcvCSmyPKmrXkanQ9um9y+6tneJlX/Itv4JNgaaA
1TZShgzNdlH7ONBX7JIr2NkiKe0guxU2EpKYjoSeWSMTHsbaPnamD8M3dieF6tEcIeNa9HRiVnbR
YrYA35n0FHN3LIIlkiACTDuVAzyjCCc8SPfLVaIUEUVBnSEEZp7zvLZCc74CNhnIncvje8Iy33U4
M57ajehB1E++R7fTnhYIs4NJxUNE9K10gGezzeJy8plYc7jvGV2zGf+JG7A/3mGiksjXxMLbmgIi
Ajafz5I6vKGcF4Ja8M7DjTNRE9l1CkccFKLAB1D/MOVRNnPL9DotLOePJhNzjxuU4lYp15s/dTAe
3Wdc6WMAK9myeSpTROGLMPHnYBuHFKdw7VUIc0ej6cFf6YBm+qvhD0RJRG/iweK1eaOD9RbyBujp
bTxB5tDvK90j7LN1MOf3makrfCoKBXZvrG+iP8HEVXZp1H5YjJLQDiTaJqK/YkvBY3HQLGfZD9WR
alzV4qlgG5SA7vla7LxUCOrwprQJELj6geqarTCfqPZ+buoBnuPcqawMWjhEZfEFoNKJHXUGbzxb
xC6kImh9iRO2L+ERufKtTpRe9MPA4RkrnFzCVGQCQyTxQRmkEOQKhhlxBFY8D0uTu8AaiOuN0v1a
fYD2wqpbTK95nroMFvO3IcSo95dC6vdhcv3qbFwhegDGHG91/x+/aYBVMapPP/DXI+2rIXl4W+m6
qi27dyZCycmdL3fH9nQ30oezqqqoi8xJDEK8CiOTkXKlgBeFDYF4PhWwW4VNRbnHmcq0w2vyHevl
QYyZxQC/qa3F0UypOqQT/1VBdlaYLKpBwlhwV+/wC18EyOSbTuG5/9uDizvEH54+KT0Sf46NrHbP
PNLJehSePSPiyqlJ/KQE9vCnQodukuU/m3vrOQgXpD/nMd31mvhEp82/7+K54Buf0Dth062R+yue
2H+eZnBS69e6FdYMbD9hM5v1ejSUtdYBmlV75iyyn52rxNy+AwfdGUKkG1UuVs5lw+8OFSq07xtM
p5chCoq5XmRqF7mAo1mPHr2038GVqcj4kgT8nNyoIy4LpzG9Yv9Ntp7hHYfH3tqr2WIYqqn+LB3L
/ZM9eNJSNqe8AHEDKwvPI0sfMyT6nFvwx1Efor2XHNIlbEexWXyefi1voB4V4nIh8WuXih3BehGX
4GQl/QzUKlogmcbJq1Wmk5d5BK3KEl855iTXsnwS3xrlEPsKj06L/Yy5C8lotLEfIbxT9f5IS3Uh
mui6wnVngC09ix9D5+viuJXO/6yncFFckTstexY+iSvOyFgrVt1U44hntdqh/SASJD576HyEhGNf
rbVFbw799wVdv3j83Jy9T2Cz2/K/p8w1vF0/oaLLa54+6NF7lMywMwg947rbyNX8xccseFYeNf3r
hA11adg1rD/5f42OlGfaS8HClFvWCytZnSk/xXulVZjZ56Twnmi7s2KQpeGyWTziskgJAaG8ZiSE
wHLjUBMPh8Yjhf4ZIAfwrkHOrDpWkRk9KRiI9zS2Xmyb+8sY82ArFpZ0ksYd/hiBEelVra706yB3
yaLsljyt+p8hZ7Ruw1AxJbNBwOm01/vzFoB44QkNUAmpkQvk4ZR4tYDaoIHHKmtd+/CtJeeR0HTn
86bvDOAWk1yx4C4jutJeNPbV9UkSjUpVZ3CNBldXgMHuiasunx283R/yiLWkJUtYReB8nm9rI92h
lCfjjGgw/8tcU4iJ6iMuJhWC1IlIBw5DelUBM//Ewc/zn8n420PWIquSH+MeuVo2CQWtLcwUYprh
K01+TxYcLgOxemKlAJHFxbpsErCJDvyeIwSEOprarFsQeVd5FZtRcRdIa80ytEI2e8RbHVR2WcWk
PFlcZL7cmXHiv5x47xXWzkojPC1T0eDu62qPXcLf4k/OeRBtLneYuTBpXU+IESKyusWCx+d5duOQ
jML+2g2Q9ET37/zpG1UWPiu7SGpTHUz0PhQM2ff1N41S0+HDcUoGzgpfrmLdnqV1O2jCkLZhQFgw
b0Z1ZbrtR/PlOQS6FVVjydgUBLfL6SpKRIE7L/fDngaBIWhRrQ0HzmFIAsRgMg6wXgMYTqpijbKg
KgNTi6i7NUlthbXQhUeLGgufmX6NHmI8msk4L2ikX/I2ZaJ8Od+y6swQS6LKGtPK6+ROaLdAUlPp
hWDvRA0WkfhIwqDG4JrcbbTXMPwFGYE5QR6SOq2f9+AltkTJgZ5gim3/UE5vtqe43v3re3O9F8Bw
G4wGqatGX3PkmcJkI9glrF9VVZaN8N++G+9441T5lQEwb1+JZlxsnZk4XptZLpSDn8JPTtCs/Clb
0r1q+ecLxoIRRmDj8EtwbHSklpAKPrPmAfaQYaddJCNnK4zEHyLYv7pw6bjWMyfi+gHhPz3Fy926
DrSk98nFfFaerTRNJCgjM+Q4SCiaX/TguEVKMsgDFMGN3o3oub+ZN+96Y9Jmpp3E8cLf1WObzzd7
lwzi70n0yaR6cO6uV1/nRDQXcv6UcS6d7t3GIE/qGrMB52GdS7rG9wpPOLN04GfLDQreGjhlHmC4
1CWJbYuzQtHEa3vjn61Yq2U21vJYyMBClQ4Vyu/RyGXl1PbXQ8tuuVR4KknytvajjBHU9zecY+LF
9NqHvmKBEdQxaKP3Zjm+CvuzV/SRFopbrdf720AiqVtHEqJlHyKJ7G7b87RHFggxIZTRv0Lz0EJ9
UEDXsCg8ZdzVzS+TQ3pLdHaTPDUf9VFnep+v/kv/Nv6zJO8diOVGixsrNSXfJFSyfYf2ZnYdApnq
GdcCEmeOBxdTUA71rttd0NhzzpJaj1HweMAli68g+ze7Q6Ao4dUsOAONNtJtawVBic1uKdAwP4se
rRTduky5KfLHRDZ7UO4XMm94NSuTfxFyOnW5TrU1maYF32DWPcKMQZVTf/Qh8Yfjva6iP3g893M5
jMjhC7GtM5QqTsz+tgrCEZ+dXAyKgkRnpf40yseFTlLzyJMZoyzN1IKZ0sALKOd+uXs773IAw1sy
ejlesmvE4de4xdUB4NBMc+OrFJRSwephdYNyi2ecPeu4P2WjDXVhtBwbGLj9yfdWDMRLNJBi4VL3
PUIISJBqDqFu9Q9ARoVtha2EwiWTbwV3L3vzKTwU6Zkv4+Jkt4RdXkPfHvMUvh45lpdikdMsxqRm
6mgabnTNVQ+wisybbJvfaIB1x/2l7DxlsDKb6vUzvZXjiWEaQt29o9kLEmMTcgiszSLzfsgo2O2I
yiaxHxV7nmOJxC8E7nzLVQimihVVDOI5LmGh6Qm5zLJj0ZPLlK0V/mEV/a/mFNkzjSf9owiRHKTY
ZT0mmvxBsdEPFYSxaacy9L0S94+PVk1eo3SuGGXe4kkELU+/f96dkOpUmGpjmpFZIBkl+tu9uQOB
4KIotrMs2wVyNpqKlHzoj+TUZa9jjrJblhuhduUd0XlZrxt7VjS8bNrsbEZqDK/26cVvMgVWn7N5
0qrA9ds9NfS5llMhiMDMpAU4+Qrfp3hT7bErbTvFo3M0MKxOpf58ExS/7IkXUPnj4nk4Zai2HDrH
LZqlTo9CXLIVYRHNgPoPJP+vxAz0g+EDaDStBfNg4RD7oKRBXiLK2KsKO3o77fD6Un0dF/FLmHb1
qp3ZOJhbyhTFt14cFLLOKP5Sp1kj9wA9QhtkEAcEakOHVFaRvGImdl2ObfH8HFnZl8pRA8Bddqfs
Sz+LeiV+1Nb0OMBxFm1eAl0hAz0x0fTyesfvcMdF67XJTG7ENOL/gZce8+RIbaLXpLjZFrvvWZ4S
+NReuiD1oqMaNol3LXCYv5EZ9ei3XRqHuSe/SLqywE3EqVabpUuD0u6VFNUqvLecAJoNYWLl7yAX
vapvC04LXQWXWd8EtS7JX7Y66c/M669eS60jjXU3dbCq2FwvtygfYW+cEtWQ3O6Yor+9e4rLlohn
DR9WGpaNshh5bCL1Fic1388Ehtho5Gax9UGQ7Fgh2SSVpE4TN+EgqTrDIIdVFXypBAXTJo9Wgk6m
5wTq5juOTp74l6oI+hMr4Leu99dwCnPJsZ/O3Ck09e5WoTG59GwD9YrO6Ml6tnSwHGsnrbW1xPxa
QdOJqgroAxUSrfZYMZKSUimfPulbUGigoIAxjaY1m/dbwrfkhZllADonoeIevVt/CAREmWyskg8e
ayaVQJhIJJXraEles7nq9aQEVZYKAelBuNUHgppt0vmQ1YqxfOHjCRHNMn81hTkldqntdEwdAaNT
ddaDxQPGmyxUza0EOmuxAu4NJJs8Nhd9OtkKHHf24bbDibd1W0j2rWuJ0Lzua+qudWXO5kYNIOrA
U/d8DnsB2azkvG3zqE1PYg793JvI/sUp/Ap3iUovvp2DvW/bV5Y0+kLSKEiKQJVRIyVmKtcEJ/W+
suU8LczYMhhrL5XYfcu9YGT96ZdvDZBZv133HTjvmumvCxDFkd8CEtjiIWk/HieEy69KPCViLbJP
eA0yyHkaJ7rEz+nhB+wtO+FnUCpYv4bV0R+rJxvUA9EiwHGiTZvWpWXKtTe7NKM/9gLrW2tVOyDK
BV5wte7j0wuYfRxIpSCbYdk50jnIjP/RT/GsAxvq0HtOPVbEfpaUobDQZjlksgKHeMEZfeJQTEhf
0+nEgXSN7eZENDxNwgD9p08jFVUx4VqytGvLAGG4yqdPf1bZC7lvoIDzi5fAQzwCF5C83JGY54H+
G5XDHB6kn82OH9yT1/zIpVrjxkCYyNbDNl9HYCiFyh76yw2U7H5W+l/e0gG5em3Ib6sr4JrQ3kLA
VFO14OdxNRYFStiiSDExJPwHPeEnjZJ34bK1TQOfwnRkxQxcXS4l49lF/3YVTsfEWotJ7R9x3HAr
6yRHHgSsRLBTV0kgHlOYRMbMEhTkKKdlRtSTiHwejpNvLzxeRQbghka4PE+rOaGf/MpFiSArILE4
XhUye0qls1cfiMGBVHysjCGVIMoT5K4zpwTbrZIR4SGzxivk+6ocegFm7Z0ddrEufQ2gf3V4uf8a
DjlXyPghEI+Ls0bs1xoiPzlCgR3kYAyHoUAp7Zw8TDup3s+y9vTvMvef/gJi7ZmJqumm4Di52hqH
cfxLEZc8/DX04YvjtM5euok51uuVIB3RmN47gqWzN3DbfGqTm+ikAqlidwvBtNsbwmrNyK+6YVjZ
2M/0fYmfVQeWK9uib+67hUsoPg5qkeRxZ6c9+3F1Cx/pGi0Sd/eLtGpPvmZHT0BWQPFeF0k8O1CZ
f8LoHvhLH2GGBbskheV77arVCZ+g8Za9x/N/9WLKVGH3FmOR+Yck6MW3S5l6chhgaoo6JRpfWHya
nEWM/U+bimZYw5hSU4Y2anBYJZkcw7M3l1CG5NAEfPykjCh2MvIzvEJ2/fSEZtX08mkXO0adch+c
uwr+2pbqO6L4rilI96M8LnCv4CshdzgvxbLkjnHVVGyioEjpndpCGKKTVs6ZAwhLEXRbedzQ2NLc
j0Bj3rLsl+ds8pv3LM9owGOSzcAzP7rNY0iWqYL1LUlwnToYs1ZUe5+nnmqFPf+TwemGPHMXPkHr
vkhl7UgzqdnKF6O8sj+TyjI1HrVK7g69z0yxwne7A5icvJq2JgWMqGlAm8dYvRlEKlFIKdhzEpa/
Zsmv+C4B+/NKdIVI6Uk/TZ89dFt00LDE1nB+pZ24uAaiITaV1dso/Bx/ap5R1YMtf7lXFFHAA1Z7
eq/QseqJrLzbYqrRgpM3zoBhosYDh4aYK+lrpTAwZicr6dcEuZuQY4/LyWy8a9Di3aAfivnQUbLY
AWaMk4/0xxEdal2Is8fsMTjWZhQk0kTno9AsIYWlX0k443P8wtaAtqZEjraU4xUGmyE23u/ZM8sc
REeZw2lYDaP7DvTujvCoE7dlbRAZVXMYrGiJqu5/qDi+A776uinSeQcSBszYgETFxa7G2E2ViawP
bp/q/K2VuyRcsbskIN74GttvhDecXuZvna8D1ysaac6+0mDtEou3nYnJDEOAV4Dy6dC5Y3f3Yo86
xfoOyK9XlgVn8wRYRZ66ka6OfG9Am9/pptAZ6G5niT+VuMb15/77wQPdvzTDckvaLL+PRJ8pFn4D
lTUmG1T5tWKbQ15iizZfq+XtLQbuA8vF9UfKbrINuXDR7gJJKTDKQ17NvJwbXnTqtuTGoNRTwr5j
I1Y9kmW46Hu1KfPvPVCKMJRKDdvOg8S8SsAm1SEDhRBUhqhwmFSEfQ4wZYv/BYFMUZcx6sIltbDU
GsWkiqKDQtdNnF5Pp2idRmKKi/fnN8xn4ZUp0R49DrL28MeLgBprnF87VI/cX+k1NqPCpsopE6A8
CKB/+t2yVZJa0SuI6i8/a4y1aHVlKJ0uzDXJYymM7yDlQ2cAHSYA2UxVA68w+ay/DXL0qfBVP5VT
gtSGss0yHr9AH/f2EHkFIQDKZKOaJ60R2Uif719zE2r23HtO5RMJdaAUltwTK2u/7/9vVUqoSENh
jT8xGccJETXV0RLW5xN5SHv6bE4IMuGEEg4Y8mdjiur5WphRYRInDySkFlhdRQfoQ7sO/FxEBtT4
h7BL5mz3kQ8jnIt4G7YmlwpC+OcyhAZz15FCb2X3Rb2/zmEGAUt+xNmzTLnOCvmmBk/yRf7cORx1
wYLeRKSSNy9k714ZzMquGzUFYR/l1yPU1gboktj/y3j5xlXjE4Oxiz20VopSX1J/siPCynhO6+9I
EIwXUUk+geSon0U/xCxBoxvOxW7amtJmUZLV0fGkQ8lV7xe2TdBxLSoPJFAJ0gWKL7sQH+1T52Fk
VHFSBBiM57yk5bdSxh+yUKDTjTRksYCIpGj16Xme+3ehoR68hFTAzGxTI2Ab6WpIEzlUw5GJMOHa
Pms4pLxfPfHcwAIH9A6HLfseVOLku5k0hPWGeDMCs3QXjsim7bJkR5a0swngpjLPa8s+9Z+UdfCb
LLK7A7v+YNJ+qzd145KY/dP6RsBJiQDcGayN5Do5JxRHcvGK10796rmhiYlgvzjNW0Gv+FlpQAq7
PXzSMv5vKc5w37PDxn3PVjRmAjPqzqKKEo7IyGNJ8nzb5U+c183Be1OyEZt2DWGpHBNbctqWjxD1
vltXWoi6mp72rZCeu5BJQ2/F68YSbG2SIhDuplR4bFmiK5/lLHTjzTTTYsjvwfsOBoiO8gTtppPJ
+UdI5pArQ57fgjJWckoLlxwdArCuJafu6sz9Xs9ZnGiuu06O2EG0XZeDKqNFuSl1k8Rev4KPSNAd
bKZFbmBtGgxGOkwA7HzSoxssUMrdS/T6LGtvY7DK9Ro6HP+WnU0BeTwLoTz4uFXvKRJIx6fhcrFx
OKvLODMbSdCleC2FXkN3RGXi3ySB29VbUhXs11KCnLgGwQJu+/EkEdHuc0YGNwx5GUffpUdZQUuA
Im//MeOtkXi6ps7hjhL1/XhoRWLpo9NMd9wPznaTEMQoivH4QW4kC/EC3SZjEuCoIjDBXXiXg9tk
yO4jQ1Tfb6+lCPgZYpvves1oq3r2oi+l/vZEI5q7X8ZJYosz+gdQBXLr0ZO/LtbbG+4LSOVTYFM5
55froXq5UAxKdXaTFrbf7hlhfAGR3bNNwQlOtaYpZoW5s8pFKjYJVgygnrMgHT8xCglA28ZPZsBd
eeBPDXLgGZP1dlyx5RhuL2/Ayexas2leNQI/SWPgHfL5AzJDMEG3U7IWRXmiChg25yuHUSryceLB
yUlHtLiPDmFwKJuY/NqVcXykyqhJOYWDPFUG5t6moxA53reXhepF1f3+eaCrnPA7ORk+/inEFtJ0
k4RqCdbmpqll+i3wCIRaj5wG/FKW0bBOhgTknOZceq77ReaHLbuoVIaziBL7zjvsd3fS6iAR+fh0
ms5z9n3iINjuvJP6ibmEh3PcJbymlOfqUrR1sqxZIL79Am1eUtWJHk9U+LJG6oIUSqkMjdia0AII
9LSzsSSRDjBRpjtdUUGo9TIeX3NApgtsG/2GcEoh1/jyoSAYfMX1MVmaU/CwLQH7YFwovwS2IpEc
ppkDdg1dsgg84ZqzpfA/+DtHWWwpKVMfO0QwDal+dlLE3R/sKxURnXg3qI5yp95f8XYoJl7DTJ43
JFoywoEDpMk8KraD8ZA0QRQtenLVg78E1U1CBlVcp5i4FPpzaE3uWbBOA/4f4Qzpdv9Tc13bub5H
LiW0mdclrBalW/GF1/MOveDC6uN5t2784RnA4ATSLfvbgBxjNozYuh1DBVE28DWmoohYOxhF7mRB
ZEv2Ezex0gvjhslNMC+jjiTBIdvurx6E0RE/Rp+ab5wmHLefwEaQfvJd/OX+kMNhoeoiieF0JYQi
Qw1emrv9ovol/yHtQFv95KDYMeCazOTjywGxFzBCNgRUPGEgEjVmmPkJaMA/DKIovu8QPoBVxSxo
WmCI6f+hU6tAUe3BeiiAjZkONSsTU8IOuuf4khU/WvbOtKNFE9k4Gvw8q/3v27CkCmFMMREuxYlE
TAaE9i/XJ/eaXeclmVTWtTQHI0d6vjshPn1/Jr/86ujR5/NBUXC4EQTWUUjKyWNVsmRjx1FO7756
d6kQNm6gZT5/vHMyJIa9tZ/aHe5g/CNibM/wwwkdH/n10dczOw7i35QMvmIepJ373oN793/GP8+d
PXpio5p2zfUlJ1yghc9zALyGhOJpKAbABXke40UgHZLKYQ474mVDS33iX+/wZTzZoYzaZq/NiRpC
+ez2EKw8/XBDqqQnX8CN5jaTn8Tuth1fLZCYidqEF+3k37bn4VWCTGfDGtFxf7++3bO5i8qIfwKt
1+Hb+cZ2hOisxxgR3Ii+YJs4GCM55I+iN7bxnyQDpi46TaQfDQXkfNRZaiJvBuKGWUmMF/lxF1ts
ekz7msRn6w4uHJFTJ/hv1fRl0MowkVEGTSjJ/dVGswLMmFV//BJg5wu41SZ6frUBEiNghRBTHKQe
w2m0YfQqj5BwyBYtxhmcRlPpAqtWNnyqEzIhWF/U80M8vMQaUJmANhixLWiG1TiDb1vvxKLXKTVj
9qbJHK46fIdgNkfrCL83vRei2pQ6pZqNSI9CS2tEEVgRdGICg6ZN88Pt5UjvQMKYZiAZYq0Mjlws
htGGJC0iJcCN6IsSs8SQDMTS4/D2giKTT9Rw5U+2ZEz6cWuO4tTZy9WeMdY2ER1nVJdKSTeSs0aH
9mCrv7aQ/XCPXYGuJPd5c7Py6s8T40abpRwlCz95q45AtuI+R7mkTUvUvt7wEizYuvBRMbiuOGiV
V7kT5+w+u/P7vNAz8tmqu1Z427bF0KHhka8g3MHV/l7QRIBQghSf1YKQnqE97PISbWo+Y7lN0jAp
BZAFM3QG9pKcSbWC6xB18UDRVp66aQCyMNdM5169zLt8eCNd2tjtAt5E5jLaHmaihjBMggepZsMP
v0JgzEc+TayVjGbtus7qOV+CWnB3GWpRQ+kE87azo7e12wvi3Z/Ok9QeB9GFBd9iAqRQnor3PC/n
BLGBiwz3AvvKIKmibiH6KPW3NONako1khvduwBcZeNoOUtUC2Elr+4GQl7fBnl28kwLxZnMoyhpk
G0wf7efWkTEBc2bWP5w0I5LrYq/RlaC4wcxCWUAe+IndWHjs5H1w2wpAwwOPvxrRVHYilI6nBogf
oGgeA+/vY1AjI0G5H2t8NRXW5xMewtEe6GKgtJI7E1v1IDBvRcOkPKSqFAELqVZnOB+IDcZd0eAi
LDf1ZcANjByHr4+cPkaHX7IRfamqhkcrTsyLTwKfRHR0wrmpN0NZk2Pr5jnqhf2aGultvPxo41ay
nS8SdHv5FFWurpYdygB2MebX6pGRDVLAFBVGLM/SKiJtTGp+SbEwhhjUtUv4jULeU9mS4YtEf+sw
TCJWOJ6aQVZL3k3ntBsk840MZj8EtNV8/vMah6MblmyWTOvPoTCPB99x5K6qM5/Uwsx75I34KmmB
PWdl4C69/rbVCMMxYLR5w9cx4hPbXXXRWQdz6Y9y+K+hXZg9Ko4jGmE17o79vqsg6xOzleFobQdl
4jVL28NEjef5p1CCrc9aO2E/FsuIlJ56rX5R5mrhn8YIBGWuKWX3yQvh+sXTZ3zf+BaQxWXM9OVg
DUJvGOPbrFK/xYbJArZGqYi/+dKjhOzJvocoKbV9NmTupDt14GdXTLnG0P6ZAqCeQcoDHP1+ASAC
zgUs3TI/grKF7s6UVLaGWO/2wr+0DJXhgNuKG7oI3H0Ori2jjFVthHJ4wM5qYqNk6zL+JhYfzh+1
nfraevAWDIPgx+/6TPnI5tVF0XNjZUOBMLrYgLnI/JSiu3WQA/aP8LZkjH4qyvrdFdna/p8l3klx
pqjnn4ByVBtnZU5waoKgfbZUkcNSLOc9z+lw9s4WyQG5OFTV7MpBU87gJIznwQTVQd/6rSGhRB8n
gDXhL9zL4Mp6V8+gQHTPoQKOoFq5TiaQJkFthcDqINbAuRCYqzonjUe/zp+aUPBkM0yz1Jr0PhSP
P6tTXzztYXbccERzhtDekYR6hu8ldUeQo0z5WOj3Rt/gkNW09t7mOQ45YAAX6ruowlLA6m4jIm5F
FrvI4TMa6GsX/su7S6B9NL/Gk+dDsPmacctacBvg5YrnX1krqoS0Ve23t+FBkns7XnGUDlvUCjif
R8FFNcjiQy/9+sU+o2kLrz1XwGlT6OM7PzvHz9OPfq54xnqTB8rfS4oxBOcDgzmQRFK5bKUnx2d+
dJRD1O0ypCOLWQxBh4JlV/YBrMPkv9ga1+cZkKcPQahY6dl+nekpCkqK5ocpSGhMEogQBincw5m5
j4bmv2n4DJlKb6rplHE1nLJrj7ICYDZRVYTLxd+5ViwEeI/N5zkNnCOCHutuFhtjXVnYiP5/40S8
LkxRtSz9xofV3FjbQjLwniUu50xmBwd95CIIkN3Z9FayMk49KFwtEvBWDeXqTzhtoydS1/OOFtOA
Zn8IYx6poFZ4RbDSbXqffQL3R0nHV5uH8vxgvt56MUeCAsbHVOWcxA2E1wDbNl9G0Cl7HJ0rkU59
NC5G1PWigyBSv42M8KGpWiEaHdZX6VEwbwGCpAIrzo3+Krn4DNw6R6Wt/BD0jmXiHazGBL7dcxkb
mpA9OpPg1SCfUk683tBnVj9bhwsi8U4FnOSVp4+B/clg5WcQo7stVGdCnH3filveQrcjfoBkXKuK
KUn6w1pC9HB2rvcO49rHdM6PM/kw9ZdpldhNCDuNEdqsIuznvMQzoJZo9jiJ9Smo9Z7v+hpsU2Nt
4tgdDMRzRfWZvgehpq2QTpN7gv6Bk559VagB+XH68D58vNN18Pq0pWmfJGZYPQcSx1xaRWFaZpiK
RnrWNFuNZG52xv7sZvT1HGyv8y1IQK6XSGi0ViYBa12N9bXlYF1M0AK/khRUqpOnBRLpRiTVGwp1
SHY1N5BOC545riK79lFLid9M6MaJijGAWzD0nXviWz0G66OrFQLGyZ1YKTQS7rzykhuHOK79Qf3v
+z3MBr4Adv3nHWERbYfuWh9dNgdnJSAPwcLHWHTjUzVATCGXLEKOeYXsxmoX17jEsTCuR2/XBaXU
+7uTDsZZJrLZUDj/rK1tLw8cL4vR1bM0azyEsFdqf9iLKEx5WyK4Kc35k5sIfOfympAqkGb/+5Kl
ejtVqv2kiRj619g5BkrzcRjBCiZdA8XEXDktbX5ZdnxsAMp7uNiFP6T9yiNreCaztowoPoem00wV
gSjeWzgljl4Z7h+ZcGF4AH1bmUcydx+jA2NpKITLYyJ7h77F/6AYJRy6NkiTIvWGE4dWiGIJC7Sm
gDbcY56zx1FtECzBCHTMVEkjfHfw4oi3sjzeBv9digmYSfayxnnsxc775+/hx7W490S0SpVon05T
1ttOwRmaA78udni+d43aH6HzXvxXXZO/snARAIo1W4twZmuYQzjKbcQNLaqvQla2ILixdiX6nVR8
nc8E0pam7MWNKFWgp3qKilADg+zGzl6xT+cnFoAfk3rIr/CPA4E5Xovg1QjQjvAK6gs+szAJAhnv
dnohp05LAiq+HLTOzWTAGUSBrqdXndCQnfDPUIwfK/M+fG1OHEQsDiYZprpMNibeReSGuwooWLRi
Co8PGNGyZHzZ/K4k1EDCyZl5RbzLVE13g7SpY8k6kj1tDoNcb5ioRrsDQuhyYyCp9fEeBWTIigqm
IgSWO4ZX48EPPmZELpiTGujiqQgIJV/x9yN9MaKlCRyXwTVFjS70Xhd3yJMVRjPLbmK45Mu04pQv
muivqWaeQvtkOCS/y0v2YfMbh8r+OYnurkSOIqthwQ2XNlvd/uH24JUfLFT5AMGvNQNFuSliAo9n
0HCEbWWB8fa+n1KDLzDTmqv/31pQVGQ4J0w2vyy0gJ2igAY8c5SplWLy15Ubv4LuOX0mICk9AW7x
+zIPAN7kfSGmGM1r6Rd4Hdo+tCRT6ShV+XizpfZK+UQ5gc+QTU1L8Nbf8QQZ9o20UR3mi08uH0Ox
HbPsBSdGrwIydVBm4JobMoOz6rZNOsMGBqc9G2tKFPde7UDJ4GCYoW+EnncZuR0Fn735+GG31AOA
v6h8Debq2FrDpUOSi5GgaRR68X/d9rrHGXoN+0R3o5CcOZq5vjYlRd2FUH07PV5hYECPLp3iPkzN
lqaDvP0bHqFmgtaN7TzYpt5eDtqrg2Q2a235leC28a3EjkyM47T2IqvK3N7sFYeekm+UA7cQdbBI
3hmW+WXR/fzxdqA8HQC/96ORsn2PcEPPqPkOjXUNGez6HqsKUIfp4R/6UQSfBtPic8nkB72/auaz
efX4wcBvXDAaHx7KL2WHmqmR/cebEyNZocYBopLsh0DJKsZroPSTvNirO3VTcQTjK9NWyBtRVZ+y
+322WJkWFFctZxzCrPGYc6tyqzMkxYJlQ1z8O+ma8Ze4OzyezVVbOJzwlxgaTVT/2yXHYJ6UEvbI
npEErS70NDfYhAdEsrTaNV2A9Rtd5Ud6ON8E9cz03SG7XRRU/64iE3eC7UMno0fc1NpCYWi0ANTO
dVWs9Wg7Do6w29PiyVe7LiC7FxxBoMM/gw3hZJW/sq9rkovKkDhrytZCSc0jgcKi0vCQxbgmnPA9
n61rwYkF5R4haLPGQoirf/7Mv4IOgV35cffBg5VVFRZh7ESPYBF+3bIhuQmrsUXFhc7GNRXXoM46
5Yk9wBc4CzQBkaWjXOegaPgIU+wvIsqsqpbSwCRXtJyJ8myjwJoxlsr+bsscqTimkl7kZ8ZF1ewV
LwciEEEKww+b4aR4lh93AoDcZ6zTRIjxmuG4w5N0/XXkMIvrIn3r2ENwp8kWC4y9JOK0v1FWh3Q8
IT5sKDIPNOAHKEHx42oB+qiCslIIKbD5/ZZi96+nIgteInvgAsjVM4bL9UVcFV0/h6QDfutH4TkS
oCAmj6sbQnphvfmVw7P6bN2eA6NHFvnk1rmzDtcJ63BCAYbK+iBd1QQ7SmU9IL4UbVhk6EhxfPcR
HjNaYs6m4yLcUUeCM7ngru5ou+fXY21JlFq8qJFwTItlGYvD9zrmNBWWxmY6BUELagPQ1Sz/PGz/
g26dad4Z57DgBRQxrE5OJfpJZjf4hSLoTzAno3rOjeXHP0FmhWmEDGWyaI5/CuZUL95Bm2Jo99zh
8oARhXhsI/uUIp+R7iiK53j4GJUGs7pZ5/KyUi4UmhBYAmMTmBrIaap+cow76+ANwRJu8/kHR3hm
Lu4ocTgRUq9gTd+0Havs6QIMNM9vUJB21xxPQKYBig6rwuUWNy5GyHPm6LnDZjP63xY2zwiBCbMi
As3KOaYfV4ER+f9FpYbbJ8M4qOSDtpbbMTL808WsmcHRghLZcV27DrVsAV5vduc5iOGQhbD3VhmN
dqhUs9nKzYRzsdAHKpLlte4W5ghvcmb8IXCxz8JciIA2WWUV+tAXIMc7yevVwrEimNL7q1rnygYI
FkIpKyxSKOzHQPrC5AbnwJjJTScuEcQNWkyTWN2DQHAuFYilyMdnxIrLUm1Qrl0uBRG56aby96UY
vXDHmb/DXpfcT/Hqc9h4lY3kkncTgp8drDjwy1h7odRHc7ReNXA5il5qxUUNvKl6/2gN1Y4FDYc4
1mAE3TiI6lLmCzF6T3alcCkgNuZp4jggMCMxCWss6Re00U3x6BADjhmTTQ3UDxb3JeB/waF70eVw
SuWwm03g93aBDXutSJjMKVTTBCc9EL1SDhtHPbr73bi7jmVATeK6bG9lKLIu+Ziiq0HyscEZREAQ
UIhoUeee2bchz5fAKrjA84NVPPKTqQBYTxXdzV2uY2Cjd2vPba32LMGl4aBUjv/tMdf4S34HKw9U
vpv6jasDmsC5tYJpVEmdbMH0v0muyUcsLsmKohQT/iuSJk0o2AYsZy2wR3u3u0UzlPyyPSCNbxbi
X8PPYYqxtIvjAkM7AWqpQ1Ky2mAz5O7SqK8WlTTBUpVvPMiIh+UIU70Rz9ves/vHPvAxlT5c0tCA
GdTHA1X673ajRNOGgkXD/x/6wVITGanFcLsUAZqiM2oE/zAWDjWQVN242yDnT+tP1S5ZAy1Rjm33
4k0C9+kS9ZqUBxoLTUHsV5raBMuKVdPT83Ck+XVHHOtNt+2nEJludlqajEeGhV2wbQKCNdWUYP4q
CHeWBLzFnZAulY+Priz26Bm2Is9mw/avdP+VXNEjKL8qMYssDxIDTklmNOYCza9W3OnasXKba4b7
H1hcfw5QNwMGpyGJqz8DI2xQEJfq08D5/El5Xe4XfRV5dvMX2EBbijUODeNIinnOW6qZqBcW5Djm
8pO129/utIS8XFzaLSgeQyoYNJ0n2YxutUUciUEHcu+ghzs+moj4VQP9wOtJ1VPf7WHju1UUfYJ1
vw7aXpHsFrmTfCZG7AeuT10RadrG8dHbK6qpXXTinPWkSndYxAZrVbj/k6T7gol4srAEXJ8jDsBf
7cpB7H2qG6kFanAJdytnJslv4k2opC6TnISSTwIbAJEPxCpxn8ZXs/kpS6NObwOXQ947h3LJl4bA
1grxxxSD14+R+Oj0+T2vpfIKgl/bHZYlNmGTt9YAwOWbrFOazHdvJSraox27pKcKFpI/9OAcNXQE
9kDcVuUvNruPLNdNO3XQhn70lrG3EP1SHEIRDvL304kvRoQgiRELYJNrQIBaGWbdBRtepjuU/+rT
D43UqLtf/Pf3YI9ZH+Vacg1Jyeshz1ChzBbyOZX1/JnxeNEWhOdb/h1TB0wW1lZEVPrXKysqlA99
4QGl9IhwjYYlKVG1NosjL+NwR/hmJTgaW6WGatfreMtHGXJdIuO/j6e3zUoOi3x8kscGuHiaLwmX
sqAQzU/hnr030gFrcKtN0Aq/qZC2xj/7j6PwmrYhHaDtlVn5EgH1QMLWkOu8lPMFGGp9HbivbPj9
TDiIpQl5n8dn9rfDme+ZIsgTFWAkndRsvKCqdM+X5hwQn2ZtoNSOsCNsFy7er8tm/fInrOPuniKf
o9M48qwfbBcfizA0Qrv4z6NaPoArfcMrgPtT7JHrRiNeLQxjvxiVvseWo8A6GjmTnVY5GxnnbPlp
i2Wt0nv0TH//nSArIzRvVVUbyPvING59t2rcYXYOr+GExWlgh6mCcYsqdWzMeZkJFq3s/uXEKlij
DCKJy1PFWa9zrcUEGI9x1j/IFq7XTSlR98p1ulV49ObFyX2FAjWbJnp6N6gbWB8aZBC2rxZMzoM0
GJVVj1WmsnZ8W2+bKi0IWpoi0bu8Oa2p7etckv5ScgBrMQTXD+mfJPHp7tUTmOUm88w5mhghp5mx
hYTktAgnf8LBKeZH/Lg+sUVYCuHOrUGCX+jhHAGUO/mAQNNOxbUsHbLedvwCw3dfgvYMuEqURBXP
XY2RKTMwMN2aMjGDs/31oZnx3p8hqXZI1cip5KaqbcF5fG+Ztxy2+C+JtzLWUZ5d6CQasSZPdOzy
dgvmHCDjxe6PXbvkngGayPJrurCPvyayfM9r0HmChFRs8nB0upafen5RPgPvkSmrbxy3B1dMdSQY
3kk2jYqSSPcwuFEDHuOswVLcQWfU5pX3TnRBfAGYz/bNP2NsjuDNZ//br3IEl2PzY68dQm3lDXQN
KU+MZUXRowL8mCRdVxaUPCW3ZQrKT65FKAUC6Z+OHksBCPOWx/oSzsOqKE+2w8O83VWrJWEnOzhN
AK3LBjIUdPBr127a9yeg4+fqwtZ6C6bSuQSQillpjN6ymono0bBTJVDAJkQ4HtL+7r7TcgWZRbnH
NPVlpaVT2poyHvgo1qR5vFb27FpmEcWe+T0t1TBAgW5KOlXndCGLQPGYK7NIbozOC3zmym0SvZH6
qvQqpMVRpqeaBwU9EXDRnH24ZJZCNQLVoyQ9UUOeQN+UP7TKmR9RdZmC4zGicAHgChuBdTBiVQ3h
q5S9oou6FktkM0VernpuGh0IUYwubUkFuth3iV5YL8yeuqIlDZcqXVtGx5Lrq9cNGDr3occn8UhB
+P9uPhJsdlOsojGNxGuZe8HPl4P7PZQ/8MRwUC2/ECO7E6LUmHVCAD5b7q12XHZLMjmKXx9jIl8Q
Pk+FAc2jLJS4ByevPxbptYLGJB4oVpT4BqzKmJQ+NlqjcNLR8Ti2wh2UwiM8pfbYXeDWMzqruxdV
J27y4yzhWLBrgrEekDu6WGpJwZNpmk487JN3YDxmi0Skmrc5jbPmDaXBg3M5UJvMRR5XMHfjHF6e
gi0AouV1tf+3NSbn3ZIY+Pgtqvy/KFRM1gMgKlyAgdmnuu+OlywA7k3uGDH8mrLIMqs3Vu2u9fx2
ezbhuRNeAC0cmJWyD4FwE7pjTRG/s1Zb27RaMmVmm0gYf2VCflpTyHFzsi1u6em4sL+/CLEKnCSn
cNtDgY7OZTHjYgtFycmsFLYhqr+lB6QQhkZ2+TTo9ievhvpSyVu1EORG92iB8vbnf7zj/W3Mhcc8
rM9UYon0Fj39jrw7yjXnh+55I/AOwxBASDVXFYGPSA4ZoONW1qVxbke0aucd9Ud6pNJE4HSoip6S
l01caJbIIuwGJleUfvUEl2YhsGE2r4XvofvrLmZwptFFDbkfZcSYkE5iTtBpeZl8apik6brfqiJ7
rn+86tsTkvh+rrGP1u0G3ghQdxNRDvhrdxrot+Hkkqc+Zk3g6Z52sqY4kiPQegWXwl/KxJpOOp1G
aC0lsyNOPga3ta9dS44S0w4pCPBd1ZxhIXI8B9e+wLAFjfJuEFL5mhJmQBINdxfzJKqESjte24SN
AUKv01d/ZPbhChgO3D3psaTm2+JLjFMvZTnYbM3wX8pST/5KwQiSVEm+wIHe0kQ9Uv9EeZiPi2WO
5rARPlLMv1/4zeqRcHDG0EMJVAMo6Ak6J6gb5PSENb36JxAJrDr6uf0jk08rhCTn3eTeY0HrC+Dy
PEWHZEtaTgWaQ4X+bF13tttwmWn9yG0eT15JBH2e0DgDNvHP26QEpr3NJwJYCn6DFnakZe87XTxx
7YsbvwWRIUO2E99EZ6HxQAoBJ3RS1yT1RXYBnE4NcF2F0CMFsK0CgEuoVpjPzHKMSPZWZS7z34gm
T5La8VYxZzNxcN7aiYCyn3U4lpbJTK1if0g+T5fuXA/AjchS8MMmqT0tdRBNnisXqbTyL5hUnJuu
LYw2ckrasORabs4OMNt/WI77dXj0CM/F7d/nHxOpJp8SCGn+co12vHvTOJxDicYOux8YLgj+0NLG
ETUz6wzD1kIglmBC2Ldlm/xjL5TRLOXwjoYjSpPifyHKMIwKNu3X8xXLJnBkiotHaJMQIzMfUEhF
6t8FS5sf8UsLjMiGlhmpdVqKgxaRGOXF7WExPHPBmP3+4GG8nAnC6JoUTvXbZfLHr1Di7pxxUKDr
CkMV/kHRulI1L95hXdjxBBj8BONIR2QG0IazyWYlG6egtIkMUCzbOvynQLPAU/iYW3zTNiMysG1S
LWxCtMS7ZphAw2f+trsuVYWlPB/it1snKS2SDPJPJyUFrHaiqD7xAm0lV/EZCvpydLmsxJiYgvzg
n3Wje0K09viQ+n5VS2xnig68Uig7CUDDXbMjx8gzfHsXRurpAcZPPYMhnx0DMKV/8+89DlCv0EGx
TV/kvUNnieR9edlJcGMfW19d4WDmNG7ay31hMUOXehQiJNnsMoM3lBzGiYHnDc7hbjCyHia/A1QA
H2P2CCcOlV3xPi42/grbezXunGKo7xqB7QlPzCNaXQSEn+0CsBJFJDpDo9rCQXBDA4cF1KaniAcu
ffLos8+EzMa3thd3Xq9SlLYAvBHyJopbj/v1WQhqRBo9Zvj+cIj//BO4kOnRAFoygXQiCj1XQl2D
KDiM0A4CTO/kXscDVuO7B8gvEP2Bgt9pXCLAA+JVYv1t+psOoSV0PCHIxpiBz1zuFBP5foGgSIv7
NmQh683DpjS5fqqj84IKAHYsmtdicaEs8RJm+IGYlnqnllCf3p6ybvLoyY6NpmTPcxrSd/dFsiez
CwNcMkrsxEUMe8UiHywcF+XyPZV+WgUl3+NGitXYJj27MUFTf8Dy7St02ZK0cvSD9GrVpD4dLPv+
7axJptIo3sNpCtB+ePTzJ8UpsN5r6pRKHO3TcZS0p5it9j3PFuCi3QxiigOyjcQ7lnSS/7hpG5UP
B1eFT/6+2L5BTWwB8jPW9eRde80DT+5zBQ7kLAerb9DCc1+uHNZTI2rlNCEFZTH1NhLjR5lqExnT
MoSFmg6sXxEjSvkFHTzBXkwJ9s1MQ2PM7sBlqFaP74au8PWnvuc8BWmIo0T4NeqWTdyJUmn1k9hj
sLexKGYesl9K+hSPidUgyaYMZ95O2LaXEGeWC/vmXZIOoRs8uxWgs37j83EL5rsIGhgcjY2NeOT2
IK6mNHx2hOQc0lJzXzyQj4LuXwGDQmJQ0HdomZPzeNgOeUFrSXXrTHaqu7QmsvGml9Vb1nnwc0bg
akZdvsh6i7HiX3y5G2Edf+ejpfE5tb+IPuV415sQ5e+jcSe1u+EVgOSajXVpa7UDcnPrwAAQC2k8
knJLlWm8Wjx537p0KeRvfS9g462a0v4x6TaDWdhdOiFXwL1qD6nUztpdaY5jaQzbz/cOGGpFeX0k
FGYQC/RHGVObXbwQOu6/Swx+yzfNC5U3L7CFnPd/U8xcHE2TEEV8IGfupmd4Kj/YxWpjjHAcIshI
Ew4D41XaedLolrL/11/RMw9umAx8hUUcdNwO9yjY7+ugEwdOc7tKLlj47hC3s/fxgIovsOT4P/fS
+G3XcVGu2+L1x+y8KgjVVBMYYxLDEILKJot6ndkPHq8hpqIhkENalNnBaErGigLJkZSvJ0qeufwa
+/WIRC4a3wGDHmdR2NC+nKEks7UsDKw/2RRU8jy9+CpY4OOChr0MUPrJc3CglvS8TovDsyvw2sdu
quh8HpGtPQWFBh9RI65G97dsZCZuj20H+61TqJnoNDzm5e/Bc/2r1oi7tJCcLOLyrZHwz+bH1N7/
vUEq1SmoF+FZyEbUUr5Stltq76E/MXjOFVJcrWMKKAcK3Itp1D9022UlLQAmj1MmgRyNrilsFllF
c+0STS73AvijRdkdlJ+MkUHi6tBHC0L1qE8vS25Ewe0dDc+TS94+d4CKdH4H22BuIo/2Lr/b0VaB
x9Pne6a/nYcwsY5KyfBlH28zkIwkSKXIRnJhXf7dtSJ2y+br1/SoI/W/Y2kKT9AkaE2PBHWQNDVK
RIkfZ80zdv2CuJsGglRo+hxKy/vUmhfSDZdQVhNoaFJszWn+vo7SNj2dDwM634NQoqwIaxhYPgwQ
2g//HEyO6pKVn3/C+qUfSF2d4NfxRgWPExP6EAaH3hLYBcZsy+n1IbFacj3895Zdq1Rl9/rko+s+
7IF+Jvp6a1wu0lPtcmZROTbbYUD6dwJr+o8Pzqj+i0EIt6SIEe0KBYVd7G6i1CkLto5ca5PlvuGY
W8Tsi3okq0UImjez8svbZ9ZGMJ76OkC2uCc7RRZGceekpkKjgHCxn1VYuEbYc74aRf60PqUZEbsf
wtwcwMg+g++shPcI1H7Eq4dqKYQ/clgjjJ5h6U2IdpdFOR8voenaZ4o58o8OLEUuRd/7EU5C6TRA
YB8mShj9gE8SOz95sMyWdfpQ2om2fUgUgwY40FLUvHcgAVvLoFcucWLmDwMnQ8ifNPIXw+x/NkTN
8SRMPdvVzK4rZo1poYLtlgTKdrbhq8jeWEVwnPZ3MS52706n2b7jgYzhJCcYe8NN1t9a2VeO2GjJ
37EJjy2hgsIpKUuP+797viPJyTYd2VOIhO2PpBEEy5Plx5HSsYtzKkKVXIoyvZZ7hRLH5zI8Ckms
wo3lhnQ41soXqfi7ib7epzJO1vDwD12Ax0KdXdK52NhoSkO+K7WIjlLmLvK9JVV20uxOPU9Qzk9h
JUBgtb9L1YTkC1t2UNOIsTw7LE0+cH5vzJhwf7lmToYczVleRLLtptLX/HUp5gqPrOYPrhITCB/2
yxuH5qYUsQJMRiR2tal15Kz2U2WkmoBM9miZ4s1hxoHhBTkSgBBgcSXuJLIoCF15o+Ki/nnJzZfC
+/HtYDRlrI2NZNJNxISJppqXN4jgcQZqmKhvufQ0SmAcuTNUk5PRLxnoyK/i5+N0QbFI5FND1joH
C/2B7dtcTdrm9fJmGTnEYCOzKGFgT1KysSd4alrR2iMOYMwnT03E4+lwfVfIvUzZ/nbhacO8POea
VLYETCCWnajvIxUZi0ms5CV95Ebsct2wyzTIrOrtlok0hW5m9WYINe01DNiwH8Qpas8zm48qQThc
NYhYrI8JrO500hK2VQ8iz4B2hr30SMyKZGer+tcabhCcMV/MqoDdDtmVsKEIjXqu27o9Ddo/nZYp
z3/jR4uZZFcCE6Px/V1j79va3FTaZcPRyHWszKDChcML+DDzEHUCMXTsfZm9B6GPjQ43xb92BZeD
c2/Q2qhHUBlZTSqsOlDlMBzTxV7iUargQQHA84G1ILfrt7/90wzFCOITKJKHE2w0SePh9MRS3aTl
XsZA4e6Z/PuOguC5BJtMwncl1UsLkW5mlu9fwiP9qA5ot17gsjf8GXS+Mm5r+EFGFmSmpkWDtFPz
EEYaqyFlyGnnASooEOlPqX8H3acT5Jt3i5uPKKlj76SBveJR3xSZPVycEOrRr308CkZuv5ipxxuT
mXDuUCITwXn64tJI0JmUYVxHdO5gXHymBB8t4tNuXyyCRX7Rcv9x9ycjxMSm3H1dK6UGhd2+ZjO8
alPlLWlzAbUl1oYScQM0a8LDz7HuwYCtPXVcT7ygzgzpJVo140bofcuzekEWA0C//NZrRTCkUVjB
beVRwNy7MzaHhI19T0Hp/3GhKI+ziM/ZDhhr8DAgSbp2F3aQY640PeoLKjOQqulBHLmVrK2SlLM1
RNXSesQNh66JUqyIr6xtKMpKmO3F4Dz584cIf37TIcPkdwPXBMjOP6A1soCpKPkn6IW1OQjuOawM
skHzQX61aHQvyvjhsF2oA4dXYRXe6s7b5eRQB2ZNCPAAzG2ye2lVWj9bvFCxvaYm4DckfP8wLxJc
+msLSusdoEydAHx0n3bVESOsU9x9qvyxGZ39u4fshk0f3rq9Us8B2bCy62W73u2c0L2QSW7CDdUM
W21DgN536z9chMCyC7LZeZfL99dASmABU8ubZx+uokGYCHkUCJjzcs4igI5s4zkqYT2hCy6GNp91
QEAZzewE4+0MXLNUKoxDjvVY5ZtCbk2UUacoWccwzZTYR3+Ld4ZlIzAGnMmlHhf6onZMIbVeDrTV
OsNHERhqDAviqLHkzADSsAzeokba0Ik75249IaNch8pqLgxKSWlIZqZSc6SrXbOmwAcAwvYcA+AC
5PB5kcr3d4kipKPkhpcPHwMVPzOw8NlWghl8NKFkpJKGNtNRcUG8oDIlfAo66xZc2ena2o7h8pAn
6ScghKuAtKr1Kg/gy6f/FaPugRyJgdPrLrWKHme/tOCm6spT/OHHqG5sOk/7egkzIb5S/VNqpof3
4HhuV6NLH024OlHi5Ewqw5QIGkatzENN3IUiwroo3TBqGl8YzOvEjCG6ExrKQ+iUIQB93h3yrcEq
1uEJid6wkz3N6q5nYCl9FPrzYTqkL6GZ4//dJlIguGTTFe4Lw7xNWL8MQL2M9IEsKAjj5jx8YdE1
QvFgHczRyBXJ87t609zMLUa1y05bIJNhDNhzzHnCMQT0YOOUZLNUcaqUKgVNybZtVGMJjYx1S89I
ck2/a9ZRYpSlXbSDuG91RiIzryzWBy3v7LtLB9xr5rMExuwhAUnh3d8duZBG7cxRLtIJDTtZhHTH
YJDu1saQPfS1lB/obVhtcScQYrs0IbOtF6TSQ1sWYPIQvvFcy+S1m1UIFvGZumkEADpGaedI0Uc3
5HgIVLpu9h4U20D7bf/Gv4G1l06pQsU7NlcRlXClY9y/39dinGN25TwwklH7m0tUVBVSfqRmReUe
JtDyPxFrJ4IDSxgDQEFNqvj6LEUjQog6Xx34zPdKLe7MvSiG8IYrCporGM0JHD4RKQINdk2lz8ce
nGFlIQkdbz8yagaqZgfxyaPyKu6wXN3Qz08g86rn41VZyz5ykcKMnp1GSKqNcisgoCqQgUsfaXtl
SKJloLkfMdJGcPmrG7dSbTTrxeTYkEXRw4LKQhaxmA5Br2A6iDYREm5eJQUTA6xUDeI6dNTSasgx
tprl+JER4Eq+ZQ9ImFUDV/yv3qicxIEHSU/wpJ5/bK9pBirQ6FlTOnJL/WS8l+FNw3rxXFEHsKmR
xVXggE9lcpW7UTfR7wPiMkj7umCpmLsj9HpEMkovkJ+crd072KGZgWcQbqxLWRmIfb/IORNHTZsw
WWzKxJ1TDjgc8xywUd783c51PDHGoCBA47mx25rLI3DiFcxnB1FCDEL8Ro6miYusuhkOg/ivCfm4
G8zrq0mo/r/C5EBRWjzZ4qb6PavoXpCsti3YbftT2zZE+KBcZ0c+tGo6r0Ulk6MeBkVP4LgvO7mT
zIJjhVhlXXx1/rw/7NTU/15v4uxAzV0R3rUg9nHbXV+i5yH467jEGA2XPbv/WDHWUaGq1eflGv7Q
3zAl0YwckfkLE+7PU6gHewoO6sjOveQuig+9zx+Q+cBM2RmgIp9I0mVrlZB1YbARd7qPn0Tm/h5D
zoH2hlMwHwvo3/srxxGQWrGIRgYrjfTHUlc43+PgD3hic9TPeA9TwudFwVSn+87ygq7CJUFKJM+6
uD6yS6Lyjey7rtbngTnTW0tyMqBwOaxTDYiMdVOKBbCGhns4NuwY7Bmav2E+a0JwF0RXeRoRHfBF
9lH1zTnGCNLTeTgWsfHzsaXrpmy5ST3G39jDecbf+EVSyLJ9tNdoE6Tj75rk0L0YROohdmaPpz48
Ox7yLfvAwx8VEWONtJKjuUDDHPapp9RKLirTJRvbv5aM0yQCbOKqPC5RIoUIUn3FaZ3bFpcmvIrE
X3R4aL/QkselYHYC2eIytWQLKEWUgZjBw6VDiHmHGLEbkpjhVlKBDXx+dAGQi3sKg5HU5LPIQL63
tIfu1XAniNipjCA+L9+SdT90286vbe3GaUXG9bF8XocCSSJdBGVpfojyniNGuTZxwrf/Kc1cNSv8
4mzIXp9Bsn/4T6zyDDCTnv+q/XD+1BsfYr8iG+eQxsQnT8PeunahpFC0vSGjvji7fOoAfYDLqAn3
xRXQkAxHJL/PAl1R8P8tbSjJzQl3YzK2j6GLosJ1iVmEU2SvVsmTuEKpAiZyhghBuzl+LuAIvqe9
3c3L1fYit6oDEmzYu/NEDzuo0W3ODJRWz+DOrtCDRBs4NALZHuJt3SWisVuyHzPxWmIrB7eo4oYb
Za9Y2ERJBfsD3mbuEkXRDYzS5mACbgXkMhx31V6EZ/Y7bd3i1pj93iBP0cTBCAm2lB482m5Lfipg
3PSqc+arqjkZv/J1o+d3fScTUUxNl1N57U9DurzEsfU0YlYOU7k/5TU5KBEopPVmVjFbjNWieUeY
ozFNP5hbmb5xWPicQbeLmUfoNCeDVteDLaWhM61CSWam9cIykDDoVLIxprKyJ3PhOgHFQHPn/T8k
zQf1Pn4o/clitpkxLNW5IBLByua7ss7c0MAhQ19Y+jzKiUcmR2wbNlNIAya3oHCPuAFha5MKkNO3
6mCSG+0RKzhB0vJSpdNxMSFh1TDkO0vyAXcWA5jokBTdwyZ7Yfp7tjjfi1z16CyyMy8Ynt5qRGAf
W4m2ihCXfo2LAeFtldE0hVUE5M+0pDL0l8emU5wldwdzOj+9jsbjF6gSh/cBRzWi0LkHmtv6jg2+
DqVu+cbUnF/ZivYWyB9RKUVlxh8eSBO2QCFJC9ER2yLV4Wlh6OVDWWLyuPv4EayRjMy0BumdhzLe
eP/izBtQaDywKxklW+Bgz+ctkX8QlOwFIm7FWm1ulkoT9ZAuvCVz120ffiHJz4jp/lcFeV9rtyPP
4cDwoEHTFeKltO3vk0mozXxwk8CSDYVsNqYPcjVI3nnb/ZGjapY1vdlRfHPudLca4WJZmxoAcaoi
+mmdqvGuJvF+9UEmPB2JqBJZbsckZ4wOd7cjjT7XSa2MzVFEQRTos1X0ZQhGMpGaiaf0jdWNDfKe
sbSYtWYl/fYJb/1JcHcLcPiPRrGIW6hWdWvMeGRLvgs3ckkuqmBTqRGH5BTgIvCbjivdfBA3mget
DHf0miDI+Ir33stCr9CB1HrI22sJrtYRqQKsjUk66Bqu+t1dHOlUz7PfyOyQsLvDfVcMPbpgHhyT
jCp7/qppPe4TO7/CNrl/OGPr6lTwEvO29pb/0ihn4YFOJzDYa5aUtFEOT86PhQcxY4UVrzmCvWbW
xVpJ49gh3yTq3ef+/FQhHQbBwFaZMhGkfP1QYq7wALXE2sgYOU+dfR9XVXcE7ZDB2jPoCZPoclX6
uZzXG0IFbSN9Z6z2jTxaKBwlF4YMT1DZgrLt78T6x3v9TakcNiNVhooQAzxi+k5Pl2kgzlkuXXYe
gC+ppOl92b7Rwjti5XkIGOXJ68roZp+B9/GxH5P8gKVQXReiL0AjbxaBB0rMipjZTPH1jxWJBm9n
/MJmWnormncjZrpRu7k9hPKsGHYJDsPMJDnfkREQPUXoI54p6E3DomUicjbzCMWd3ZYbnxclCl1k
GlCN/aJw6UqSqBWcVEip+ITpfGIF3v7m+MaRagh0tx5hfqy29n5ERAiGB+By9Dcb70cTs+eX5xz/
v0vlhaX11t4qQoVCdqjboe2i89p1TrPGaxboSok02BFhNXgy/Swz/yvgCDg6KFbYi9GYcBLv0c7h
DSLbv63tMMcmoRAATEdbRmlitAVTSlenCYpLohoREOkGev9MsYRaz86vIeY09tQjqREEIAPyVurP
NUtvjNLrhJuSEEAp5d9xrYgV9MKBBFoGdKWsNyBMvXEkXqEECiNhnGB69iUpe0/NTGAYHnMF2hnu
mDidQpxT0hXf13adZiBrhsvVgtHbVLPfFM8BjB77a5ctM/pP1SuszR7eZlNio0gt48aLC8OWFdiM
fS18d0TuynfBCD8/fnVOYAIczP0flFx6qHJOggrgV+CwJZ0lCMp/H5JnjBmjy3S8GRMGtuY/yNY3
n7iKzOBCEZ4h55nscckqRUZOkqat72QMnMNGBo/I0D1egfkZOgqv1hgFGCAYa3nEKVcoiVqKCJ8u
wuANkMC6w+YZRFc1xZJnuwlP2jQGCj8ATxOopob6FuQFZPGyxff+NejEg+HnGB8safukWPUQSAwj
bBFE9hLTvtZNtUai7Z59feyeOXRiWBPwkcJLzHPiWqgEkzBbsbUYTTxS5t5nuE0+AjMsx7nX9JjI
7nITdmnA+JNhjyfLXVkPUF3EOETv7iDmaTLnXsMFCah8100PexdY1baT5tES4yhNqweyhq0UHoay
9wOAEF9fKjj7ZdggJo90C111cdBYoi/uGVSXcSiVPhhlPE5o57anVr0WQGb1Zfoz1ybtbjNTD67c
yO9iTaTT5nsRNVsNtlhTK0pLI+OF9+sU/tleFGatDYuti7rblkv5Vut1M4zRnrDxO5Ni99Eg8JJo
CE52GMHhnhNe4pBETjYPrydKPCpwjmcPhn1E54wkFYaDfjDZLxONaN6o4JILWIKwXVS1bWPeFK4J
zBznyZZDgwX+pmaxIl5Ga4xO3Znm2UIPnwlwFcXZ7wGjR8b/CU9/tOCHcTRhD/KuRYupRy9JhWI/
GS23rXwNWpatlGK1+yvtAgPTzZf/2rJQNcLMdokntZ5P3XtbPsMTNEiIEfr8k5vlI6vrRajcVsJ6
DDQzFFaB+A6iGYL0jyvxg6brj1pik/ZKngAym8xZSfJhS0aduhFiHmINYJjJJel9VN23RWT/iMyM
YHw22/EaKRe8LbwB/W5nTvWycl3ZnFeBO+KQPVZHuPrCRpJH/ZRPn0b8+lKPHUxKPN6VkngqfxRI
9ONIMs/FNt+WynC61GJfHEXaI6tJWdo/DOBt+EaVbeYI/whdiH3WGixfBtddBDkK8Rq2ml29OJOg
SRP86cr2O9ILdhg/xR8ZVknp5nEyrLcAONNMbYX9O8H9ZoWb1COeCDT1tSklfWbGIqw0UUv6GGz3
J73iIxxtvQmCk8wn0tQhBI6n8nCf3a+ZbWgVFb+KouWQMs7dMfY6jJ3S/CAANLkKqbk6PQfcIjwN
rzuH/x9SGHmPj2imaQglCjoN1Kf/j1var/DiyRdM2ojxNow9c6BclbA8OL0suoQi3NgfTcQi3NpQ
EFnyp5MK0FFxUztf/hQBsiAnBPbIlMS+UAghKB8eNl+5lgkaV6iPS2Tm+8eqZm8iGTTXJ4AOeubB
bFbBY3g/Nd8uIjJN3PciP392FSH3UnKoUgdzICev5Xqbr65mSij0bUKrea5slbt+rN+Ipnz6QQ1e
ldmWJado/T3dOnYBvFwPih4fImIzMT186sUQQm6aSMtCvuN4WnQPTa8tfwRlxp2D3XEbCZ67yowt
wb8hlYh7SVgOOpPE+NqcSkBJv9Ybg0A4BizwcQ55QgXIlM9GTfHfkkqTUYnrcp+FFgScFHN7zwKb
5ATvn1dj81yDYgNgBZmVmfzHkHIrMIVsMdxoc0odfOYU+JcpOAPcKlaAubKvhFI4B7ei4sY2fxms
urqHyqeUCFGrGJHj2y3o2Mjy9L/P8fUJXkQJ9t7uiSbQwNJOYRh0wsQAm63b8p08iyLvV8452NXs
r6opNCMcoUiX3LB/cn0Wu5I6JyNF3ZRFI6XF/DV6GF8N3t5DDdcOMeXvfhV747qRUbKqvZKk2ycF
Wt5Jb1m2bg0FLbfech0lhg3WInAFWeYvAAFSJBtKhNPid2ZVRmTHBfNtaZ6YplPhwH5WcH9cJDLB
5qWFQdLPzoB+dVUxN3z1cTDNrR16gafgk66OkEvaSwAcZK5pTRq4fpuWnxWSj/bnxTpGM4PHqUa3
bFVPKK+fPBK3AwhBskyKpaLEkbY4KI/poRTyoE8ULy5RLglwyu1wMoKmg63lyrjRVb2aWAAm8JhV
Ks9tfYMOe7FHF37+JYWwt23Asf0IQqvNI5Vf1ccJqdUDWl6aS9F17/r+BO9/M72M/a7GUHk7Dzdt
vex/pN8qi+giMi0dUd3ZTKPs9Hj6VafD8L6BN1gtNL8mktTu/KMXGGY3qOIwBFoCYdcOqqH44SEB
7gEgSk3u/2cY0z8Fr6kaNaFbusJ5ZUSMpS1/p88ZUsgNVstF9n1RQXw3CR1Mkrv33Io3rjUTgnD3
mNp+FbP+l4X3Xg6p5nieRv4GQ4zdXrrQ8TsII5moHb+Elwoff5rgO8/5nB/Klv65bd8VBDmj8UvZ
MC8KSajg4q5yB6k0M59HduKZ5kVGMv/vdhlTY7X6Kz0tZobhKEietZJy3ahCpFGDqm1ZaNOS9X3M
pT+Lh8YoUHyfTv9BXk+vVQr2re501GwO1CCpdgdJnAc7LUaUWfKlUSipLdpAc0/Wh6TyjN6MjCWo
RamA413UT+YfyfZBf7z+FqGtxy9hVxSXRtbrqXGABOSpXpCsGAXpX7W3JSfrmMWUBUQ3z99W9Fxo
s7nEJS4CX2jWl6DmX+eiLu6UqSqlTVsAVckbHNaD8iz/lPxFFobvPXCxH6nILASWjdS3gzomjVAM
WFCejkywViEpcV1JekPyIYRG09poRCgSlKy+QCBatcDOyZckNnZ2MxHySXap4ilXVgWbuSMAPlSU
fS6aFKJ+tnC+E48KCbhBAIWdjc91WL5QBwaMkA29t3/vwX2TVD86Dq31nELWUk+3pJRhAolDfz2F
fGbTU18BWU1je9W3a7eQUgsht3pjutZZ7F3BVqQl7FSB0xYgVT/Eldgf5X8HbikIRxCBRnzt6SPF
/SWQVPget10Vh5pvsrQTyj4x0bdprXUQ5USi2x9W2EMZKC8Ji/GXj17xFqcdV/IeDaK3dpPurz8r
Uec/AzSpO9gf6jZti5HkB1IcU7uOvGk+hWy5ZitQ7Hgaetywk4+lCPxrPNuXL/wpCnAE/eZbQ6SM
Y963vLvU+t89JRs4S9XAgUW4HgCJvMnezz7BEOCHHVZEuo4U4yNFU6vCn1/n+BzGjMt7u4sZIMb8
L08/tEuGe1u5Zjpk8D6rkmGrLbWNcgtZ7zBtSKSZfftwqEzBizdsbeZr9sakiaWg3jdUXp+qVW7b
aesFaEB4guz77MbbIyScszDDtk8iwZ0TAZQuC2jrcln2UVoMdRvLXZrfA1YbxIskEcXEGS109iAe
SPEC3aIVnj891xIEOLA3cgKPqxHEiYMHL8z+4jLK75Zd6DgQsICOvlmmbWS5i54V5JPqK3Gfs67w
Vx/NTIEdk+ua9NfOm2QB/HSztT06v2IB9LjSIRuu+ml9hpig+Csrt0NUVEFQjOAJqRIBJJQqozqt
YQ8OkCbwFKJ/2X/xMCTv0RSws+awr94qdm0zF8E8zGv/jGmuTqIfRPpAI2PPpff7uYMW5+xueZFR
7sMlSxJ3b1CRLaxZicw8sbiFj9YQkhvR9QfQrAkRmIsROjVW00bbtDy88AWari6ZmRAVRVZNdtwg
A370h86O/rEHtCsdSwhUJtPF7ZL5tTcKO9brq/AhhuaTk2txdDxkZ17UuAztW4H0TjbTIlYD90bM
2W8LAlbMiDgcm9l/I1mjKMcN8KcjEeBInbyIlg7doCiN9viSSgE13yzsbr6plKmV+10DfGMA5oaA
2KjqmN6Yasw/7n2BwoOJC6AvJJ43OkahJUC3kMkKTkKJR27MqB+BxrlnXmr5JsH9VkIHLezHY5Az
hPlyMP6RhuQTY69vYK7tda0X3nLpFxz0W6xVNNY5Nq4XdK04qhmbdXMrzejbSr5XsBcPJe8+bgqB
CWY65YP40YnySzX/lfOVDK8zhfc0vkUBN8bvp46wVDmkK21nfzgobxCLjGQU0mHo9Q+OraBz8Tm4
68wNg2hX3p/M9k+ecy2HDmHGkvcPPvg0fnS6t4/rDzRL7DvxVhmNYMGoGV+t2h1ID1JQZYdtT+Lb
MTkyJj4hjMOj3vxAz+XPFwD+Knh0DlEf14HHzNgvzko7hD1VbILnd6ucVmZUJKyuq5zOliCSU6v8
5J6Hw7TR/dX8e2+jbT61GZvF7gCOK34xn5ZoD7ZmP8KqAtVS8/Ey62htS1siJV4ihZfFhJzXFR17
H3ylVfHmOGFCx0g3f4Ov9tkPRlbhpj03tvyZNI/pvDJn7Un1TqbQriBr7cl8hSFLshY/BxjVyV6B
qznVRC6GH4xijsXs9LRTtcSir9iYwB79GvVG1ynkxledE5rJfvYe8sLD2QIopHW3P2u68uQbgOwr
Mry2BRCr0Hdh83eh98Hc72liHAdax5r8D4M5J6gvebi7QtaPfFWkRLBbSdwlRVBPjk329HKfrVr5
U2M+ssmHeOVDn8RX7bP+5dyWbOdLHk8Hi0SrAywdvfvTaOuVC8H6NTsrSNX8EumzsDiXepwtSWJw
5QX2pLLGpJjOMfE+rx1pk8em5v2eIXXHuW/em4+Kd3oHXeuI/cxQ7nweAbppi2Cx77lAeHk665Vq
FNzl9f4hCAWvqFz+CrUXgqDCW7MMEAevKQKb+/LKpMyOqsP7NPocadHx9bLg4ehF8J0O6hk/sVDL
GmAt5/hVgBkdiepDIHinCfueFejFQ/JDJknAARV632tCfvubYOBO5QQQHiGfYcgbp9N3G84sjc7A
Ukki88ai7OaThAJdG3obGduSvMaN//xlcwS+qikgA8mTm8It3EA1Bvymo+30PDQU87Vl5ZZUhhM7
4psaF+dtgoInpqkY2U8kmqMPWeCR3JSMZQuNV1aNhrXaYAbZC7VDb+VSABzpsIgCcqZXIhakMpnM
5H79NEtIRdivQJ+7zfXFXzLMtrg3YKE9S3Sbl7xci3/IpNX5KPUuum+FPzrZTFtdC8ITPcRYH8ok
Th3Qm8CFqH4ysciNhWKuvv5RUxbBVH8uB118NIArffTz3d04VyCtub5GD0Q1QPl5ZwXKLm1D7zDx
+bSqcXtu24ivemO7aU5Wnq7krvpwz5vYGkC3q7eil+RFu7XGzM5Q+UkbZ4LTysuOdQvrLEaErEE1
4nClAfmoJS8/tG2qXdWZGranmHZI8CYV35fCJyuR5r4yIBi3CnXxv5xqBtKKUFgYOPt1BS5UrZxm
UUd0x3u4cENPiB292WnhRGgEAhCSCNtwZ4vaAgzpGSyBz6kZSgyF0IVvp5a+zYPhd7Ul+QqgCumq
T8dLKi3FypnFW6axUah43uw2A4zRFvY1kQ9WleWnXHgq7B10q9GbdjKqH4VUBOETxafsRW2yTUYg
86mwaNjPfMJPVYQXWupMq/PfRkPkQk7S3xzTjcd4h3SvSPf+v7SyWOUxBVJ3u02LSIqAAMx+u/It
1gQ4od9uD8ZQfRLITTHM+/KHrnLn4gVAP2IUyAaNfBzZAPbuxJu+y3kmpDujgpjiHJUTVVNwagfu
f0CKGqdPa5GMnK7fQPPnJLK2KIa68qe239UP+QmO3afsVU58LoBVIrA8MHRdTpQ9ecl3cRekJcVM
t+nAnoJ9AO/j+Mkmzr5Vjyg0h2x9PpNSlamg72dsmWtbLgNh63DdGSeFOew9MNLjMMaCQses5+4T
BfUko0g85HfEm99bvzceof89MUKPvBOz8F3T/DyTbJ9wzPJ5hVdRwdQj5sHz0TCQW1aJ/uWYDptN
T3BSFXpy/Y4SVI2p1fCMi8sVDovYfBquN6lwF+CNzjRZnhHbuH1KK8vsiHzBof6MvDGnvHbMV32T
fISMI2AJ9nZd5qFeflboo0rieTDQc7RZoUCOuD9ptwcVf0WNQ+j0CLY2krLWWZKfFUk4a9D8W748
RZ32oOG180nR607TmB694775GjUpvCqr1FlBE9EXaD2wRWBH6KdKfVlgdYMwlMURbRbQvvd27d7i
eKQHGtQZ51jBxYH3CaP10LATXxKqzrNcC8kqOCICJC9fkUFAmajtNhGdKnNun3jgPV9F0YPkdNDE
LmPHhst9uuJObp7M2VB4TqfIjs01Zki4Z9MuAY3npMU7Yk/+5i8v6naJLP1Osze/3P2AA7UQ/5Oj
kNHzoVMbDrlChM5UzZzT4aOtXuQo6hsVP3YaAnKTULoBjVxkIytlJmhFle5UL4HtpJQzArO/0TGD
AY76A4ahT2CoH5N5/ycSFKj61rV0cItSuOLnrrbovU6986TeSsJSTkiEaDaAnK4NP8XRzPUOXuf1
b29W6v8KmKcrRIaKGsmtmw5ndMOCItoS8/95NkaQLmHlLVXXbuckauPXakE2vJe1kpOBtf8TcXS2
79ptzp/IEVn2EkyfNh5zHmFOriR6HotxRt2ODh7k2kk9clr9CmXDVZJV6RVxT/Dq5HpAwnw2n8eD
6s4Mlux4Q3KEES9ZHeLu82OOBhpKUsfgW/X54xbJShD8pWonDl7LG67whTClZDsYHo1/63Hnna0V
O9VK8o6qBmidTQEUNnklsuVmMW+wFyGiOGdt3FOCYiQ1a/jWviXPV++rkNF2y5NvDacgG6b2Aru9
dlr59OQjXtdhdrWwIzvAhdolvutsbtoLuAuXgpvvANStik8TXJCElvIENku3QcRKpUHOJL3wXRwX
zsWqu6z3tv+0/SXfGn7NHvCTlrl2C1Z7PudvgSe7b6oz6C/I7J9bFuR4Rlow86fS6giligpv+aIU
VVEMQciQHv4f2uTSMAahsjjxHneRFCHr/2znwKm5hDhx41gjSHNgioldJC1biuqnOXfHvqgIKjpk
al6+Uhj0m1EQtYHmqIpMF1eBmkpU+5xaK6OS43FD4hLoGIzqQb/VxtZlohk5M1KqjbMbuOgx5zB8
nduTLHakorrPsC6koKSFCMU13dmUwiAbSAwxsgZTX3oiiGAA3mPQ7sqxyV8OsK/GFpLYkAgtpFIt
96NKQBu6N5y/mZuhegbukSp1yPI96FPaujjipi9dHukHn7R3B0RTDZb6JavY7W7yXdPKSvzz3h7J
mngqJttEKlV/GalhybnljT8JEYV/W00PHokrvY44mfq2Bq2cTPHzJdZc5VRQ7KW+AQz733DIXou4
mMUk4v0okmwJYzectFCb4kEsWUDaxC6tUQL1VAU5JQoMfAPfD9U/ydhq6/H8Tf4/CgghWrshmi4G
Ay8zFDYKtDtJgJVMmQfGqJHcO1/cdv0TtuKE0LmAuRQv//+VVsb/OowOjrbJ7JbEFWvRLlfS3OIv
FQkfNz8trkpzGlnEtFuzh8Yv2uGVv7x6OLRyXRWQN78h921d6vVtArqCA4X3v/ODZonOjG67dohf
GcLrqdvWzGo4dtj4CgWiMOySwMZfT8iOOXQVECHwGwfHhUZ8HCJfnmdAfkSoAVYzxrKwF6d0XSKv
kgyiNPifrPemDORAzvIDes/y4KyZpeaW756LWa0TDTVV9W4OsXt81hafbhx6JAyQiYCLTAK21Ufe
OJou89ME68sQVkKnsgDz2HEKRR1UIW6qa0wzYQ+l5kbLCqp5FoUg3s0lCPXmKkF96vQZbG7sQmcw
iOG1QD+dRBXzn7xqyXy/RZaXsHjSdNd0Ok6VuFb2ovafwM5UoCT8/qUpUpj3N87xPuDTz4NWTJvq
ueXIZmFIN/Tz6Fj3j3ZcFuvwLqbiNvztMME3WHZwyTmKlOAiJJDpIV8t8UsVeVi9wy9LAnVh8XiJ
qqX1j6KluKYWtRuw11V2LH44A01pGT50Yp9hmTnzSqk9WoQCW8Wz3iXSDuqvr/WBxo3IJuU0IWIF
tZW/i3le5VStal1T+zx/ZX2AZqFvY7fHcDVt3TjWpd+OdHkbPquc1Y59aboORFkwcUgHunO0LRx6
SitUQa93XsiNJLqspYTaRUE+QPYokcniJogHn5Dlf2xstp/G7h4qMkSzGYqT9eiUL92DZFTbZRz6
31ZCsu46nEMtS+FefR0PC0ZFUnSLgS+sfi/LBziic684rBKmKSdBHK3IC2BubWiywxH3A4UTMGmq
SRUW4XcPjjC+4fWgOKgIvArdCFphTqMqPri/nkmVULscFcmERhhrotbsFKOIOgGfbNAmUB/IQo9O
Cgyy4nqVU2fU7bQ6tqe5xnQFd7mnYTSjfxO/v37HfkfHtg5y1T3SrJJf5xPyWWR5SFRuSTpsfkte
cxaOyZ2qF+XgZNoiRBvgVP9QSt/tPuwt9gPsb9TQhJZnxzXyUyQkD/PNQjhFc/7MdDvMNd6XrPKD
b4VjiCaRvRBg1ElelQ/LSKNEUNduhAVly8YJy+RI2AyRmlXzbS3lj38jJOum2+S/fDsdgCa/Ryb5
sM9n3IvTJ153tpDOaTA6MwPjM/o4dpUIRGAh20mU8v79orr6rvMQxct12yuWMj6VB+4lgxtnZ+8y
jlH47xiAP5/PxV7xC21ic5tl7U0JjBG96gidUEJ6TlexGPHVZVX4KITqQ+0pb53avWotGWoTEodc
yRbsew5qyb/QP7jYijI4CFCzbNLAGM8DP+6UZGC5cMtWD1I5NH2cCtJAJt3jM4zswwtwq7MAmgOO
uQb+WNOZuMz8bmGOW7VsMOtkQtkjQkVx2kn/hvyeepZSBYqS4IFYxS5/YAxTz6PVjAfugbFhVuA1
I33zERj9BOPf4UsIuQ+yvm4kZfaHQM3rdi37fY2eWTzbHFpqEmZJWPtcaM+oQnwsBXNHpVHvm2PT
x6PR6yquwjsEA6g5TnVPE3pAFeHalgnwRe02fyBuRpDbbrcTJ5Pe9qYhShAOVym1ZY+DDmSZ//6j
M3XpH5wHV3VWkI0k/ggU0F/y3nhBJipK9JvGYXys3RsmzWAXH9NTKKpCdHwqHYY+cxSAlQ9lY+o4
8TDkS+BDR6jAX7oH3OUGd1piNybMHz8M1k0fssuwgnhzIghpoOqztFXwOuKnBNOW77oGoCQELipb
o6PFOUjtLFQ5/GthhTFnFI2LalqHtHMQ10D1b6KcH2aj/hPqOZNv5cN7D7gqj+AYDJFjrmMEqt0B
5Q86ND6I42b/n753jJQ3v2z/TS8jyJ7oT0SCYAQFqZxlNUdW9+8VI18tzkkehNGSyBdee3RFAIhu
PqyS/dlAedyoWs7G72nWqAvPnGdIQROC7/iKorNp3mUjocmPxOl99WyOgwzAty170BFvQTUR7wom
LfwDwX7kWAVFaXBE8nMr6lvhdkkhEQhm76vFYe/knGzLWGzWNQOjqe55yl529wN10fMAsQmjNLxx
hJ3j7IDnxSxPuA8HeBi5saQfYpww66oZjz85VxgIobtfACS+PCP0ROd4HfRYA+XYEb0xnbRLny5B
jvOAxxOpAxZY40QNT3hW5RPX4u++RPyXTbfXo+4yggT8ZUxG9pl/tTJrKJpdWsqEFHtyqBlmoHO6
k8IOCwDZ1AkDY95DpsQ6DYXxduFfmk8c4+QOcuWQMyu5NKFsqEvGW+v7qX/+6BW2Uo1lg8BcKbgE
XpU+7PDyEWBUPOxoFZOFnMEWYEpqh9FWejrF7Pwg3RxGDUvtRYb3fWhlDiw4wWkK5gRdYqgAQusj
XucFqMQJ70yJeKvCOTnogbFZw5igB3fepMhu1zJpqKvwkei266H7TLWYs82NtUgXF5MAvMh43hKe
Qjalca1vYovtOATKZlXdncVR1jgRQc0fT5F4ln5AUM69Dw0B3TCWZFSN02vNxQAI3wAp8M4J+3XC
z36JsEW3OzneLyHB47sCbUOxiWzJWJyLswxzyUuu5dSAr6n8nybzxE5QnpwNIWdeBBgjEaP+ggqp
7aYse+nPfamTu+LeaFSz0JdqJ7N2QvLMyjfBWXb+q4RYa8+jGkwbqAjh57+5Z6vepi/SD5rx8kVO
Cra6fUUTZLB6N7c0fCNy736rewItopz9nlnkOkF3Vnlzbff/OVrwCLwFYvAaFqGAW1N9hiinie64
cblziN4O1PC9qaRn6gEcMhWViIIqPXSrDdTIqho7oSxBo4iQozml8+0zjbyg7b9ZDWS2wSSiRNF8
gzsBHfcRUG0mo0LOiepLmC2kxwZUn1J9CujnQHM4PAEdwZWBST8n4c4plSTB3GXXGRK4ADf4Uv+v
yxOIGl7tv+t1xOdHOWbTuTMhV1H6+xe47ciptB06GDevQHYJJA3mSQ2lSpJNvtpT1JRg/EsLluAP
3utehg6HCvgVQrqQ2Xjz26zwD2ZVjqsg/CjIR7hTsaDtKbAobtYKm7CNCNV5VFw/WOf0xS5t5dbP
bl7kAW08Xv2L8Pyla72G9JCoCAwmX1hrG85//YfJCtMksFq2jlxnE6J3/5UMoZDS4gVgcEz38D/Z
6xRvMWj2t5gqQVEhhV/8ISEMMjT3gq2InJ2kwSiERToIXH46/KQ2rPXp5CgCOxEF2YAIlcT6hjXX
2tIsipnYvRWUmddMwZlAnZVjclGVbmrZRd948Z8MqINc/NPAtWSmPozkar2mqqYwEzYBZg67Ir1h
YfoGYT+sR4gVbMqR9fNoTmATg4MQdvdiItPGi1PUuyB7nVdThL2rWXUDwY7cCl/R4a4EqASl9daq
hd334AZDVEiuAEfarJmqn26V/hZVd1qk7wFP9TcKSlLmGfHBGctjOwncvSJQBQlvfzsn5JP9JDaR
tkOfZSOeums6mEikhVKYILaBwaLQlfx3vch4XnOZZiR19a2IzEbpOatj+nzh5ttEFyIBJWd8MLuR
Ntzxp13rrljSr2aRL2KpMPwPZB1HRy1SOsS8ktJr8yDcsPrsXkETgfPguA6qqvAyyElyt+NOcA4u
l9BsrOcLlvCBbye+y2p0BSm74bleEJcQMwmQ60J/pn3kYhhwqhgggcG3n/f5YO7CfX8OG9BR3533
7nBQD/GF1VjAtbGq3iz/2O6oOOAwqbOXg2r9TMjmHU9JOUfDGbG0/uKW1QkZ7pfg97syl4VAV3yS
MhsQZffoLa4SSA3NCnAUjIrs15nIzYdZkWpW0olBTTZvKDETnUU+Zlb8ubNUTjapb7S0ehs+cZBA
yzLGi+Ke05ZTGZFHaJRv70TVcn+y2/cG/jVYdTnHMskpbOPuynTUvoVaOeBoehnoZjd+Z/iknF0f
N6yar7kopIijcFIZHc31MkvKazJHw9E3bq5ETNx+/VWKe3tezowMKzFyFe3XjRJS1fOjsAY9hZru
emWxDfaiRfidnP4SdpOqWEiPfRqXzLr4w0fkBOJBatr+ONt6+QBYHG4sKcAOvzDX1CSdtu1+nC9E
zfoUnTFjmwio5OxP5iHoSgeBPRClYAYMgsUW9orFxv4+Q6fsghb/coDX2uGp2Kx9h38YKDcK1O3H
Qgp3UH97MxpC+h/MZecqvMXRwDEemeZY7NkWxohznj0qPVjGzQKyIGlIS5fe1u4OjRI1dl9To1fa
vhSmoW02tdwfogOsXpOTjo88AZ4F20QyfXSMNBPyDbew0u4quI6OnVzb0aT2vyWCrDEibCC6h77Z
LR8TCGcg2UictYZiEA1ZzRHDG7GMIosG9rwYaVpmTKpq84X08MWp7rIm28qImheilnanbABbkHUk
b+x+zmjdh9wHd7HyQx9IoL3Xghl6kfz54xjJeDCGKXPbKSaJjRPZbJgafYnrPqcg89DCYUCyZTr5
woOVVOnCQ6SenCAy+nmYv2jtBdw58aVSiiFMr+qVpjAXqzmlzyVn5wweua3OBNo54KR8og3r8MNt
a6JBaCvI+KARe0wiXfL/rAbOljauzwxqCbChVl9grn49jDhK5mWYMYd5HXXP3TkGar+cF6CBxuDD
Bk5X9W0bo/IO9iSQPWVUvQRcGtLiQoAxPiwuz0K2LqSBAuIFvthdzBU4OxPllIbdV0cz3cChmYLs
h0Bhdsq60OkrmnFjFgr2FFEkWmhAQd0s7deyna6Ie3YAZfNFeFmOBVMuifPnEwzRUq1oTFXPPzrn
R+1LErAdeC1RK+yHGzFRO3lhBBogMfLi2B1hP+Q4h1UP4DK3v+qO9niz/McJ1AiDdFdhdyZIQNOE
8PiRXYSEHvoENYMuDnsj8WpUw8r99N9XPi9x6c/yXmTty7quYIDYLyGQLv2kxcw+MROZL/kv8+hb
HAhe0AOf8z5bovqBlHQGCYY/0EKQ99AhW5s33zsVE+FBpR7+0dwz3gIuoLmeH6KCXKQw9YvjewIK
jD8dfXnmPmSkmZsur0XN9L7NnyDMyKv5b79YFLscXKI728Bn0BBetHqbffMhK8GZqWnRZeZtx0iM
JaWJUIdhDu5B5oxevFdRPip34tHX3Ln0O+x2om2w+LJpseNlsXMwZjqIdSeUZmlZti5NgPhFDL5M
oDZ8WADruG2apDhrPfzn/bzv2yFe0hG9bboNGI46q9adoNkkGrLoyXH/6iS/qeOQZkJJkDwiJ8dq
+7qH3lnzIoLLR3EE0wi90S+Pq+osfkG9BvNYqVNfgfDHpBdZBCgARPX50daG6Gg6IL7kodMs7Urd
3lETslrY7TyDLdg4aEkhNpRe6SgTdRMRmslsrlKW6sX+Gquos/v+GfIm23jQD3e2S4ZlXiV7erZ2
hK/Q2gBXZ4BNbo9JhLMnyS91OQxK56vRy/qbPCEPJq4kRwyAOrh+/kl634OgOsp+nq26pMjwMpVI
3KHTXP8EZ3lASeVllxvMiTLNNX8HuQXUMkRjNjao1tAupjm7MdMtU2JqrUkvPhvWSRC76yye6BVn
RMX7Bik4ac6xi69Hp5ZNYNJ6Nz6k9rEWl3qax34flzEI7czF4BiwsXWTzS2pMjf81FmRj1kd4eqm
+byl4GJp+JFMV9Sm3TWvQHxCwsxP7RWFCqhAGGElHJRjeBYPKGnwN/nKS7aWb2wNwAsInaYbuyia
oRIjhM2ZTS1PWP9hZc5d6erVGqLGEyXWP/EOfmTSHN2oKXl0JhdXUyyQ31QlGbPTgBYaoU4b3yhE
inKuEdxRlTvRVh/MBe9mD5kla/sy34qrlSntmPe/DGPMnatZZKgaTpqnNFSUuAzhpDd6VqyuG4Uk
Tdq2ZIDZi0DcTvLX7IrftPGGjNXRx8UiqVAkwfMo51Mfc82y7B/xG2WuztLat/wmWyBl6W/Z1jWS
unCMs3YGc7os2x3jUZs7do6lWVpqyy1unmF8RujT2H1E7xt310+60x/u+AiP8NU/PBW9s5Xyx9kZ
Kkr94WuL36O4SocN2TsaP0b8YlfGwuLZ/k58KWCiY0N9LwR35x+5uZbJEJVRW/TwUr0W77GqH2PV
eZxhhASuR19TOCAbpTiwEWz/5qgy1Ck8ZquEpUZFqxC5Ii8HShxzg0dH5UiCDJ7ivroTnVBo0kjy
nxRDZdecGV6VYgQncqeESRfRfPerqyqpqhMSOAPm/u5A6DOEGQKuXHjYvIZuWfsLBqE9xb56jxx7
VL7sgLQurt2qNt1TJiywwph1JAm8vyIqYX5myniMMIiO5Y5hu1XfGNLp8svZ9vT+ZDVK66ii75EZ
QZ/xgU5l8YeTtHycnvKWGgdXURzP8R3y2MBvbNcs35lMQGyNk4jg+PerOM4FkbZGJfNuA7m2fSim
i71zgwsbAtojr//M8vyN+F19MGc7r7mu86xejlJyr6BWMhb5b4fnhQ0sMSMChO8DXb/cQl/ktoXQ
Hq82mNInYFli6CRQpEjjtnTp2zDLzf/liTBoDdEleYYzm8JAgl9kCfpJhWysfic1inyKTwD+xssb
QePxhw9gnFAzFvVJ47D2bb7pHSil6MCkij0Ka/tBkOAQ/qWi20pG9XOgoK26PIWOojcpjp1P6LQe
br0k8hV2bfnlGQyxt/tPd8KTpwozEp2b0uq9V/7YVeEsBg4FV1JiotuigroLv5qjpsiCZS07K0EJ
i2U5gDEy4coC08KN3iCT0SS28cUJzpMpWYMqEYojjIAYxFCklFZ9sjhgmiJsD6AfLx2uXoLqWuwB
RvvVd1BTmTk6u/rD7U0h2QFh3ZZz7O0AWmcMCpYRNGHdKiZfdLLOMoRdq8LBONeE2JJPSv8sa1ca
DKeGYS+8ZYUZAbzDckvhxK6aIGSe4yuR76WArRAgagzs+cTIT7PG3Sy3wQxJga2KSA5C5JKTCHrt
FAqlao3FEy1ptHbVcCyN/buaQiDWdNJh3hZVspGMAPDIkzJS5K1YRiXRXi1bTj7YYRDpNExzZQY7
3sgXyUxLrCWnL6LcaHLT+m2ntcVTbRREZvGeb/njJC/lnvacGMUtkXtjSLIplA6k21M3rYqOPPAT
ekqeADzSJZ81L1IVzzPJd9hq5aA4j/Gj7wZdwj7Oj3w3eePw1vixCvnFhMxIVxo2V2ZJ7KA61MJZ
Er1vGou50S//8ROyxf1D0kWElgTxVV292M1vyJeW3h5tmNSbkuT6C2AGbupPYNZEDN0h2RaeYs2y
svkPmSeT2zpKMHOcSG3eQuOvaqd3gOG/YP3Ka/pD+GkY/XxxmNJJkBQ7BFbWClaPx4j35GEePYsa
muN2ZmUKSiBJLiAdzF6zvCI83544Nnghhmo4oJcJ1JvPz0cipS/5rhD/2tG2yzfZy/Rgv4t2IBj+
KfC+GubSK+J/CoJspzGT3qToLuahdSUM7zhjzz/R5SM4F+4nL5+eAP5y9C4ODx3sBsiZQQOyP2dR
xLtNNV6H5+U8YDHINiqkUxU8Mbq55q/0pRH5TAd/yDgS/4PqUsVc+0Xy6fw3eYyoLnYVwelar1/z
bisjY+vRMZFgSZ4uc/e35UfiF972sx/q53GGRCW+QuhYKFZWDs7rcYc+FR52Xl2Y3GhPTpuy88lE
DttqFCR2sp9Jns+sv0t1UUlDvZt2lGgoXBGuEAjxHGBpJz2fJSkAgB+BV+mZ5XIj3GVEUFKS21EK
URETquloH7/2N1Nk+w0oH1/RTigRgRTSDsm3Dm07HqmzENua5FKs8JgwP/xWodRlAthSIMBMpFIV
iMLIa6BDHswmxuWn+5FHm3rLWeYq1n+LfDr0JX0r+zv2Cbj3IIF97m3IbDpbcFe5JLw0gpMI2k04
xtT6LGw+ddbgHsOUVOjj8PJr5SuTyX4rkYaUPkEzB42noKk0dZyK1LHG0tMbLdmW95NRjTMwEz4u
D6Awd+dbPdk53km7cUMCIXRPDbnnMjRnTQkKpdNvX6Hv7uNCap1Syawa1zXsrOv5J7cxp+DF65/j
tliDKVd15VB/0sJATBV7uRrHCbEFUhX4uIRpC4edNkebQOpf+Rxvs/iKxOLas2a2OUOr3qaxJJWs
LCJSHhVBJU0UT6EQu2uJoLab7Wj6tA8s/pHQP0n9cFJlodYTczzhVWqUtemjYYecKl8YC2+5jbuT
iYErQCg9rUltDIpDbwysg994kulUWWRfGncO0toblqmau287P4EZQ2I3B6A7HHo27sxDr3i7PbuJ
O+mEGpbbbOX88O+XJd0PHFvK5MtWsSWHbe/Z7acMW03a3HMdqajOsGCBX87zdvjXdNDyuJpnsQ9v
j8l865wVnp7Bvw/t+n3+bCkJlflqDDYo4AUSxCYT1RlNgj3QEL0ovphad3vW734e+wSxYKpfpVIb
3X6BijyY19Kllsya3o5FET4eXGtWgsRB1DNuiV4B2UJ+RUNcPhT8LZ8HYDcqEMDg7ofSD5SDD9Z9
HyPq9a2y7m4LpqUM3WYyiym2l70uBa1MCGIYEowmI6BWjYgjbJcKXLnkrBx4taa0diESJfyXA74a
PAYwW5ERCFZ7ueRuGTpyOkQBt3dpt5FedBB8cxjFRZPTkL3N+Lwu4H0d/sprO9+mcbH+gRU3nv3H
r7Z3NeTNDYd6GvNXf/Amg3giwBNnDhDWdFMa/vtfB1LNz2+zFr1SDYDtGC7eabe+ILZNfXVmYmII
MfaFCXfOeIFzueqnnttB1qJWpSbcvGr59TRR7AHBizxj9O/no5wDwp2JlFjx4wJYlHCkkFtts9ij
9nDONxGoDYS9hQr43hUQkLbb6XEfj2B/20EzvPH6ZG0GPCC32jO73t9yffcneoZQPFRsBmfKeyyU
cv2eMnlSYl8d2vbsmbbIpGFDYERji5f69v5GwR5/mDDWUOWHLCaW9PidTw2PfknniD3AAvAxg9+8
zc01UJ4vKA8gjhWoBwie38qWwXV119LXHLDrwA4uzLMhNID8uDAqojGWQzhnyL12KrvOP1XLQUvO
IamE1c9o4qE8p1G7Rw/+viIlFYY2Db5Yn0jcvS1GzIe20+d3OTGFhykQ7+YnbNQAhHtDHk0hx2Gv
Ysr2W72Q+sH4XRHq/md3h2xETnjFxQaWmZlg8OJBc+SZPkusO5bsyNJygyKzOTJCB4I3YTsk6sZo
RWCH0vVywIamAFkURTwU3WbeGRgnfmUbFU/D0iBfjmTSIVgtcrRWd5aqGtNkxHF02y5ODWLQ92wP
gvXESZYp8xxXUTkL/l4xNvZMKtL7n5dOGtRpyjUfpEcWDi2htEeorSAArX9rTIuydaRBwNG1v+IT
Phib9OtVhgy3jSmBg9I+VGzukc+gB1e+ecpAh1Q7+/9907KHaRz9PBIe2/cb7Y/2PY49RMfi8rA9
sl4HqWu2MAq7Rhf5ZTWgnTholCOP4hsITbwuEEDW6q4cMNMifMKFzLDBhwbi6Z7wE7sW8Qv9k0cp
SqB2rz60zuUGZOe63OZT1qDAkRnFbsJC+pZmjs7EHTRCum3BczOU0XHc3JOm5Hu2cNuNdn0GdIkI
NbJlT/CqxU/0OKZNvhR4vL8XC/MTTPzT0nBQUgyKxEpd0f7x82jFVj3IOuuaSLkJHc+vkRFIbG42
AX+XJBNhLYfN89cIz7jqzVUeJGe/dkfx7+F6QjE4ExM2Q6Ukyzp0u/h27v2jr4uevIGXudh/H5+b
ZUCJTHCCr5goF6nVyr7MiuHWmnnuRyQZe/dFy508dJIMu5Hk64drK0XsEX1Rs4stLWDHkwTGvxfL
B+e3+JtLFwyCeUTL9mhp9dachL63S9LMon1tUcYQK/8EW9NmrfssaCY/yriPNZ5BheVAov2hyYlw
nW54vlCWD1RY62qCkzoodjIpkS0OLdz3raNFA+/6OUQOiurogXq24lbKVGFqRJumhUgbFovsL1wn
RQhnj/2Y7mDpU2nKCB9+EPZIiCMToyGdczYsujFIcpWt88O62S5/zI8QNq3MP5QakaNOhXY1uiRB
pZJSdGXz5f0uzpdeaFDwz8X37tO1dQsvYL4iYpntHLhc23jOD0c7NFbXjzhgqsLKJiiNjU3PEg7u
yH1+8dhEJ2EYHVyAsDd696Nw/RFhoXbIxOxvLUFm4MUECTpIRhRR0CRN+7K9ByBEA9vBdGOq0b93
++uAqDww6Y5W9q5lMw6EIpNkAw+SdLrnz+h9rZF9fT17wdXfQ6lg8dYjDQ2qTyCDNozyjrS56xVP
JJOBokFSm3zWaATBCElM68e0Fui6QOXiMD2pfpYMa7HIBz0VSvcEd0Y0/bSIA/aQ9S1p9IFyBYpH
OGX0hw2nVX7I7Q4H2HO4hcNHDD7MkmxrJOliH0GP2B7BDVVLUMPY80sXzeYrkGmlA8v8axgoSnoS
rKw1WAzRr6rYKgcyTwHBZtBuC1wYR8wdGJssf639aCG3u5RVNkO0PiRYoKV3hU/Y23+sznk5l7rL
+c7k200tTCjExe1VWGFj43yezZeJJE7t8GrIJHk3dkHZ7xrYtBhsxDwmA3o1ZftGRby/jNmrpBKY
OZpuO3IsPjCoFK3WcsPcwkrBwJ6MYt7711did4pW/6Baek1yn9qVudc3aGd+07F2cQ9jgwW/3has
Wfpv4CCJRogomtj73QpvBnife7odwoT3tINKPg57huEr+Xyc+FI1V/4xXToSWt4JABqKv3v3SH9m
2Au2+9KdexAGr+BTL+w18EYmjoupce3IhdjSKfN3LBa4EmyFr/HQaUCJaahwFVku2e2IBrnHoy51
g1PTOr6VYHxmmmWErFUU1bGm5oQYz6GGGcyCgwncIPwqzd7UVG+mfMJk0d6lEdJGfRgMKppivatD
j6yfUfXBmA4pA9UwqA6aGq0TSWUQ3i5khF+c+tuVxySOAOWgEOvxJcqihNQ2VFqyjaBMZDHtvaBu
zoougzI4ngHi23YMpwMXVey3bMnwI04vh//shCOJD8R8H8I7LQBNNI3cq/oQHc+A4+Z1k1KI6TPY
WlJbBaegRfhc89+ctMpvWwEryQ/GFiDvHV9MOKttSqOD3mA3Uv5XLF5WQw4LAYjFN9CQ17m1PxyT
wriRYfdxneA+ylf2tSAm6xfnXhaff1cjXh2H9M28y6vyQi/LcIWcSZnttX5F+ChgESvyfiOfdfWS
ROvsq5kl6f7fdM6vC/0jHlgJ+oaQ3MEtroFYlCWpx+Jwa1FYRyQCkyOBxyRVOdEPp2l7bCAdw3SR
+HEEiK9tBvICYGEcMuMrvA/y+wSl8Ga3Mearp7j4cUiiOAdV9T0evOPSbDyFfFnqSUIEWBmqozhs
pucyYRQVOxGuT/asLQrYe29jNvQEBUFwqMiGf75+qo/YwP1FgaXzBG6FMIceG9/YAoUn38j3rIWm
MV1g3xSC7EDf8TvzuPcy3UQAKNAHwrN9ydNL8aW6AkzSnSNvXohDktseNQ86E5g7kHO31FeP0Tww
zVbFbntDFOANcXQY3GO5avrJonv+ltxHM+XI2yX6t0dUllNHILWoOZ54n7KMSj8RZNReMHvc4mev
j6KUnGcZUJFgLbCXhjtphsUxwFzmiSnnUrTVZuB2yu+zhh3Sz+WwvypaEtOBiLDiI6iXFkYQxMeu
Ns7KmUY2zRgxnS2isOaNQ72aP0I3ElQXsln+CtrceeGhXjhR4IU2pFcf+KztrTFHI2AZRWMaK/Pq
cOXuechM7EwFxtrU1vXo6TdI6y0f7kpGKuUuK7K7HaLMaVHY/iMENaYKppFqYdw8Ldrk5NPSnm4M
XgVqVpWGZ3WDEnyRsVIYPBVD/gmAq+OSIru+T9edn/npEULgnKZIjzVHPOsn/NBN498/bwTZqaty
bsEzHZ9N2pEtQqtxqM+qKrObiv0ndPhSoaBy66BU9e/QR6K2aREQwOONZBZy7QeWNILvurHxpu1w
n0rZonkH6FaVm/6JPLk/RfiIizz0alU6EQ5642d488j3k3lo4Zgt1KUYThJjSCBgexABa9QaLS/P
44A7nflg4XeHrI3fM4cy3bNElJvRW4G1nV95ORhTMVrZNo2Zo6m0n8HZw49zrY/LdLna2qVP940h
cthZhSUlKfx1IzZjpJHU+i9i5Io+OZcSVQ/S4LtcTAN+N7cqpeshAslB2Ik4O5bM26GlNZQ/K6Ey
yKdXZK5IhC6ie+EfN2wWLO2Mr7cq8VK+zz6DKyV/IqpX0YHQuhScXXnVwxnAVQGBHUXcX/8zLFpi
mxm2tULLCrMC66v1EPzq53eIk83jtBf8BnjInXDnf4BK4pu9Pa0BsZv0JIyvnTA/aReQ/064Sfwd
a0kyBpJt2yP+Q4i1dPSnaqYi70M3jlakUvuwBnY8YiWe/59HBpLiBy9bMDHA83VYXsYPC9POdbLN
LnIZ22FO+22vSPVbtwqVk8q2ypMdlHA58pDusS5E5Vb9kWH2bFZwlL+f1X/jXZPief0beUoXqM/Z
E4rAx7E31uDnPaZ7Ni3zTTVecfPNIPgbtBFWHu/wepHhiOIJ/Y8ckuNwWWnJxqzORFtrQgEZRe8B
TKTkIHFQ9xQjeCdtMbrVJN2evjeneA+wf5PyCX8e6RYdC2KfzW1gnYKhrGd/MOpvqRPsqB79ZfAB
nsFQgOQZoEQ96zVcxNo30dyh0ph5yyD32Ns4I0LMsUvYblrfAf3hQwtRyy2kyWrbbcrH1qFaCF69
rdRvezqWB29wH12q1vbLxnH0HX4Cr1/TfoMAKz+R7fHXd3jcbgj28azTQdfUHP36LBLthkg43SGH
khD3+9fjEQYAtfejfmHiG1dBUckKj46YqIX70xF+OynUVzcAUT/KTHZwbNi9fLIID5/Rfif8roqE
xdTvUeLqDGtKE/XI9dIAQKLTxmvYrjP+g4oedBhIlpL2gC4y3lbRh8t+drDGOREYLBgH5oArH/Oi
D+H+qB7bAGuMZIC0v9ChxzwQ0PzxAfyWJRMETmenscopD+xtm0BMDwo60FWnaytujEJw7YTTHM4j
gI6fABTPylzIkP25vbd8LWHdxCpup6Jd6VstcbFX8uSKwnQz/X1mSZz2x8u129y0jYAjfxvd+Ior
cJM1vyxBfxaJckO806kltA3LbsDZPUv89zvdqQB6uohrIJmmbwzmYwzeQJTa13TzfJCS59fII+hP
2Pev8UaQVDavm7YZDGfmwmJ9IDYN1e5DFlYB/q4Y5Vt4IOy+VijsoyImT7azPXjKTt4DbeMJV05F
dzQ9d1L0AJ4JrqBdtuJtc6mvsyPsDmHQA1NyuT5z9HL0THHpKfS61d/rOmUW6kbjuvWW+6VtLZVn
B7j0tPO6sZNwPQv1SzL3Kcezwl51v9kDciQQ+kBGYpOSQM9g7ut+jgeA0FN4yXkacO0+Jaz5rohO
lYje0EDBrq/dp6ebQ0m5thlDImhaBVtRQvCFf4KLfg0vOYM6T+2v+EakmjXizhRrNkgcR2QeqTQ8
z9RUlUCTwyBB1f9Hd/z0Ai+RF1snwZT69lKiI5NcA9CoF5zn6hR9UdBQOcCFyHiEPhh3+D4ere2U
g3rEfk5RHfbvKat2OZ5XzO18INQ9sT9rxZ5gNtyEiqrfHrWNyuFWNxu+G72gvWcn95Rl/eY156+U
84lVTrCh31aw+yqjL2BvGJWzNakkjDZowPcyX1xvMoaPLLV/Py4Or08u9Z3H4+0U78G4JSEHk/KE
A00RTGGf+49fXCxZOcJ/0AtxXLq1v3POw0CTPQc5sQyTyzqVOrf2aGF4Ahihoz+e4tzjVuIl10Qb
MlIn6UOSItqnayHY2gJBM4LsmA0WAbA/8LWNEpVoOc1mGvLs1tlj/CaHcW2ZaRuxkb+xvSiESNyF
pmQucbbBvRN5Dg4atuWgNUICu1/ilXB+89D+GIy0k4wEDcY5hqlUm//1o8noQYX+pWTzMTvK5IP+
fIpFMgVQDCPcgHVrQ5CJVWKFebjbWul66ZfF8Wibaeq/2NFssAsN8VfHyBb6PRf48+b2izWTAHLm
KNg5gJhJpuzAbHbxPMwvMSQwj+MMmXMYuiVb3ESFhNoFt6o3AeEwWbHEEt7+W9J3lL6dhRnMdmbz
4oA0xc6bQRwVe9fj2S6Xqr0g+CNbRKRPWreIyflYsQL+m9OqTgg6PCpm2GTFiwNN3YkoIjJNWEek
xSLwEi6mUgqrtUu4WJ+6BEuuV8qk1DP08gYNsg2KlU9vJUp65T+5+RBHaxA+by9LWJs375UAn5KC
TkYo1iyn4Is/W21ePNlDZPqsdVGU+zKYCfx2wt7jGItSulyQSOOH74y2J0hmQ+TWtSzk+alT3mcK
VXFSdUUB4FmvZSJ6VXE70rAZwG1pxVlP04nui+rsg6Xq3D5cMrbj6huaaVav6r7D9y2LdFBoXGj4
jRXIYwckeYm6czWPFHK1Kun7ymrVob3HPyZf/c4QmfOJDzv+X4YVmjgNqqMclG5qmi6A43dKm9/W
nFmrcCDgvfG6EJ07RMDjLyT7wipUH3JiRSQX/gfy1l3cNXhlrLsMOW7wul+Wq9Vt7F5dyqRzO8Ya
ACUXf2HDWSk5eWRKNTceIS3WxkeOSC5B644a+11wvl+4Rzhl1coubOu6/vJh423vaI8Y15yjdSzb
Z5QmEA+bhNVtAZD7JHn3pbswTy1XnZ2LUUclyfCD1qDZ+XbTg1JOY02RUwnmApMndCBDyUpOK2nf
8tmLVB+A7gOwtDXtMRhhTynqReH96wr+V6IsSkyV495w4r0Djbr3oe4yL89Uimjz4Z3zw0jue6n7
qS/CrRFNIxr6/KiXMWqBT7AB5A92W7zjHPRLPpm+I8hky/lmV/UOaQJhzhLmPWQL2GJFyjIKU0qq
z6RbDO3WDJBavjdI0o7DUTSlHD0OeI/quNmr6qqU3HN7E7ZRl2lrngUBd7tW2AKEOL7jNM5ReWxX
A7Ra269I/qNATsLOx1wsoLaSuxNM0M/UlQolBpsIvauWPlJIHWsOLWJGvyhYy2vNSXN2uS1OHeue
mldoC0gSmrzwI/vGgfTNm9s2bGfMO0LnYgNaakYA10CgdNomHJQhs6s4lVnArHa4Pb6CsG/hEwDE
3SQZir71jdJZLwL1Fp9D0HyzR8N096ciuyKtMaR3jp/UGspdHocm+0tSLpRnsPddMfx5dXI7CpSm
8ogS+6mXl7+0P5OLTnEaJYlEcP18O9XUJXS95CAPo5zqsw59wSaeOM1waacBt/sE37leEztgags+
C1KdQnD8HmjDlO6stwHfVbng8pLrddOYdhp6ObGhW06KY4DDQeo0z8yn/qhYC3z6mG6SKXsrxiov
M27w8nZPBmZsux6Jdx8PwDI3i9C2fQXy77HJzNEVjdGw/PHahBfUCBw0vZm/UtzOCAZum8EzF62b
eMxo/HXe9e76hq4kd8H3H90M+Hicwgnvj1RaBWNnzVt1oqm4aqOu46+qwYvZOE5wNzcmuyJOMMsl
jjmoTuF8OsN0NNc06EWIESZTn5BxFr8WfwHT6RQjCVODiCnWPLA8nPU+fUkz8mmGLf1wm2A1wNRR
n05SeNqMQIFmJqPceIwp7hf/oK5SJurFDfuk74C5oiYWAasAg92IawIp6b7WEJkmkqaXVogSvt5S
PLYousl+uv/zvhYrJGoB/GZSRZo+GQTU+5t7DX/PhbP8YxaCHn+HPyF1iaXnRPDeAfZeipIUp0wo
qlOOZSFJefTP/fnfaFzc3VGNUNhl5lYTSDfbO36HrBAoiRnoBZBn8nnVds5FgjUtpUSETUA/BDU8
F2CJpR6bQb+6yWuiezojERtnTdDBAWpHnWXrUkV6lYxMfSp1lF7OZP6J9X+fF0WetXV9YmgUBP5h
4BQS8HjmGhyW8cfefiziSeu7oqr6u9gfyBxUGVTtyDxYYQmGjZkfoKSa1pZR1ymP6jfMWJO8e2rR
GMFFfxaewMuQm1L+O1ziD/+r3BO4uoGB4SQ2YWY8Ura2zcQxR3LkBYp0lBG2/xIefx/v9zy1W+AS
9l0K8Z92lEZsHJiTmpd91FECYMccgM/0FrWG0oec9Y+mf1AsY3UPoyH2gaheILlbB4q1jpjEjpbI
DYNuqiQUB3dik4ihpumolBUkJjEEXiZZ3HIA0VZKpZ2AW0HkKilB3Fpd++1r8bu1QtkxHioQWdVR
ttUF1rMI4FEdwND/IYSX+fVXDlp7RK8cIaEwgODNVnVwBcyV7auogqtVBppJigotYlVw2p7JAcZD
p0r74RMtmjWOCDsbTqn+8gheSZHRHzw5FnMcwJFcAlO6D+bqqJn85qpCVhGwY3GiLOxynbPibREk
nGI4WYoFBmXajsjqcoysHtrxEiEiDQjDhmYghBu9oHC0IGfo2Onyp9/drdwy+MFX86jUhGDMZnsR
jzUeD2ZFs+03qBOpxq/v0d0JN21otk44oH+d1byKxvERi0Go8+j7TaYM8LVO1i/tdil7jN2n47zR
acRULl3tzQREHBRw0xBlyMUo9nmWzRRxWK9nQBofOv6zmeUYQUFxKVpxLorCZxUP0VZs2RdNdFvW
+FX1gN77q+2I1BxtGLbYEaWkMp2P4s4ybJARDIXhP9ndTL0dAejojiFvzbtttxPdXdw1BdtZq4pK
xS41BMP66sew7qG2tJSyEPHb9VXvYXFidA0Q9EVpc0eUfOTrJS1oMpcXr0N8cD3Jf2IJQaWDtT4h
sfLdoasUpbsgVdc/Ho7mZwoIx1o+uy1iDnp7qUNBE6HjDVir/DvctG07WW+tFVzqDfx6b8Mkyz/f
gxJs5FG0h0HT3K0GiAnZ/m74Ei3UtLptLI6npKARKE7ApHl86FOrdWwNP+VnqoecbrAgutAQD4p7
pXT2MvrQwJKlYQ/R9XwZNi7bjaThrUDKefUzJG1v0gdlBwchTgHLgHOQb41fE0+2HJSJqS+1qjSD
cakizY9lgMlyoRiqgTQLTW9IJ4aqdF0MzpIvFXNQCUjeASCZCWyZ3HMebdUQd1DxRX0oe16ovJTS
aESyj9wDX93hYx6x4SfPR9H28kRoG4/RVU2BcfDyZtSiXudc8Yz40A9GcfmGNisXu3ZTM7rfFS8a
vLoGEunOgmRZGLf2x0+/r4x3MnMjDMQFWQ+7km1wpoKbvNQ4pQTxP7vW5gN5dW7x6kFTmeEFCQAm
HJWKrvkqW0tIucyWKonPBtfRU+PQ+Ryh1RX8Z3oO9QFGGXjyBJLLuBCsGZUfewaGXPSa5LO8YheO
OC6gVmBRWA+11DCVDHDz20WEppOORCrKBWW4yIxCGSE69Y2EXgrMb/DWLRBxSqdmfNBL1E/ZpWDp
4KDVEEijte6+2sgDEyBFKjBJyIBG3oU5TBKe/FznJ6ebyANa+oM3SaPYGqPFrV1I8/DexkFKR2M1
khNHLLeYxa3gSoZRIJNTINeaP8C95pU7+XlIeIBI9aB4TytEOof/6r/L+xNUHaYZrsmRmMB73J7X
ZM4pvGWryt6LGdjpmM7kb9Lb864dIkNS8WOJOE22CBcSIod6d9SJpr5GuhyfeVt0xH1Uv08jAMkM
6VmRu3n7JUfUcsfXC+jJhSoQTBI4L0RJ7PhlwmFuqLju9h+2x5P/m1JVGihp+D6OQIpDOIKbZMjN
7hVRmewstpyFqv4vMO8PgkV3Nn+ArafhtA0OrYstJEJCFizl42WqRrX6bf77Q6feo8zsFgqEhBZ6
pbLhGQKL0tHm7j599QIwKr2c3+4UeaUa9WieDg0YZYu/1UhZS+QSZBujOMmVzwEjpWORr2vBpkJA
iQfGO1o/hDwJaOzDX2YHhfoZPnTdpOghEAXbm3K8STzmrXFwhqbJeAAeikfOo/ja/7N2WMvfusMX
lqlPRvnEY2h3jJtg2hEc+X0datgOsChJOAUdJAGKPIV7/ZiB+kams+lUEXdKeSx4mGYGTq1kpiZI
/ZWmnegEINSgqlYmtSdv9GGPy7jcqi+tV7iJySaD7itVKPxX60Bq3zbVH71pisQ1Vf+nkFAqzZY5
0pGtCk7Dy4nXNqlFBWRr5IVEzhI0ZfbXLGQT3MQxS8qnJZqSeHCYtAYjEiOheym5Wx7RFTDrKwsn
ZFpQme+6NMk7KRv5qRNXlpRubHUxx2WfO/rDIc5/yXKs9RJiFAfETGqLGNJfDaU5Z+hZ88zqCECe
JG2Uc3WzgIdxU/hB8bG3XIB1gjZ3F8QmU1ABLmQFFyqmSdTHWbyFTmyEfoTMlLNcsPZOJMuzHlYd
VeqJ/KDWIR4tIEyW1dtL7W3OktqsjBcS2x14ZeKFu+mxAgWqvGsaYsr5eTFG5VUHhtoKRBPNOTod
9v+899+3vK2wES1KugU3LvFP7w2myp8HTsxaz7oLlvQBWgyzuVrisidAy/2J2cFUdDi7tGOO3qIM
FaKjhgTLiVTN8fcWkKv7yfSy2TfiJZBGB/K50or+94eufIE3WXv6/oxxyNLgUlJ6eHoY3S8p6Wd4
uoMtShrTyrPDt9Jk2PVzLDSQ/gR0Y6ZiReoy3BPTigtb6IwkF2+TRXjPi7O3ZsjieQ7zvRizWE3j
C5VQk8u7qtTI8VRHKJSfrlCO0vX6I1nGCPHC5DamwYvEVS01xAJ5uYXrKzRiOEcUzHrGaWzJmar9
tuAFJAcyn5dbra7hMpvfLgsGMR8xk/ZMzHIqgOHNS3W3h70BjgzZvw7NEgIz4VRJonz4nmEt5c0L
AFMiWNuClvmnvKMK8vOTYHVuHHGgXQVCMeNVgcxnMEr9qvQCYdd8FjatEeZHvxB57e7nUxV13EpM
nHXzKg5JL+cCVrrvMiiqZLvpVjzMacOUXP3MqqEih8Fh4dO+GKqE30FNZ0bTLOoEykp0s7Fn5Hox
b+YbwDMDqqQnfcMF39S9feSlr3G7ttZLV3VTiH+ewwv+VMv73DFPyHhpTKGBhjBd4Yn+4EFfY5KE
brLVxMg6zepMLgwgVDE2J5+1BFl7vUCY19KAimwyCT1QZdTsCSsto2Bn2NAJ+r2DVpIHJ6N23DZU
uHqadYM+uQyIXdZyIA3iw5fTiQtjuz/M7nnD3Yc2CyqAk4zgoLy/Jn5YbNq0BDYlPg3uRj1IGE9k
5ZK8paZwyLmPOU520zULHpQDlana51LQoZ8bz+aAetjZ1QsnU3nGrBqA5qy+XeWsx4GXyeJLqXZa
pV+gnLeqkI2VID20RV5XAPdvrHHBajVvcqAAJj6VxhXRmzodf8rwz+P/EUUSQm/BPe7n4TKt1E1k
Lx2jGw6ZOYJzMraP5Qf3B3Uu7C7TcV9RuAPIkM42FnG1F5ZRGSh47/XcglUyr9CHguREzU0Jbzr2
OpNjFNyW/cJEfisMNDMx164g6R4BxoyQIoBckOwX1TDE8D3Sq8P5e3sE8BRcepSssgpSWafONz4p
EwAZ4wK7ZsaVc3lAo8nVLPVmdsMaKyUOKUlrC9mMiMpPal9owac1vssV80Py6I+mLUNa2CGck5pp
IoBgQMPakSOD6yFUJkwSKwvxJ0UlPRx8jimGd1aSvzFkNqRuX+oPKjV2Tq3ytKGKV/wfSjkGXv9D
E0in2Zo1di3UUxyPfo3YFi94LIESsKoVA+ePm4dd2pKS+Yflz0Hr+vg2QCyzKmL5faIa31qb5nMS
dDcHlR21V030FakqC0PHItb3Kc311sYScoee+f5grYMCDN3ulIwTeRomxNMHHJC+L+RdfmCzNvK1
l/Z0W8uhrpLZAox0163w2KC0T/KdRRMGv1n4uyE0E3O5FAgjnVqE0PWLcQa0SiG3kl5EJ7n/VRLQ
wZn9yUV7uD8X0ilI12y7eZnlKNN4FX93i4ygL5FNbmrzLmIFfTo4Su4039zpoYCvWRJ2XGMOPDty
Qv0a6eIIJ2jxcq5MCVqM2GzPenQRdUKMw/ponCISCqGWSivxEss/Xlpp1O6q4v/mYmqIvJDZqZlU
aFtkTZV63ieJd9WU1HCHdLh8TLZ381P58WlQqbME+7e717O8Gd5CHcjw2KOHDBe4KxL4Tac/0Ag2
IUeD6odVmzSBRpGmVtvoaI/sjsaLXVwFpz7WIjSn+FxkQOI67EbMFafzDhyGkb+qynMTYPOcTz4n
eQoEeECLK91A3fDfVIcb/CkFfUKxlgsee/VZeUXbgNEMTXah83ro64632RGMyZqjO9z5U/RG09Lv
y5TrW3/aUO6nyphtzmcZpsaRPKhdOeoDmYHy66uMFSnpCO3nDYYaJHtoq3btFgx4Ih9aV2OxHt3x
biuGolOz5hi8CwM6ALdidj3YyHHKYfza9olvmIY8AFNst+E/HhPtpKOkHYdFNWegMu7T01TNteXr
AbmqSHHWT1afXW/69XhaNP6FZkLRutr3WpZwznVK5SwQHUGMDDuxExTXWQOKTPLxKmmON57XoXvo
UsAzhLdLFz3coqK/3ioXgsBR6ucAmv/nH8utbjzl4Sjm138qHvl3oJO6Dvd9uyCrwTK4E/c+htTS
UJhCFDbLpRhVUAgpWkFlyTWX0+oq9KTKBQuZUeK9Pygbj6SbzHz1vx1Y1Ev9Bt3LqMBfFekQmuxc
DjPoR706g81sao0a5E4Z36GCg4E1QO1j78pnYjewppxaGBKfIw9mdMrDsYdCOxAnpAlf3UZWJLjY
kZdrY2g5Eq9rtOHlXyfsPN9g7yiPxamRUy3E/nNmXpP7za3uQvRCYWklDrsx2IJAuvTb99Ohvi7o
a3M7CzC3fYmxwpqS54xPp+6mLi7xzBVGV6J1P4paBz9EDDHMqPDBJnNXQM/Ytz8TZYraNtrvECKP
ADREgef8BM056y5XLpuS+HXSz+WoWqHJ+gzdmpKZL/1st2tGl/mvAitvM71KKAjqjOVwvd3BlXHb
YkeFrSE4HrgJ0KeJ5k/W+FvGqj1IwYOWc3Y4Ug7ZLX3ZqIRBxaIJ0xAZapvgIxgYir2NegII9HTD
i7VLBFUGskkd2ocUpEt3X5oZ+Cx4MgDMeQMI+CLzRjD+Y7aojjyQ1/Cx8otL2EKq7T8mdv3nwXU8
IprsoUOZ63aSJHSzOG2Yg1hmZKQHHi4dCnVnBcS8EIX13iNklHh50E0yCHjlsqXUffpUBK3HG2dc
x9vicPJtzTXOMsLyPjxTvYZKOV4Bk4+cR1FNSiyp5GWtJa0AAcmMIkYtm5d0wgyBpPb8llViqRZp
StwUM0rQiUS80ml19oT4+cQSfGnvbXmXHbMX3Yqt9C+v4KSrEDOJ3xsT1Q+r9OXIQnfhUF0j6lQS
OmIwx4o0Sd/15dVtETTAxP4pVlHV1XWLykQZyh20oLzy3JIBTJJZHkEN+AYTJpILKIBqd0Q2f+PP
OHvHnaXSgJeEpwOdActrxFI4WFty27sFSygC8ewJHNx/MhxDXBxTmWPxsxi7nTRCrvxCeNNxNFFn
++uWKVglNyRm7646d7d1uoiH9QDJmBDKyGkvwK4/QR92wtxpoJ0dv82rRDgM9rQeY7/UNmntAsnL
OVdL/3kIO1sMOtk7sGPflfKZK8gTLLRUdY+7mHxUzQD2AOQaTIQKa6t7xnblteaE3QoIg4pub0RC
zGyuIhu+gHUCmpEcb2WDPmvAFY5uMP+YUrQMwpoA4Gb7jSglrw8IxaqIkaEvkmj/cwdpMazYzFZ3
3HTVHiNTTOKJ2rhRZitR1tXws/DeIGPs/ywvmRkYsWxpJCgyqy1MzRSG4RWaDHNTLK3BDk375Cfi
HKSR70H7ndXaoDwrSjZ4osL3wqayiyBcdAm6CqdDbbrp69bhcAiLmf7kJuVxIDQlLepJhjyKhs07
qOjMufVhDAE9v5+9kfJqeVYN5tobWSZnrR1l4vEc+MaxiQYF8fqGIEhdAOL92bWl4eedC1gITErK
9bhDWivuxbabl2/Q8GQViAr3t4ry/Gh/Z0LDkxlNH4IW8vtxpKuqBTK11T9qLsfP7njvwMg6tduC
gQTjWB42AGQmGeRmAP1dswBteCEE5ZRvBi/5Xd0wW+Durx9j87Dt7OEnSFWIu3jH/Fmnrzf7wumL
uM+PBs0gfk+TY/dLfpvi43XRIp3c8qgsfVq4PfRDxsH7eC0zISJLi2ZHCl95JWkOfHtsxLMYFJZ+
Yf6qtCvBf1X1K8MZZGQVCg45hfQJw9aj4XEfJ0usX14tBTqDFtOd4ZTrvU2hbRNGBKXEEx7U5IVU
nUUB6rRqmwaTdUZ3JlUqAM+6HISYGN9TUQXgy8DZxaQmUm14a4qHUmUdtxOmX/rbVcI8jKBOZSh3
QWIlD5S/C4bZ/9QrtBt9PVnbm8Csz/YZpD1TDWywRjexjSx/ljqeWV6Zy72Af5f6MnZGaFUTKdal
G6CSYp/5HC63+uMx5kRPwS3V0Y5NNIq7EEUxFJR2hSu3IgDa1DUsX01s4m1Nj1laSz5IAtlOcfY1
0IEzvSDPZ3zIAT08U/Erh8Y1fDBnUdoJymWsVtNn7Rc/w/EQJBbOOnqGKtMHd9IZ5TJ8Rl8a3vPA
GO8OhJWfujFQWw0XyrBgcgN7jD+9YFeS4CzP8xJD8j/YipTuUSL8QMkJBW0Yb9ibR4nZFeoDOFNQ
+j1uuZ2/X2bWR03GycKjF5YHirgPkxFYX8V5Oc961Si7xSsOiJ+3PuiWh6oMX/SPy/Blvap1f7mJ
9Y0ZYuoscvx8CE2zKHf4wLtNZO5CoKL4m6+odZvO7deU7Qmbs/Hs1DPks5CZJ9OX6OWdZQt3m4tS
l2ieapu2pNLobanhf0EnveOQ2cMPdG1u1y6EKT5p/6ynsarEOuVObj5i4+4C9Ye9omRUWWpj4spe
MEYS5HKGQdGSsgg4TLL45qmjtPeC3PHKkhoieOSqIyGaP7aDSkXMvN6+HD+b6NlhnL8xU7LdpLvp
9DPBroXNVto69ezvD+c9V5XFRNFp/qSf/OT7qXP5tABDTP0rRHlvv7yT61MfSbk7PhybAkT19Z2p
UdtJ9UgVUB5j08Gg12hQ93rey+91XTFH+1ZbyydjfWXQtLeaBgzZQf4bAnE6Xgb4Q0UXluao32WE
hwlFm4I7VjrFOp0ddlImAUS89V4i6YzzEMXFDlCeXSjuCrpJ1wUX7TZk0H9iN1D913OChP3xU2T0
kMsKFzfl2rToVF+nNnJBSRm4iHciQg7UwVmlwukg0oDkFKlqLAlb3VwOeF8R125/j/Zu3o7S8t23
BU0dxUhWa379bePu5W6cggW0r43eB68TKeGcXg1THZjxa+xYp9Od+rFWrxgNOg6bqyJQJx23vXai
HB/Wr3LGyy/wQI3b6secZ0clWFwrlzrJhVR+9EkUQVq2sfbYBFCVtqqXuZxiklOXlBjXTe7bqhnX
2bgX3MA5v7UvmH7CpnGcL1NN+gZ3lwA6b/y3vpLditwwnUp2INLFfpUg1uPCMgZG3SN3+J7k0My6
Jcx0bRZi6cNFU9fBy2Kz2loN2DgQvilEIxncFLC50eAmxiF5lcKLhVNCN1BRgE83CwDbT1tvIu4I
CzdqugA5ZpqlTVdMtZKUVrbeKfh5DSZlzq8o1sbFuim9nBuVm6S7Oj3xAVQGbCvYFM5DFxeoYByG
QEBHJXce8N3RisHM2AVSIrJC3xJY3D+JsPlc6ANz53O6S9GNo8FMyGhPz/xuRkoY0h9hte0XH6cz
fWz/kOafNAtjYaat1lPQL08t2oOhA1nLm9iVJDLWEnpZA5zVOeOq7BDa/biDTNio2U7DvTPis4SQ
W22sVpfrp1i7s+ChCPmFQoaBajy4cZgyGkwN7owcY3oHnJ7Bfa30f4A+4Z76ZYvKe8a/Hh/761K8
SGlzfpMnDHW8n4AiLKScoZkoMReE9N35wobfIJpbsbePtXjUek4vfqZ5L8uNTZZ9fQVugovTG/9o
pgVCrEHM1wG7f/RPNpUha8XMa77pii6c3fIDqoorOVSjJXaVCyxQRsbWQb9Wqak0JQxn4XF5HXbx
m3jfk0MaMVuT+1FpjyXYnpWVXqHg8QBdcY5a1M7EG/hGtS5yg2f4wgV6KHTAQtNn6Wn3SRZN921D
ZfmLg2adGJU5kjpiX3KhQvGQfliF9kZa7mVVHyW0MyboXv1xfm913smxaFr2Zj5tVIQ5NR/VNSma
NfbqUWTi7U9ra8sB5e1twaHncEmL+qIis7Ukld4hatPDY9YxueNxjXclKsqaiQlQ5vV0dqVbUamD
EllkeF0ODDPK4gr+Yb21DM2cAPrd+kF8wz66lcQdmVLWKsBkPmPRXmeuwdvunSRz6ku6sohEdQLX
hsNUnwYvULkwZN9dNrDQwFaLLOxMy01Lg4dcdSRRAPJO5NMb7aVpImiDAQaN7lHF3uwYl/bsz9Ia
i+RW/SqIeShlZdnRgh5g4AZ6UzftdK+s+/hdyZuHFZgMXQdy3LGLAtfZ5yugjrwdyuaUK6v5uTBI
ucdklXZuDdHi4vuhsfhU65NBMLo/mBcxXEGx0meddQVXSGo+PoQfiUz4cWEGafHUebziD55pn+w+
Zg3LMzoGSshIPspQuq7NR8FsoNB81SxlwUq7z1ePEn8tAOITKwcxALjLSWh906P6MlH9rOJ3ZQjB
8us7cpPpHjgazyPAA9HV2UjhUVFRb1eoVU7TiO7LKwihc+TxRp9dzbsHTL/RivclRxgy2xWZopsJ
L4YZKyyzj6BdoaY9evcy+YwAUYdNJl4j4SAbfXUhtwqm5ymXzdUTiiPG3NAcYUVXLmnz8fhX+1El
gpaoDEiK2kCEw9FH6x8kG6gfU1fLOKpwdv2fYaZsXSTq3Q8RQaSEXcipSXwYKYWrq4zrMDTkmoxE
DKqNg0HDuBB4+nJZRzrw7hDqxamVrLuRhLGqCeleahFJX5x0l0cSlvKBfwq43XIKQHz05ESi8b7F
iK243FGQOY4+KcdLbnHQLDW3FxFymJU6UD4ewP4u/+2R/YU9SIWWtiMVNpa5SnFeCtYGMPzE1fJG
nrMH9wIySNwCAAvsXtUML8uMgsv4QqWYWF30ketyP2jyUhDv1H+sWGhOriuY6QP+peY5l6v4nCGY
RWx+GXlhKO0D5EOHgTCG9c1/IikuuHWzNAWwjnI1ySqP5ub6N6LqP5UN9BVJLp87ZwQK8jiNe//M
uJnKm59RDG+sHCiEu92sbzOm8eufV2IBfzXBKi2fFDo5Pmi89wzC9/CmyoLIuSsI0IjeYgpxYWuf
gHKpSQutHBBNwFP/XnJ8SNxydvoDYrXc5GRysDs4Tjhi1ZZlzS3yNABlPgDOFfiYUzZzTHQEGMjg
Fxv+UsH0qS+xIS54G1op3yUqUqp12f7yXxeNw86IUyhscD0dJQCu7+ViA3feDG65M4Nc2of3mp/0
gmuKeKTbVnhqzs/nNOyXC6jn8zJrL/jjWRzsFuMQS7+vMjS94Hk99xw4QXdeUxSUrZw0puaKEmcI
FxScbzO4uLWyVOBpRnbtjXZhDTFeYB/wYpHJqGgzYkiPZpP63Qi5jYDZuYm+0L3YrxsQ/eYTB3cB
lxs6JYBt3WDbwsxuRGxDTKZSyqtqJgSoxXkgLntmQAsFjHbJd4nZ1FritIJSulhxerUt7CHLuqOo
narZNeJvN3PsrZFD6mHJJ6dPOXQaSr4WWy/VDSpC2uc8wjZDPRR8bsjD/8bzA6UEGC7C+/f61SOR
5m/qvPVpByY5o5gTqxgtN3/gljrpXkSpZY7SU+xtdeGjV9A+2M1lF2TIeyBgM1yTvCxR/ltiQx/B
w9eJyLTE9UXqOW02XQrIIxzxf5iIAi/Sq7hkIykJFpIUMRGpLOwPh/blNZEj3nh7YIpWXgvbXc0e
N8O+8uYi9S6JytTaS/w5fkZ7/27hsdaSpD0gXFScnTprYjpACQM4lNRcTB2fKA3r1cKoSUquMi4Y
rWPo1hx1Pq8Xjmok8HYtw+BpcUUbiYYfnhUJgcBESmPhn3m/+UfU38rD5UKftHsKQfEczIzcpniw
UyGpdCdG2/eE78OTdPrM1Qpad6snUlhPZazyJFipGtPdIfntZ2fdUFEmk/QJ4oiCRBEziTl2xuZE
onimWt5MUMKCfMIeBXdYx5lF8TP5QvqVsYTgAnw2ZrAWU7LhMGYzv4sjU0Sj7P5DllC4y0SE+Puw
RflgYpPQb+LOUurZI/2iokGIOdN1nSLfvPh+0bh101f5PIgZkCNv95KOG+sBD4pbuJP6Ua2ymhl0
dbS+AMvO7XUbTmvlxk0yl2tiNazASftAq6cFkTRWvgOOWFWnyISCfatuxWsVY1Mnjp9W4matcnqK
ZGUioB95VMF9mz3Y03ErM4tvTtJFiZz1JhmdiHa+otFrRURO/UFs8BLy3NsyPUGzoBM/OXwwJQv4
lguSfAci3h05soTlbPs0i2UrLTf+SAfwKbxvnOsRTat5tBGS7sZgXUKxgUWrAqfmRP7HbLtZifA7
81NTR+tAskfVlpOqcExXVGB2HcGd7oGwpjE6F2GASCuYBiB2EaFmsuHSiH9/Bzz9mRre2kf3uxoU
PZXirCiSwTNzIXJZFw3tZKsiW3HRxHxCnxIi+Q3JJS4GZZ60hiG0lXAN2jExHhJ01ekNSyglgF/A
IMn6fDBn6g7hbKrKEF/4ONJsOCrm9cu3NwdfVa9Vh+agfR+KnAM1kseOjzX4vQN2n9DvDkJx8QdW
KaFE4Ft5bqwxn4Ql6hSfpBFIxNIE4eiCcQpVjC0+MF/apYlbxfbeuCrhmCjtiy0CbzQUYYLjtOTr
vzMh91uSpwyuM3OH1Q7L0XQjnIQ0ci8lKriPhyaM6Hw5DFJRT2cxigfGYQbS9i/7HFVm2wHW+qNZ
0yg7cMqQYxaKpTlTW9Teubt/IfpS3VezkRSiTLy/LJX+PivQU6aznb6TGd2xLStuyv7PIAyegbee
qQOIe1NffY3WickZiHbrsYlm7lq4dyet3H3bfY3D6dw/vpAs6LcqqSBttLF8yeNdbXVgtv1AiURU
tZewFdpOkL/U3F1B4Xqcy7w1qWlVP3QTy1r+3YDQ0OIkQfLskfUGZq9gzOGJd+zGBegmOZFl3lBQ
ld9eiEaQSJH6/b8fe6dx4IdCarq2AFEH4f4d86O3qi1kxrIxwUBV8K/bTNos5n+VYo/y+zrM676e
RYdwq+YYG0Cis3hyR4IS3rTk3vpcXANI2Wy/5RBtJVIxb7QGE+7ThdsnTKZS+rVgJtl65Sey+o1m
bg9Buetu5A1iekKjipZCJtymyB8FDYUOi9+AXyPnKWnugYsDNpbhFVKeOE4YXLilPd/IzJpmCSKc
Eigcd1FQ44nreEVTwxxr5ZgqUkL+OWrxDOLpgJ3uJGbnBXvkTvMheoMnOiqJ4zVHJQT9ht3v800q
Ok9rGdZ5wCY4ALoTh9xjWbxLm3zpMYojXF5HJQ8aN1/sqiLKylUuVpkqpBe8aZ7So5elq0IbcsDr
tSMEPhPx43lDAXO5U639GOvETfxodoGbgoh91ve5RzxJyictt5+lmWNNc9q/7y5QgdyuCfGZnENj
QHpmjLH1Tncoh18GG2csWXecbniBIDl83gN7n7Fey7twWAOF81NPCVCl4PqDdQ3i2sl4YlkOjJbs
6GJCZURLwhg04guc2op0VZGzFkmUhSCo+L1VY7a+p/DEH66K6PJS137gkYiykFXyLP0aC7UKNxKY
bQBxfdUFcqlIMiZgQIOsnBMBGgtpXsf6MtkJpWQA25lxeScEjAM1o6p7evKwjc2AUZ5qYEuibMQw
nK2sm+0uZtSCA4JflAhjT2rPUYDsQTACYm32svHriU+9R6sxIaDNNCSOrvoEC9LQVwyzWfn7b2zT
d2AI0+VMZknp2HQ8uWN8BLNga6wAJkiHCDaxHyy3kbsLsFdyKKyX5qx+inH2hdmH3XP91No2oZWA
WtKGkZq0KcYZ71XESU0HDdcciFgYCJY+/hhjTbiahIQPLcbPoY2x6+khH4gCu6A8CNl09zfuHm42
x63JF0DA/0X7C/Y94Q4Ioe/ZdyMXQyPaS3piN9tuG6tR5RUQIKnTBGHJ34Xee+DhR9xs2c0pYu6M
56+gTYoOVBWNXqOsQoalmV7CpeVHGKuYGlr7/fdhb9PScdQqDND//QvwLEAtOu7gmTbiTcvr8xme
dr1FItbciKpEj9Qdxi/E4yQw/r/Z007HU1Oa8K8c4quUQs29+saYgxbAeIzNxe/q/WBRdvUjBMnd
F+RswSzLqO8Cxj7ediVM/spZ+KcNJwwWLaJ+lyvabrA9wLGlyH8AmgLdPkeU96A2R/UbyBxmV0l2
/Tor5w2DLjbD+nFEDITJk7/lhW3JFipeEAlPDA5Fm9zvPWo4zXKqkf2oI6FV9H6xnyGjyv37up9c
3yqhlt50VtOozb2nFkiIGGcGpTC19qFLZhFL5Q5B3/KBJeN7Rd/8qteb+MS0wq47bG7577ewiArF
HgDgsxT3py75Wk7fspAUfkAnW7Np5zvsYTzyls28ua7trVnk/eZcrDEb7zx0fENCQuppAjwl+ZBs
x/8mCT/Quya/aZogKEmMJGTMFBPRK3ivKuffANHYPOJiZvsZQBpAAI+1jHLyg4jrFdlqEeKzNt8i
TuPF4+uCng+x1/BIKhaawBcs/nXvI/mQX8aVCG9WaTkDbrwnMiMGerUJUxQmgdC75rJ8i4OEHKRH
6vl+5lrwerRpHnG7fbzdPQ8TS7u7m7a720NT3JvdMuQWigKJvH6/P+yE2W1JQh6mqV+MUcATMjhi
MqHK6OLHCAzLIEBoUuNzsvIID+HAf/FHgmtrQbpWOes8q5F72ggIZL4VQKOoY/jw5nH7jpt9vFbS
MFElcqpm/FmnJBIqaV/c4PRNlspx7ykfVD+Zh1CJDRDUE4ooklGlKw4WgbW0SL7oAIdNdRNFwumB
0xXRY7FbvRqh8sW/XlboP/P+6bfZQk7vb3iZBzJ9iZD3SB0BGfM6AapRPQF5hxGUlez5ibDPjB/L
f+d9i7aKLYbWtkydPh1UHme58PZV1/rhSHekduf+H3Mrl30GDe95Jk1xIp7eyJ42fKptoXz7UGVM
PeGKzHhgF2Sh3XjPIlEqU3d2WeECkOWJVnPhHd3Kjvkc8JDYALULqFWAngHQIVz/C7CBrvTAZrQ6
/PrEz5SxD3JwqnRNEnvAgwnMAqa029nUEFpeE+TKM8G9bQKNUGy+9jv52Xt3fYM3FWysmiBMmD0+
WkNPWfn18URaNXfxwhXajUDE2/KOPlaGgA0kI2hhUoGVVbRVULWNI3cqvPYOC/dbF/Qxy8GeV5St
Oo0RPFkYM6390JsFl1K8L9e7BJnZZ599+nLTEH0wLlRoP4EZ5oZzxCrcnMGPbCkB9xIl9M/nvuZP
lT8y1XD6grmCYXHxDE/4A4F1PxSA6hZk3BFQaE8IYgLs67tEPdQfPVQ3g0wqJ+QlVFTi/LADe41g
iygoFWKuBL4UujBQWDErCM0K7u+J5hr9Rc+KlkfmY6MK8K3wB3Tk2ufZYBIPTvZqoz3LxZdGhh1L
3YlxtRgh2e/bdNzQHeHp6DFVoNDWWyjPS1zAzwY9kx1eeRsRycHW1MSgklQtaotKv+eGpuN+PkA3
RA82/eKpA2PO2cC5LfrvexemPd32op1XJGjiSbtLtBwb4jekmJTQ4M5v6ycT3EkQQeOur99PLDl/
zZsDYda0fT6VAZy5tBX8FkNWbiZs7XjbIdizUW4ab+ljVbeGkWTeAq8Qd2tnq4P3uwMBvkfEl8vr
uYBdSzejL/w/lLdkDXTYE0f4RdOcN14c9bx4/SiI93+d2Op5oCK6pv3hoBGBFYFWFW0xKIEaJ437
Yi/U9pqfLNihuNHojpfjFJrcpR6/CeKuu0eU4hG8YVlI96tRqJlWWYbLPuSJ4xCslrlmsgmgOKzx
4sPl5Lw3U1gKPUCpfcCt0sK31SARISh12SRu2cnGe/go+ZpIFpMXYqCZi94t8QjaIs+r1+lXsb1p
XZf5L+K7VSEXbd5ifL2ShkXIbRAq0DBoAxXLSU+WIBLdFv0+hfIwWHJiy1LKwsPkJSi/B58Brpul
1OF60uGa/oVVgaYx6wRMxT6kK0TkSNtIHUG7z3/o3LcwXoOr6QYqdQqQGHcdmg1ZfLDU3JXvNx8l
ftQZsP4GrtIjrjc/RXNvP7fmizI6zgbSaQ911j2EEw+gf818M8okrZE8rotldBKsKlPqQ+i6mJ79
JHPqxVskSnzoPRYz90vVo/9JSjO3cZDJaYPBZHsYKynXITYPmIu+TVyAisfmB1c6YEkNBvcqigtq
EvMJm22V7oPUlDGKEqsyM+gpueKskLBAULsoWLdgIG/pFr54sNp301/EyIhw5WOUitwdDzQg5qDp
mm59zdap2gwgIq6zacL05KFJXyWPalKVTfZD6BO53Lho5269eBKRM3yrd5ViZ+ant9CaLNPrj+An
aEgOmZin/mbAFG9oq7v0UDu9mVAYNygQ7JLLg/RROKjzsAtIONDufaw/ICjqop7anjiYZsWHOAKT
HvcP+K5TRnndI4quKkU5bSnVYmdXUlvtYJy6KX08Yqyc2xyyE3/7VYorVUpuzaRnxbNhVI5wGRVK
IC6nb2T9SXo9+ZnQux6XSyrcplQVlgooCshxPo8hQ5wXRRt5DTCCBPQ2ml2asrpDmrzxx6yg3Why
TApQ0nsQVN4lfo8fA9UuU9a/i+s/pyDAC0OIVRzD6REDXgLt9mJgW78dXasJ+cSQKryuAWUjvYv7
f1BpsDklYnKebSQ2Uet1BtBOrKMysqF+4z5AxWjWpv6nzOFRrykKRJf2dV/1Z4HZpBAZnLBV+SE+
8h2xXL9oFFya6T52GYOWCYmEhSBk7nGFFW58Ch7I08wAyPCrtaIaoBNs0H4bZ6dCM1qinUciT+vt
7daWSIvWdfBDHjhfO15K5ovdxjQJcRRSwhWUJHxlCe56Xv6nIAZKdbjOtCNAP6K4ao6Fy9EoQey+
+pIt11uSQ6v7+cBy4ajdLaMXey8uOlyobTmwKxCytY3tOor3+yUQvYEjsSAx0F/H2MEHuIILZaRp
n9ZBGE3Mxc2o7vUR4OeJZI2mFLXfMS43QhmjDkAsReBz2wW/ue+3Fm/ZgjH2uHuBMtfBAte45Yf2
sYY8IxF0IJt7D/J77hQuY2PRqnUIj4rZig//f4qFUQRDhywFPwDx5ICBqCPXSBHJm8ao8Bojx8Zb
c5PSX0e0cBwdKkm8GBdlmXvi+TRe3O7A02AmHMbuVoOt5v/sizrXLzOuHTGe9IN1Kyr7N3yIt7Ch
AWXMMwmX/uw/5LaVvj3tVYjPHusluijR0PEb9RE4OkAC6W92X5GUZKqtz2OrFFaz1XK8w6xeTXny
Ucz/o7frK6R/nmH4vKh6OR8ZwPXlzcYb33Bbq2i/VZWiHMVIWK7Uvyd948U9MRe6ip7Vu+WYKIwx
kYSlwJ066LRpHu24nucVI8xkKqArQ/vUT9hLLW7JeWWg7FfBxzFwWUrr/ZmcYiqX92PWnl7DJbUO
UXLOIK6O/YpsXj9m5Gpeyf31daL7yCKfprDzfPcmUvYtWdJlz18ku0yL4s/tHhU+R3N5RXPlw+cB
9rckiaBcmgSmoVQcmDeO6aAYCcBae3FSqaY+qaHWu6+sGviS6ODZgDX6HftNNXGAI5fOPSg2742T
Qx5LGRTXgBYa9HzDRwFhOE+Q+N3b24TtcvbmU5qpD6IrOXTQwB653v9nZbxpda+G265PRkSAbqWg
JvzZlgcloy70uUmWJX+NA+xpuj8dDlqIJyKXthAPUPvPBKvW3fXWj0ik7qcy9Y/St+TnpFQYA3hE
qwAEATQoPAu52oc/1wvX1SryPSRugZ6Nrv+0gvqjIxiCV+afDLNQBLFAjOwwWGAw7Hpcn84ZoT/9
9qNlVs+SZT7vSurgJxV7phLPBQ7whhPJEqv7KCm3kFqXiy3pnHjXgZCMoO6rAMsACjSE8uHmGpaC
KDTVSy6aaLfC3W2J2tkEnRqHf6Lmji1f5JGBikxK58qKnw4YAhsTCsuj6EAx+p6VNohYkC0mubii
aIqKAZ0R1zLwfGtvK6ueZrOaymMjZMYdYabwCBJgcbVcfbMeuxkWavZUmUduL/iTqzTmL4jTMMRx
Z3qvymeHGMJUBaMJK+S0lcmoS9Mb73Vn/N4qsOtP6delucJ8/L4uWcX+Wn5GjT+3Wtqo1McuNbTJ
e/58sEBzDZRUiGerUmiybJ1bLjJYLouY4nEEsBG8rsdp5Z2bnjt5JYAqnuXjgg8NQcEuq2GPuVix
cvGr8CZ5n1R9ElF5wEU1ONUajhTaIijqa0FG/aEAYn5bH7dAlMt40DBfIhV79ACh96NcuHOlSqG3
mdXQA1nhjlzITl0Tnytb1xxV1anlI9xU+WBxYUno2uipO4beMAVxJgGW7Mw2ufjisUmExYliUni7
+GouTihyIQIg3/+LXReu/tA4lZc+qaZOygiyIn49a6MewfvwvdmtPhBPoacbLqOiBRdqZWo9lgEY
SYERAmRUgBr/hGEzTveo34CMKE/xdJlmNAySTB/d30Lu4s4oYnJagfnVLeEg06KPCyCJCoOsk94i
HtnhFFMiMKLEwgmsyD6J/dFYdZW17Ucn/prnt8Q3imUXruEsHEWPS+E+82q3oVE7PHym3XPTG3tX
2Xf+duXpY4o6crevHLYnCwGFmUYLEsn3YY/jxzSaT48fjHRd9ThY2meKZHCrMFUn7YoGrkwxNvmA
vdntWgm3vfSapiAL1cPp2p02dqq5s2/f8WWA6UlQw8Mcd8kNJfwrlYvfuWVPwaRZG2uv86lyZBV4
573OEcf5is1JBBvWW+pewh40MA0CuMI71Ji0jH5+9LP/kQaJ4XnldEFm2dXatUlaKnEDo69+ZCet
syrGa1jSLZWsLvDPEwP/EwrM12aMb6PAWfm5WyutuVy4j0s0sIZDYlX+5X5glQdg4SjdbbRa4qk7
ulxQmu6I8o61umCgQhyg2JemW92eVRis9ZcnC3v+LIUfsv5/PDyfTYiB62utxgMH3ZhDHfUFISew
KZBnt2vfuUtQcdFlJiY/mRoDPT5ZBw1Bkyx6D0RN5dHSkrc3JByqB64xDtuiU+3O+7IVECiv3e57
ZwE+b/BKVXB/5Hxq6+Htj02rjnla206NONhF31jSybQs1ae2GX7zaU0IxmVEAlqVarJFS9QTkNOI
Br8m4wrneUYDDsOGs4CWfLnwkUxPDHDP4UURyrucOjF40NQftPCkZs6+Yv4dl2yn2wXblFTBZR1h
NcdssJXCOOhyjlPvRiEEZgsSd4+htlx4wifqNpV4Sp7nOCS9iaifg9PekmPSB82qWfkjHwhzEtsg
JQQVRHMCh8GajeHW+R4VLuQW0Ixl2dVRjym7LW67MZGOpyCQ2tKab2rFkacWAajfeab7m3NXelj9
BnG7TB6RuZnzidxhTeTrOHs96KQIOuY5s8ZGvduhNmZ0HKCyx/q+D4xHeBzc8RCIuBQPrsgliO7Y
PSlXpS8iTMSHN1Wr+kH2F25E2opPTZhRSJJMQ6BHhXlaGo0nqwm5ZWTh4NHD6zyEpQm7B6lQ6YMj
2nlVpoTVKuS/rIgK4ICbYJSjKe4Mn+uUWLyCMegJotvtXNgVLxibkR6NQbl/cgA7su8lKvw21U1/
duWEhNYza0cQAqFd1JHZduXMsX5oHEFd6Z3XEV9s3QMQ5RCciBTJaCU9NJZFX5pUCZCsxgxL6WZE
jUwAYCJ9LHbSFogCOUaXnHPzx5BxVvSlFEKU5Kc/9eCmyCRm++KhOkzuOR44Cap8tGd0cuTKidsW
ZJRTT9rHMn6hX5FuO9zjQqP6DfuIc40/uxX5g6af4RQenvdVI3LXuSDYmH+xajBpa9TkQDaUWI7k
WGZN7e9IUdb0MoEfpJNUpsW5TxyyoOO6iGMn4mM8uVmQHPknSK49QZs43vvZLJ7VfELsTOeQkmAG
gdF+SkWLr9FlBTY7fXwWuofcE/rRIigRUkSDAD5E5sVLAhm33AyouWIM3vRe4gE3MAEnvRoNqWOq
uC/SkYQvJi4/0Uwgam8+URNQd6QwJgGK8CyaaS5WoDrHZbztIhqGkxbewyUnhDvSoDphkbvMiG16
wFUTe5DDzcJiw8bR0HsuC8UYYNkXmmdKPjdcZxKga/HGQsliCA/czNLCK0wxpj7HJDcRNTTyxD0I
a2vvbIGBoxxvKfFvFMiGg+E0y8MRAj2BaXDQkZmzfo3qu2EEKEC0jPzYyV4c/S/nDjjRehRKhkC5
5HCJx48IfIhh0meVqoyXAbu51K1RQWlHBi4ujZ3JaCVSg3s9ks4mt13Dx7Lh4ihnN5XtEaneNbmt
kMPMgVfvvHHag+JEQGLhmxvYdrj7A0yNYNyPVI1W47cBnBYBt4gGqRisydiCvr0G08+hjVKCoZUj
MWm5d2Rmf1XxkVBijWvR1jKqDAzuUu/HgTODQcOp7HnYo7HtrjaEJ2ErXwifajA3T3LN7P+CSPdQ
xLjIMQdxxPdZufri1C2bi3DjfRz4QqVW+wjQ4XPN6KER8syhV5OvJY5gIB+XzF/9t3QmjTyAem7I
xiCxGssA/UM9XlKi2q2nfAWQv1sQzWL3ZdR3OJlCRmn0+biynmjpVKXqn5G0hG62966E/Nhx8xO3
umUgZaiJKQlVDBhrDWNqN4BQBlvTkVifwlgr6fzLS+QPD3kGb9kOe/9AlxxSEFrZiOhGeOZY6aiu
5ahM5LSZ/wTZ87g4BKFHqO6CDOv5W7R4D2fV13tNV0wMHgt4FBbz5fXrTRaTi3TcxwA8/nJC8lLD
rdNjIMFsSyO4vmAMQ3/Sdi8FM2yatJTPU5tM5g+Sh4PZnFu5Y7z+4yNit78DvZCluN9vKNpiuy0T
U2Tp8zG6xA8LPeBPvBhqlT/u0lipAjyrCzMyB3UJjJDYH0zzH9qSgg5gMAi68d3GUr+BzoBVW+5p
vpweoca6u6DyXmNQJuFrzEOfS12NcxGaV8RKZsD37nKbRZRPgi2+mAxdt7Ojdt2Ij/BfI9d1b/gs
jfx/FF0zbI/RqOEp/yRYQHmKIU636XzT7ZKmXFmA0qlrFe7GKHmeexYXzOkXFV9UJ3kEq3gM60jp
AwF1iv8377w1fQLGJVQbfXym5WeCI/rSyfudkoQFTndB9GPupQ62aVcNGILquxM5liaq9qq3sOIc
rax2ObENwm+TRmnaXrYw8FHeDrVWmQjw71t9j71GPR9p5ycLo6x9B9hlsJzniWyHvmds4+oZ2hAO
gZUnrZhNsS+s4rScOEGIY7FJqR/ahmHSyRURF5sX7pXEUp1Dza67tmkwvnMJSGM4RzNaoqbl4eEf
Cd4yyGjV+qdapp0c6BpCiLGzuPGmjhMKgjLNsahEJ7ut5agbucH7NPs3y69MPAHGEfqohCOyNU21
YaBKRxyAxxG3lE4JoxfFGwZB2SqNIgKcrhliTi9dcJEcaHYa8u5HZ+TCKccZJJHS/8wcB2aLhfe+
Cq6EkuXDQReoPK7vWDprINL9hG0ZdHFsAB1LzI5OAMS1yHYKyhsCI0WoNNsaUh9+93s24mIzBPRM
cWz991mL4CmjGDjeg6AgUN5kPjctS9c3HGmHP8q2WNagdsrK25JM7dV5sXcoGBh+pT9mapgtHJKd
FEXxT5S7oYKNL1JLsQU9N73GdJofD80uiioXwe5BK/mMUyId6eCxyBX0ULKLFejecZjSntvR6Tt0
P35D9HHVKao2BYAVGtGu20rE2NGwZsS5qDVXvbTO+roERlS8PVFiaE6htffzt6ljCb8RI0gH9grt
W0+apS4i9KZ+GEEVYNjhBRNjBCFM4sZu84i/jHms2f3YGJTqSfpY5IVETLrRph8V8Eq38FPa/quQ
DIZua7hVq2ONgezFRARpKLSoHa1Jkki73y2tGm1BWLLxPSQ4JzfDlsdqes6Jj7Ba6PUlxLKqQ05n
nLQS38TIRAxJ1S4R4fN820Dy10vds+qjZbn+ERAv2kJqNpDaIxnBUOGisaQtcV9hiFlC+/osT4Jo
pxIeZl8zei4okLwDsC/t5slTEg2pCdvNz6ef61vmyDSysYoDPyiyWJP44T8oMKkceYjKyoePH0rg
aEkgRn1xVf6jBzywtyG2gPFKDZ2/kg1JwQGPR5S2hlUrbDDQtFzcUiP76476Iln9HmamsfciLUu6
f/AqyV+kumaelRdr8/dVHfXz0W78XkX7DlYiAHUPejfodhsDTIeuUjHrW4EvC4PxzORHrkIu49Hj
p5Lj+pNvPoNR8pPQ/gMf3H/UOyqtxyNEf4DaSMStWWZTVswB8l6yxmxrdAkfSRJjRqFt4x4oxv+W
HD0YNa1CJSuH+o0xx8uvo7XzE4fhUC/k0L1/SzksGTAG1GKei4uI3hmwc0o/bimJ7V2TipsdC3iX
TwctzSRF1JarnGiwGQgRzUPQvEAN73wSt6ll5PysQhh1XRI76o2N9fmZC9msgGX43KszD3QLXkiv
Dle1fJDMZuukvTnbwkW/khaQMMAJbjJOjJJZUYPYG2XTJhvA2TuCZXR7DXjvR8PkGHLvr1sxUFPh
aZW1u4LQLB188KwO0hjDkcqkMy3vkprQ4KetLt0TACeelCXtOz4ZvF+84BitMWTGTjRcDHmQnima
sXP1iVuuhjMUUa+nWWhVYDFeUwEqUaq8lGbFZ1B7Kyz2d/MGnM/lXV5xlB9quS8M5EpgpyVieFTM
vkOea28B1rQXEAMTMn7UDmwJUC4qi8Ws1ecu2U+XzxuUnKcDGBO+fTZF02ctFne3c5vOkILQCXRH
5H4v6AK0WtJ7fZ9q7AXwSz3bHIR3WS9gw6qFqk6eUvR7VNfJrw0r1DIDfaMoPvLO9VrLL1608xM3
aQnQGl/T51VtiewpfLgmi3GhH8uax18vmPQosL57YUIzdS1q0zCBmV4e2iVulL9tNMRaiKW5qofA
4Bjc3S47oPoVUBIC++b5JClhIkDFDTllhiCA9bui0VWD8XKEF7yu6jwApDpCcIiZVJX9eH8vM0HO
JqLPi340t74ldhK+nS6yPoe8Fx/GDNuhzFN/esYQ2NCpwv6eM9Tp8PlRBAtMiUmHrGWxhIo6NPwW
VpP3Z/JSuJct93gbu5E2YpnBk/+1r2Sa1HuhVaP8Rsfd2IDPh41pDj+9NIdE5mRHcoCoFe/v57C2
nwRzbCkXRWIpkVLwtCstDTBCj/EdW3Xivw1aPr6Fe2EDr3paroybcOLmJ7wEEskq55e7g1iwNQbJ
TcZxAjRwKrr44lNg38PEFXJ+A6aFqtUJAVcuIOuUYhbHSeFVGqvQLHOrJ4zzbOWDtw0Bn/ybeK9m
YylQHyveKWmWboGG/VBzOp/xZLO/NTMQPWogcdTFC9lm9VmwhglLbnuw1A/TnKLUnol5A7AqGOM0
TnFkXnFPslAzGI2+LVciULjSCf3/gPRZv2HjRMMWgmjWVYw1S23jdwF1c5qKQDdde8wI9f/c2Ecy
4BRqhgfXuZEDKhL/DTOJ7oVozZKq9USuiYzHpSvbpAn45xyINhfVa/bKUPJW/Pn3gVHKS5EzjMwb
rgLCsxWBsTY6ZUyp/jGquwKAZ2Dq7bxlejwt51YBfW+60Ru289t53xZigZe7rpr+x5JP6jukzM6v
oopss6zW6ZHTTXuC88injkIWjAFRz2F8DKSgjal8EduAhSw0ki3CfSbUrxoVewYSU2RUbo5X0ExE
0z1H4pTZLhPekxI/qEmaZSkKyAB7L3nOqKl8+2momsG8TFWA7drcNa+Pt65GU7p2hiuGZNx7FoPs
71mT/dXROYtwhGtX9eWZcDach16q+vtQrZTgerq5UqXTi9pKQNZXCd4bkv8ws9bQq8CF0h7oxJ1q
mEJFD+A+FucKXGSVrjh6VS9ArF7w7yptTBbLp7+uzrawUkfSPJCQvgewn/GlIJt9VeFl47y73c9G
2bZCHsjVC++dc01aN3MhCaK0i6qadfgEiqmrPjSOnmjUG3CfEi0DyQyjXi0mpLy8YcWjCAMK0sm0
LpzHTuWD9ExdmzvQ5KY1I4uBC8NnJLO2Bfb8NxZmj5EiiR6mE03nF81h09WiRywBnj5qSsa2J/vc
Ce11/1QimqlyuJ6ETtGW+sAxHIIcV0A6aOgFC7djt7Hzy6CdqJOqK58TLbvvbZ0MJJIdOBQmny+J
pVZQk1ohOGuDqSOLryG0zn1KAhrSHTZEyZWowz9mu9P+xEyFC8bAPQ7IxeJcCMIV5Vg9GpH7yEFD
TK8foa5eq7Q89R+iamOea2ia+dR5MoutzCQLbDAqlRfwT2LAn8jHH0SxGTpsAGm1vxbk11Q9Sfi6
spHq7A2JeKo34kE/DDZ3nd2Sq8dXGviS5vqG9RkadmFjsyt4zfjOS1SgY9hEVKhbeBFVF7Qg6Z6f
55qVJKG6OnoIXWGVgqjVbhT4EP3K6s/RLNcsl/8OEhSXb1GUi35K6jtOgsBmuYqNLto3nJ8bS3S9
W+86UiyjrhXxmW5ADKvcNVdkbCHCGMfTFOPJXotaLvk1V2rQBsgyG7Auk5awDsMKJYs+jYOFomoQ
Ew1RlyY0fxTyHwGWA4LPM7rxxdQDNgK93NZqeUApIq0trk7moG6cY2R52ACmC16zPKL+dHQurTqN
AP/wK3HPdM1J1Avpw1MYU0BwFxkhr4+saS/h3qdISguhjTMY7NiJHmN0fmCX8PnFuTCBU4vRJ1Go
O6k0jnqVpXiQIweNyL6mYpKphKTlI6r2ze3f1j8BR9AWiBChNa1D3qRFCM6FZFB1R1KSOQTHsOh1
FkW/2mdvCdkVLhff2PQKoG9kNtvdnWlT1lIsvOZyomiUcDgKt3N3CMpjfL3YNeYFbeEvwej3RcOW
k0DWjYFLIpEZ79fmYrv5+Kp0OeHvvPpcdSqJBZLpXPEtv3CmCIPnSUVUIBEHTPEm5Vz0CZsIT0oB
pLTUrzCWk8z3Hz0PUdslwov8rIJPseKu5MYjJb9h0SjLwMEwTKX+m9hd/EynJsVZJizsDz8Kexm/
QONBnZOAdcjlOXOuWzVjHxGwr9k5N9o5SbCFMWHwx2ScHs2y5NLqaVxb+EqEyo16fqwCmgeAvmPI
efAkDFO26ymrYgVJzaXfRzFjGMHDBHEOhPcD2L8VtQu3N7RwMaUqHo98c+gzpJQezzndBUmSQdfl
aJcl46KditZD8IPY/x8PKHeLzhC6WO+YnUYH6EGewaGv6OToUCwyVaIvOhtZvGj1zL9bMmUBqPxq
uEON6UIgq6+fmt8Me7jZiHsD74EU+Fp33h7UI2vQSHotu27uHShqC4O8IoUHbyh8vSrzE0fzVtIh
1+ZuH7HiCXx0prnoGqYKI/rldI0d7phQE+tpNeMisobVMXDZEXE3j+RAVcniAn0Qt5G1686A4lD1
WXBcUY+IdDgXqg///uM1LqvpGDxv+jPSSpnTCHA9fknOlR5n6vv+gGwU2kpu4RJSkThWHzi9AYpp
YAVhD5KgPj98AN4xSIG2mCIdbDYtE+8AvbXM+m+yY/TdC6FYByHCFYKby1vAdJWgjbYo22zxM6Ge
Oj8gbwf5tMzrYWE2h7XQ0rSIIsiL8G2hyq/SgHRtZy/9YPhgTewI0NLYJVTX/FCxDXATVxUKE/RH
1kIq5Xz8tsAINfeoTROGWkghlgwCKr7QlqGMLOVsB9B/0EGMhBdXz0mGd0mQEcpa2T8aekyMA4ZW
lKAhvvOKeuVQTTtGEwpwHq6o9DEKO+2qAh1aSgf+/obspsmcO9fY5XSY7ysrX4SLxttxsqZjV4LM
zXbK6Zm1Q+jxSzQ10Def3GmbZvHDdyD290YH0/0WAgNx0tZ6865rtkUAdX6x/nHGBYScjwA0javP
E17FJK59glcOMBziW/NSSWND3ZlfLtVPI1yyDJ3/PT5dI6GQO7W5zohIdsbdrwLQe/pbKPawGrCF
fFIJIty0ocX852R8xybJUZCfi8Sck4OFNYrAlqP+mvgsqrSH5l5435pzqiQYiPbbjXMeTg+1sA/w
KG4rP+oiF/YZJeGoKCFvG9O5yBabA/WQRZ5boFp0+BFJvQBIuldYm7YB4F4vhlTfpxFWlNBJgaio
Y/vwhEoUmDyTJfyiMelhzhd+bPqwZp53z4/5M+fACwNFVTk91zLPSiuAeeRM3nk8+nWgVRYIybRg
1EzFFFqWS7Im6zvW0Z6sC6n8VM8yHWuE/8PN4Cs+9z/+zxD6oqZFn6lVrRFdC+SuWaqNKJqXT6rt
ayiIebWptUP9HYgPW56vwpJogLp5HKNraD8fsa85Rt/FoXubO8gkvGabqb1ybt6m/boE5znklUhv
QYL+ZN227ssMT7OmxbaQlxTh4cjZ9O/oShc2R+AAQMbiVUcjd/n70GGU0tt83TquKFRwplKZx03J
T22xmiA3/0UBBWmCIqapq8Zu1q/tditp7PWnSb+EEFOLx4qvKirN0FwNm+iBYi/4l7Yhmhi1k2DB
PFaQENZN2Iqige8o2le+HShZuRrqvw2JbJmQ3LSt+OWy+q39yn4MEjWyVYaRiRkbQg54XCwH68kF
gRs0ikniFt/1UY4ikEuQEI2Ss1P2YdNWUn4zQEriIvte1jHNqsSGXB1n8rTNLRY2lVAM7jMLv/An
AQLEhIB/gIaXfo4/+ORZ/J3qcvFD39Q24FqeAHJdEMzdMetykHA7L+Y84S9iHnPZKXCQEnFS5fwQ
tWXoGCFAZwwrbeKaJIuRIa7BsQFQIPoheX2yuYrfAE7k05LU33oHBsVjXgLZBWlJu1ogAPg0Adv0
lo5mYjG1Focfa0wnqXH/HoHR+l4A/6lchwxaOBtJS7WNHvl5SwM0gQB6D/QSj43uGO2TisNvlBaQ
Eb70W4/vzCLJQwygK89GzSUFAfk5hkOUL8Z+h/2tjAwP8DAzBYyCEZHUhn/uQ1LhHS4kpNY419ss
5nxzDzx3bz2G9/q9D5yFb5DzkSjnPTwcJmlMYch7WoNsrbAVtf7Q4Q7KGLWQAw4xrBedg8jgYU5q
P2cak8Fz2TsxAKjbXCkWbs4ThMJWQaz7oa0Jwz+Oic2ePRYRK3LW0aNVwFlDAMhnXk4RILGkam7H
mhc0OUWjq0VifIuC5TkuX9pNQs7Jo1Y/U5VBTOgti7KwFgq1tKA0SsmOH/dZ7wBkGB6EAC+OF7cm
H1y/r8UzifWO4AZCwfGLIbm/jn1HYpoNY9TAOx+ZSqZApXN7yA2BAzEqVs8AaoffiImn6ivvqLku
KmK4bbkZpoPkIYfnfU3/zfiwilBY0gVJSnjH8sO5msuc9/BHaKW87YEGpwIdlZ/uvoLkENu2yIjZ
VehB2O9/k4qR+GpeOy8Wh+hf6BTsMWE290po3IIskwiTBBYkExtjfOXCuHPfOC93RzubDG3oe3AH
CQ7Tx1Tzi0mKdkccn85Vl4kYaDkvdFknTqw6su7p/9yI4pvUM5d2FT/cEt1HUWuGtJ4fSDLT0A5u
lZPcLQtHCWoEHIvr9fVhJXqul5+wjAZqE+To0nktRGxwvC1/4MHEnn07fPV4A4W2qx6MA4fJu7yc
SlXIDgxgq8+m0+ZDpv0/gvWCRZu5Pj4w3TF082/xJMLNVFql9rZWY/mz8lmc6wfg+wRTsrOoHX8q
EmEeq9FOggQFJ1qS1IakVwiGSaKbUURaxANpCkQO8q8a0AuRDT1NVF6TsM6Ie1zRYDD6KMa9Xony
ta4cM/qAV8JbYEs3rlm0XAiReGJ9dK7FPBAadNjhxTqDbXTt9p6F8hzYtX207nbijySXcsUtNQJC
y9c9zvaJ/sn3iFGVP+1XiX7Hbqrnn+YRg/keOwLBfhq/88tYXZdJ6KcWRk854Jh4BgneLXKwWR63
NK6fQ+yWcYjX/r1EOmuasTeNAYvYBWf4utsGADdn4jKkTbGimn5kVhMi0VC0d+R/uvqk/riHszSF
UaQ7K+XDmf6nqtK8xoqAkswRGRsFcL+7NoGa0lq8akej7Srr6bV+PdepjUvnXpUQMqpnh+fhA8on
e4USCJaLAHTYsSb7Mv4z1p4RLDjaWyCFe3vdJKmqFH9liwp1OGJdPaMkmsmt1FFJY+3m2P6+UAqT
lLeACezI4pN+6wcN1MFQijAMr+XdZvUn0krIiT20IC7PeY4jeIkwlPGEUS3sdl6ifYpKu92Dl0yl
gZ5yKXpL0qg2lgaEv87XpYLPOP6z932iKaqmehwbeOmGdHeiYTSWUFpjIdYsvSpU1vHd1FPzt273
WxZiNrtIG2kr01YBjlg5qI5KSt+Lbe+qYbxtoKvUswTKi+gdyICHbYtEW9dYOP+auXHAKQ6TYgaC
yiKMfKT6vUc4BhzWrHp8tHnmuJvZIuljrtHpYuXgdToNXfDAc0TD+yoqBLIfWiMZr0JZypOkWy2K
b0ZwZwwzHnvju8h0ThdAnLhCrGtT7TO7Zxig5S0pASsd4i2QGcJTrrt1KsNGahvAxjAGzGZjcOFQ
XU39yJMp+TXXL6xr9sraiK2bs+aNBLQToR3lCc3WkPUGIf1O4joDGsK+i7YHFqXMnemDjLwz/OdH
OrC8IZ9inb+dJ+YAQCQQo2NTo7reERvcdCEBsowftc64HsNrYbjJWCdjBjc6kONvuE4hR6Hyzknq
RfeCgURRZj9lPmhF0UQNbL/pJxLyLgtBWF6XOEsf0YXb9BEgNvMuh4NUQTrn/mVPyUjaxv6yrwxS
VMVhz7pyuErZDrehGU7chVQWCvHXwvmc2fzO/NDJROv7PKH0kSBKu96Mmzsn+L9eI6EK7+8gTw61
kDWFbFJbhhcMuc6kAA48xU2GIMI4UivgDNlA1O67wsO0h+tKVE0vDsfUfPIxKKG8B9BoxBEeXj+4
3LrM91ioaqf7uN5QWxqVVMZ+JJ8bsrsYyPml7qilw3bI5RvALnd7Dduf1oVAlXUgVsxL67u6YNH+
W4sIlxA1tNoGGRDkwzv4ikLoQBsXx72IfbVhvleA+f8GHTn53tHtYSey0mhUikuayeGNTyo8t7PV
1Zv3ANZ5B5j9D1dGD8wM0bYcw7xV8uapeEEvIvhoRihykGjS23tUzs6XN/CNm3Nlj5NhyTFb4bxc
D/HJonaRJqihXS+FYwRsY+dGbntSOj2tCsS1K8hDvpXUXs5F0TZEuWmusaifmVVPvZEQvU3vemMq
pZyYpLJAWTZIAp+MqV4CNiXVFvNPlnY7drgh1jmDzTBp5M8bfFNPkI0Ryh34PV/rEG2YxtEDDokH
eYYvGP19K9M719FSt6xDJyDYNUcwnmiWG7MiWuKAnyDhVYddxVErXojVW1I2j7o76yXyRlFHtf4f
9PPjtdGQggStnRslGyplFA2TyTAbUDx46AkVhJb0jEf9eh02lHrA5SuZwh5P8p+KSB/piN9j1bca
rrOj9mLvx0sWSG4fl/SGrDGOhR6gWw9jJEMmpt6Ih3NKs+0QpiA9xiI4WD4xTZqJQCDTCuWaEHF9
dKSwHkLJOFX8hU7YzybvFZeyjyySWnaxpH6xVVIlCijv1yXMiLwv/CoAJ6s39eBLU8r081GRAtn1
fz29SfkfXx9Cw56MKE68br5/Xa9UpUtLBXfI7u0wsHZnDqJdaheOUmPG2PLAdcKK3Dbfit5QDksk
zEzn0gid7hf1lv6fFGYxzv97o1PkrA5cb4Y8LbjqJ9aKasA0B5RyGkADRWJGL8jPgX2eIKHnwOIe
EPOPx9ZqWolY6Fp18sEJA88GbWYoa4SqgRN7EH8CzVdKej1GXtK9PjXZZFOaqhycIjmLZpIUUnzS
II8FKwCu0XVBhGg9XVUcg/u1Uklm4Gb5G+uyaC02OyxQoEHNPwdsHWXTQKgRe3PVIQ6JFBvjQfVI
Prn8H6/lvKHMS1mGm40/c43w5RkdRy7+zZCFqQ/RYMEc+HieETKid3RRJapxZy6CPq6l0dRRAAwf
aq5+OOdAmUhkgsUO965iKVEm9sI8VruUyUGXO1I7gwFcfKs8okzKit7+A6XQsu48iDyBOWDwRqfb
MDuzLLLueHa5UUOS0aEDsZ2nUSA5fCTQ4S3aHVWjeS1IsoHm8yN/+tl4csSlEleMshR4bSf86kDg
QIEwKtUFCzgPq+wtYPsFdhJuOf7yjpfhIHltvjdyKUoXLdCNM3h5krsRHbrYqH4T20EOaieq2Y2m
Bm0jM50PCB+FHEZGiWq0TGuhBx9YikvyChchJcA8eDhkuZ7FDjXpq2RGvBu4S0ExAQK33OSic5+C
Tnf9nT+6XgkgrsnNX80WIZnTlSaQR3yP3LFeMSCS46dqD0M8RXPvjtcNrrxDkAwoqO58jQY7hgdf
BtNyFlboAHUGfLMyMFRKIrEFg3hIJxeRvpgwWEbiQWdz4j9kQnAV97Zl8EFO5Mh9dKdwvzwqT4cE
Tdv0SPnulhcdlrhHOBLSnXRz8rBuf7jmNDk3ZqUjYPJfbbhoRVQ00beaAMM0MSNar6Uo4Av6lLpz
n3fp+AIqau9zi4GRMO+GrduGnVbp1N9p4V1xDB4q2k7CS/T5JLffsfF8+sKwPZB+oILSiWJWZovg
7WxPflsumWPrSfVHp7YIlzVcoOVGlDXL6UtQ9FwtKjrEYrRW0lEFgFRi7uv7p/BA+bV8S2AXOhmv
PpBf667yGim2dqDY08KJWF4CN6ayKW5rp03vuU+vbG5GnD6XAneakYfoNxqHiV3M/FGuyMaod4R/
nhC5tnovc0ZK8CMRt/jQZK0cEgG7EpqJTgGUaOX1LvaewJ5z0uojWNHjMa/GLbs7TlGw9sXrqkJ9
kvLPlKxf8BVAP8hD9A2fP+kjSZbQnMG1V5xqCTbSojLdC8PQtBhIsB6CDwh0X5H56uMd8sJxWkVA
2l6lGE9KtO0qUTwY0tmWeJCBPfMM+eTzosG+WD+7+bJIf/G4vRQBOXlTE58Jy7l8NVk1ULUuqm+3
Cm2TLatOoASYxjBsLrCNZP/8u2k0X+cz5e0Mt3L7P3VXBP3OkaVI27coHllXA5jlNd0LfOIBna8c
2lF0fGVj7iKxb4buwxSVepyRRktcqPBNmBwpVUhoTVqmwarmVQfBZk7kplbFT4RA5wDZjVTZlA//
yh1y41x0NZydzBZWTyBKMhkZuedpuCTMFGm4M4PViIMCO/CHFleXlCLTX329bkBdFQorx3Qlh/KM
eO877+Szk8U2LPDdRL6ecmuyAalIwpAzb3P6HjGwhc6W9xhCTzYGEteikjFW5WTTP341Ed4krfNE
LOzotmd1ILJj15tUepqKD1pP+2GLHiZBLItd6zP2c//Vjqix5GKerSdB+Frc7XdwozS53TfLzEIK
cH4pKZnI0+H2TvkSEOKFnoPdTlZ6hXKRP0QZaltw+0kjVv72PkS3Dbi6Kef0T/UlvUrYxfKSUqps
Zur/di2vJnFN0xpW7QcqWCtWi0PurB/VCWlgwqmz1knJSlCOvWmOEixS/QkmGZo2yg2K8qfPEW4z
T+I4CuLrK6JeTC9rzEXSiAvtBdOsCCTcqTOGaz5313BDxthhYq66cayHZQoqg7VDG0oDvMxMB7WT
szdvCa9Migobp3+y5Bf4jftcfYAu95V5eU3NR17SOtJhVPex1hr3UsmRszki73xdfKAK8oRqqdjh
nSk6kT0Xe9q7V46yXi+WnChZPa5fn0+DX5J1nnf4NYK4CS39UWNEuB3LC8uftJkkEC91+Zr/VCRP
hNRvuUvxbz2HAuU+j7nvMT7mPfiVQsLJGvq1J5uTfBeKvBKJentUPapCqYMNvlDxpReYIfk2wt2X
mLfI0vX9JsypZ0LdExkFX5nD7e+KMCly/tN+7sbnOg0lTTHTOLaoYqZ7o6A8HEOJdNFb3AMV6Ncr
xncPBrWOnCsVyZ9YIyd1u3hAn5tOOL0LJDHvvBnUOH3tJM907jr5d239l4dHTBC3l30iBEuOrrsQ
nWwpV8doV9wRNPLq6sD9X/qh2V8v5YS4uPdF4YI1Ujwy1RE281p+VMPjb4I5bdso6vmhfIsWTNSE
vKbdLz7ShIvcvJYCV+VsFkbM75cB7Ka5MW0UGXBvAHZr/BLPWIHsewnRQqzEPAwVJG67uCiJ32AK
ra6Lkx5kUZ5yUMLZGEFnhfsLxhuySXTa8QmVjd22UA2oSDzbBVNdneKpOP+fwDnIX3Qe2tihT5wC
FeAcYNRz6zwStOzt2qqbG0HGCHJHxxcV1e9AN0kwRYV54PYUFYfTrHwEPvSb2iaUrA+g0ABZOtch
d7YSNxyrzsTckTAbNS20r/yPmzvPv5G58IXcqa2BkLwvuVcS8mhVpDsQtI0CbNbdApnKzW5dlU+K
a8PwnjVE6U4zMQ8pYUZ6fz6XVusPiqIpLEySfIUWXAP6+K+3/gDP8XRBO1uEsE0aBupCqgSfb4ak
lf7GJTDSSD26uTEOpIChG6twppPgwS7u1amVa2pRs7qAcUqeMpjdAwAAGFJqe4srEptjQ3zOqFfh
1SmuTvqpkJSUlnhpOBxK27j8LaCezDnnznWgnEwUca2wBZfkOsGkTaAgn4ryjzsJ8line6aWDORJ
jU42kSEFLIHBD0H8U8cXJkF10yEDOi6eWIBadlIGQCV5yLenZYOdQ5F9L94TU9GUbBxIUrfzqDHp
SArEOjOgLw1rYfndJPEk51WIZACY3DBM4byGSOWX7eFAftPLCQUx3FPe39kO3/Papem0lD1oN8v/
EOu/mK27T7REjYIN3C2jwPKt5PbpHB35FJq/AZe7jvOQmZa+dsPUX02hmm2LMh+Sc1JKFV/ZPPBj
36Boo1Smq+lQ0jRgI1J8K9NMMCZVS/UMMOLkvUZqVjcX7IZ9rjvdRe7YoadEuNfrnLUY4RevBVXz
5QCj7Y6ZAZWuAu/2n2GoIYH4xF2l2smsZ+ir1OAnNKyLofC8icEZKirOXVUS/aTNjP/Fg6kiFX6l
Ogm7lPgYgohbUZZkgIR/c+3mJ21FfHTzwCLcb+50HmALXxAKnPKn/hsuszp7UsjkNh/LGTybjhPK
nFs2sMBvXn58F9tIaBYZUmfMIWZt80IM5w38k17G8IcZ5q9sdFxfRDaWgkaFsVPS9Tb1QN+/1HFs
Tt8jPfOhWwCNV0mcihlxXc/mOmMVtmVEqzu9V5S4pEGhji7wgN2trzOI7ce1DwUTBc/2QcrNeHV0
V/R3HDjeE7HIJ62vRAnEETZ/yddaMxzw4/BdPti0OoqwsjIRkD2N7z2LR68o3NpMwFyysvmS8Bn/
J0istj8jDPwjTAG7YVA1woAv/p4+L37roDmj+wNWZHeS7A4RUV0NHDM8wyYhyZMXKljtAywQE1Kn
FCpRqc9KDG1Wq6Cc34JdW/GkM+K8x5RlMXZKVd5m9U1BYpM4zvXoFPXertTkWtwvoFYTHJcjRHdd
gYNLkYZ+xgZdxf6itsWzjryS+SLJcNirBd85f2hm2bR9ziuz1SA/XwnU+b0AVt9RXeqYp4kG6Ppi
vASEJEcEbom3iwhVZCez+iXN4i5Oa7qn/ABhhijAQ7i4QZt9xQP6SV2N4DUdKExUITrj5AnTbeM/
xXgdQ2LiRvyUWKK1CAmP665Gm7blBOf7qDsSh2wVYlesooa8mXEc4yjItSIPFmYIKoW4g4YWRC2x
eFfAhtReRsyU0fcCPfe/irc5+P+qTUGl9NxtQaiBv+c1/V4TvIBpJIkjfNge5VeNqkODZPgIvMX3
mUgpNFYMecx479gc6i1z+2Y8vwmI9uMZcR8KK5jHKIY00ZVujSqBSPQcQ2LCudS0B7sMd2RPOLut
ZQvLeLEqEKOTuxDryUT5ij7BAzwuZoQ+McL2XblDMf6UozZssHYUaL8X/Tmgw/Ya4UNr49TB9Qs1
wM9XmBroVzYbwkBLJGBRcYxDOBJky7kum597GNGRPlTy0JPkj969QWDzGWhjQFLs/zvUoR0H3c59
ej1WdcFuk8r6mFW7a8EAjPdiwPg2bwh9CfOOEjaKXSZzX4eJtSc/bu53hXn372Ue2wX9UPgPKHzo
p2tkApePCvTMkyAy2jElj5FyFV3P52PoxIJkY82UhFzrxkEAHGC4HyAcQ5L8MMpz6W7tyFuf5gB9
AS+GS88zFtdVXprob30MLNwfEmCufr+n2H22b2c6IdIBDWvD4MDG/7WcUas6A7n3sreXc1tdZhvu
wEJZFR+v5CyMZKBBYpwDNf3PXSeXUXNA9LtA+vMyP6748kHcZBmTbf09KM6T5G++da2WIUr7bTz1
xkFJCliVIJE1XqKP0UwBMdKTBkHT0Vhntk2vEl2g3jaC8b+Fhb22u9MTZm4ltffKiK1G6zmwN+BJ
yv5DxH38boz76AEHcU9OpAyoANUE+LhdCE1n50YbCbzrTWtbi5IzYuy4BJEsRPRTYYBEhcjBFKd5
/ZoprWxNx1DuavLeejPZgeg861bCUZL2uKjGJE9LWk/2pGcgeWbnf10/lSf11/pswWdWgXh+NZsQ
jJkKF2/qjFMbVWoB9sxXOrfFIw6IFLj3f/HFmBC9k+UUuxO7FtAxv0/VrhEKwUFRUgJpHFIN4Alz
lXDCLNpBjMnPFfk5ZdL7TksGEqV6SOayTMxyvaHqQbyUdoqE8HKysZxPhLaYylzsbvtf/K7q09/d
9y5DPeue/SPWZ8ecPahwMKDk5ojjxqhpBOVUZ42ZI4WXJgyJkh9AtlFA7KxW12ZpyQ7oyZSUfBn4
q1DaSs9FOIF7c0p4NKSNZye0FoxCZ6UOv4lZKSfjYntthSedlaOv2SzEOMdo+F1lPL2ktVLyEcVx
UrT28hB0xQ8+GdQQ8Yi7BGYM3hETaKHwrh0LQ7GK6hCQbNdRIBjuEfzT32OHtbMOLtuOwauGtFXV
+kFqzb65ZP6brQ02vIKq8nl6H26mZwrNuonROp1Afph8LDnv0k5ud0hbbZ1iqbXQnMCQunk2xBB7
bZaajtsesWSNRAdRT9SHgTgbn/PwsFNUyqkX1SuzjRKnTQnmJ/gPT/4eegvkg9T9DSpwc+6YPjMX
CSEcu093B1RTjhbGeGTZc5E25EuirewEkgWCoYRsZEVZ4eotVOSy36OqM9Ljj7g1vb8mFHJ35KUd
xBLzIe3Var6QFvHAhojWe8uA4A7y+4c1wqIVQJSKMLyk/bIWYuLBcJqEZyY+g18M9rbIN2Wyn73R
w/TFnTTs7XlAPlzMT06IFRUKyywhWjmmCFsuMEFrQSyjD+4rgmW03LqU/ySn8l6+KwDEeO5D0hhV
AVRYl/iLmyhXQC+EG1x9l9JOSLuU9J0snVG7mb3ABYis7pGGARLHw9dgDD8SQtd3IMQM4EU5ifGZ
TtQJ4YFSnl0UqR5Kj9aNlns/iWiQLoh4TgfAfFnSiC7AdUbd9yo6fXCPJBHY8ns/iYz+voTGaw6Q
D5AWCGuGz5GUrjDMdEh8PbBbnyqstjJ1fhMqLXzjSGOymRKVnk4UJO4qIhgyeBW95QoN/n4ggXbc
flBZ079wTtKkqVepM4Yaw40GOcAMyTY3O1jB8p1gzo58JuQFPxAmZSe2V4kGgJKKfrIm+dduiTSS
BIw6xJz/4bDooViS2vZkXyTUY5XYD66X9TIRuwx6PtgUeF5HTUYk8Kex3rl9ebRpa2jmjr/9jvpx
JoG4M0EGXm2hfpUuMbd9cSPykL5hIO9bWwTvNakPe7IbJrFTvWi5BDL6GNpl1kQv/O1tzAtY/DsX
59uiT9dTVuehOvpVHDUfYu8lSp90XWa8XT6fqDFvEQwRiXy+uV7+m+jvOBHAyRU12u/wxvAZsPqJ
hNFnWHwcDvnTWPsdsvE2+wzS/F0e6fDO5g8cNwYuciB6kAoBlbrkb9AKleIvj0Qbxq4ZaFB3Ao5s
XGaSbYv8OI7iEBCcMwdr1KRIvmcMxugPP+2/eHoWJwyVVooG+94DA8CrU1X5iDQZBwWRfjjsAkla
NAXA1VxuGQ38Z/dBNIewu1TsRrtVviqSQ+ewUoZgAWSa8fbw9XvbArQ2ZOKYrqqBn/xX0uUTEmcV
RuatjduSzTHlqvrhFS+3Zp0VpTcfMITfQmQi2PLKbo9q78T39Nwe97zGfjLBlPgH6nI8/zggcd7I
5gX2glbr5KWPSvwgxpA2j76+ruGUVEtpZhDrK9/IfCL5LQIdu4miMpCOzN5AlYuxuTRFYNYixHUw
D8MYM5F9O6O0R+U5LeiY9F0QpgM7jCGL7XOJ7EvKw8GGEI9lQKEmgaywhN6fB432yoFsX0sWXgvm
OB5b+rCHWsy4j6LVMYCs/cQgpjENZGvQhjR5416RRLk7s+uDj/QW0iw1HMDbGSIV3hgJku6uQJLq
P3JQhaw2avhV2s6fJJ8ZiK4SWCQ8Ka9oOnGkTWzRfoSz608TgR7Eovi0sPmMtEPaU5JHdTyyRPFv
CUOTdUw8tZRowgb72eTnpikW1ebrCmegC3Vdvdj/0Vqgq1+CV0nIxLxrX93Mnodl7QmTqek3YSwO
ITRWtr+s/wrfq/dDgRsbxWs9m0eHrNzglqsvJoZRWztTC+wXUO1geeXbkPjxzKGiYJa/sStb0Aiy
IdcWZ3SE6Be1+XM4EIweE8HZI04r8ZR3E9DVfLZFHyt4fTbOGEzywBsv/pFvZzgTolgbU14WV8oD
HzgdpVWqpKFvl28G0MUxsKCNm7JuPybxNPsqkzmneUQ+H/7Wlrn3ZXkWfnwN0Ku5C4ekhkVzkbyZ
ExMKg4mQfRp2pwmdfvodUOFDaa6ZK2JAm1fByYGLXxkxbyFgHGAZmtOuvD8IQNMIdwxJaasqxd/N
4RpHEQF1Ffs5+TOUC1PYzc67sE4TykJhDrrXPrIZ/ePNwRagtNyBEwszT+JeurjmUJJdo5wlNDqM
S4eCDP55x59Ah8E1NYpYjP/ji3JsHxjafOG6xbAJktaX5y6rhrHB0OmH98AO9At44AJRuATsFriE
/kJsusWVJc4EiT4NPAP7+DrP9cAJzlS9GJjrT0ibYSoFYQb/iZEByZ4zBSjWtnDFSuFvSxRs0+ZI
R+PUFH9BEY1BCjV6C8z7HqI4rDRHz3MkhwzZnxiTfUIXooeJWx/YxX8EcnCmrRfYsLekXm4XW/lL
PIyWIg8yNg7+tr+lzonZ5Ww1XnT0F5/uWaV6XSpQGrl5SGHsv4lxDeSCRsCBlihcPGpyp3E6UcHE
39ocVh23k44uSGpXJq6Sk5j/3Y6WfpaXxHQABywqVVNDTKbPc7zpG7wTEVO1ccPXgvWb29CCwmNw
+uEk9mqJXaczV3f5TEVImm3FXRTZiNrHuhTvt/xPsjho34EwPp7xP7q01yUT+AcRQxf1GXpj6k1F
/emEizW9wV6CIDj31QZsTQ4oif41KTb+w03kikZEUuS0ROFxP282QxYx3hx3n91IJC0OU4VE/q9m
nGEs+cRbKc4gnXdqZtXm/Rm4FwvrMM0f3wcURXSf8tJ2gdEwYR+fxIxu8+Lfrw8B94brTISLkjPZ
VzWjpi1OYbfSRm7EUb0ylNiMJr/uprO6o+2wP3B+HbEImBF1DI4EBpUREWIEa0a5qZ746msHIbmi
XjjsUsr83YYhGFHy8Z6kgESWT8lN5kDMXNGLwHBrro5wWkYEZel2OjcDfb4OzqlxqtzL5tLlokvF
YFOVRdMyPi2mp1RlKcG0qDincBXQ36vPmnbte+Vl1qkYVfguVvEgBRQwZ6p0dvJkNDp5PqQVhYwu
GaRwJW57N2CAr/gWgLA5WHqonRn0DqMWt64oJV3OXeahegjXR6B8XRZ5cVPyv4xhUVr6WfStEDlZ
7NqfzDfjGW9DmSvjmFR4Dk5dKe6wiAn+YKbaMbFI942XO6f6pj2rLyM/CBoHYG5hER9+0QsWJgrf
LZ4PyHlbbKkPooWQCxuZ3qJHJiQRKKh6n1hDOxmPiAttLgdydvWxPaOmercocFjx9mu2co12J1sz
rANKGEY6qFByWYfzZa/Mons4GNOuI3ce3nK2OJ3VcW+OaUpBQ5OIHn6w2YLMypLgCe4pUx9OFhOM
oGnVvG4CBDBGbe7NMDxzlg2rZDkVjYntblAY6MfIvBinejQsx1cWC2kSqtTqhZCWa2vGuQC9ayGF
lJjL5Q3UT/A0OuIzECHnX4HQANLrxtkIWCdIW0p2mlshFdLJsvQOUvnyqBbmrtxndWU8n/Cazkfh
8e4kdi2GQzUbEW891XBfgp54ZV/e/CWjNnlAD7ma21gayVlj/srKUVAGJ8irDsY6uMpwQiF/DZ+V
x9SnAueYOf6avNrYgrRpDyCsbF2Glox4vJRcKl0+rO506kKk8hxey3rLeQnmTaSYBWiofnd7zovj
Iyk2EO8GoidoB1fIyEP39lSOfbsyVVEAKjrEW5XqiGktQ5PJy4sP2L6Gfj/BliiUKEgCK6T+RQjF
aBIiSKFxIensDeU1BstzkuB8PKdrNIDdAc0Rp5grtvLkWk/aBrV3M1CgvfQ8+pxcWEcpouHbYFZr
E96EVvZEKbwc2uqLM2Akqrjo6g5dFuX7OtBjbGtUTO4XzuRl0akqDV5FpJwCog+5dcSTouDAlL2J
1FbtiZ1dfSw/F36KEPY7V3DjWNmJTB5J/MosW8LCnTWlaiSdf5HDUGILRUd7tj4Ve5sGUCpyqgo9
Q3clcv4k8iQD1t7m6BvotmIxzTVqP9xXXJ9a6c587/Bs70SkeQC99XquhNdPrAvd9ggl/0pNcanb
Y3mOIXj+4u9nRbpAzob8qQah4zRxig4qbFQPnqQtE9qbL1NRKCoK/4qZcCVL4BqWXEe2tSUCTZt/
Q0YgNvXkfFGowT0QGA7QPxJIHgsdA4JtIbiLIY1UJK6RZjOW1oBkymnQFq+QUFx5iyCNjnVykL23
Sf//yJIJtYXgp7n1MGCTijadCY1IYAUFeNcAkoxOfZ1rZ1l54QoWbvQqQSc8pnKWC2g9sK4DZbII
tsuA7nUzmIMaawMR79mG52VSz5kY9Xfbq2O//bnAtNv4D0GOIc9Ascz67KdujTHEEf/u3ueDPDee
j0btBCbTVHYgO0DoJxz3hFU1W8wucyKtuk6OMJQLEcaw6mEkV6RJ5RAkfii/aOzmArLnRL3ubDUa
qbLz77A8JjxOQESF+9Orf1xG+5wByOR0JHRk+/P+QWW54WAcHNnio/5zEorbFf83dkBCVGIoNlnu
M4uyVuiE0ASsKWoPAzaRBRhq2ViXbIW80LDxfsI5x6oBkxeJWV+8ZrJH/2oOOsJ2cAnM8rXXfqN6
VonTK85r+yacWbOFzuu21s+x+Veb5IJfPaTpRj4JE5SOoG+gNASDIe4S1+huELjMimoy5SPpk/wT
Gzblt2jGRLKCCzpSDQTU9/BroTQY5DLtvQ/0/anUZ6OwJDh+s5TiLNv9F8REdfxjCierpyrE+BwT
O443fNE+7xuqXDEqitYagoN9ywfpPThJf9cVEpA+4uDk8pq8f3CoBopCzedTj+ftkQt7juB0gDTZ
8/7JQCL48svunD1op+UWI55TsKlbpKiPmBfggcPyvJG23pWz+NzOrxPBxuwPeU5T7oPA8ATJJ8BY
cWx5agurHKQztGVx7q9Dd9UMRwumEzmdXLzv6m00w3rdgdU3TsIG9xKBo4Rp+SIm1S8pjsCyY5N0
VwO4BuiHozxcYHjQ51CMZ8HESki5gfoxLeN7cE62RDDuBHjGmeKYRzjzzj/+foFl6TYL3TBzRWN0
Fw/n0V2VXuCFns1KlUYNNAPFu52ZXDXtfwaaGmZzhEiAkB7m3VK5g3xr2lzuMImvk6SN7dgzdSpB
7jfx6sAf6reB/qwe1ddy8iwIMPv3H0hFyo6ObgGiRm7w2hEZyV/AwGgRMpsCs8uWamqsQwXdZMwS
MqxITa7bHv/vdX3Ql5mcWi6rYze0+MMVrzXJBA9cndbH/aETMS89vJnJwKg+6eusnVuQH970GtlH
s1BQS/Em/yC4UcVI+x+o1PrpQqQf1eYx9NELaLVQYRFhnq9vxatIjnMMwqQC0TBb/8o1jmg30L1d
UC5KfS0ZHiwGOePjZbqfPWsusyoDqH/xtNL+1LCVgcA+KwPjR2OV1hJxbbfrsWtjS6kzYxrZa+Sv
G9Xc7hUbQZ48MprBrMXajAoy4BJtj0xLmBVAbW6TOs2Oo5gyx6O2DEVSqbSZVQ5tX1ZnW12B3YKj
R9pYX5Dw6A1bYgnDGgVZjxiHQBuF/NjPdvNmwH2hGZ69vvUyAOIFa7OB0ek5PP2yF7LmGee+r04p
KJfoCIUp5zePqCZXwXnlHRGNc3MLySYhi+PbDfNKL+iaYIo4qZCtk+kJeHmvnyqnOIyqMWpsR7se
NylunLXe3elscSlZrpefYqGf/xYCg9Ckqlj3ZgOTRGVmpjT5xEADXjUwnVYZ8wU5oA8OMKOwkCWF
+yiPNrT4zJAeWjZrUO9r2zfoW6XdGqkfSiVDlBUugHUE+IbSby36HtX+ojg3KfGKkCXwQjBuSIb6
dT6p4B48s2V6E1+PPy2JqBHTSxqsRkSEPPVyU0qKoRx9wItoQ8XMr/xTnwpTbenWUJoffhYfdURq
ljXlnuch6TT9/+DF8x1aamZCab+9eowLmHVM87K0V9WBmbA0r0akwd3JT6rKCao5tUoJTw1Ksk5X
7VClr4ax0EOCcCQ4yEKsAJr5dI6r5hvqEazffdPvh3zs8nh0rqvrO3JzE5NVrAuLRZ45ZWSIUTFM
rQA1IEy1RNISpEg2BX8a0HFW+VAe6nom4FiE5GUdcDEHbefFxbHaZs7853sc2WhOehFlgqqmOYR+
59eIlKqWqN7mLMHmWFiCjrTCqtPhsJtz4kQKl5zAWp5ysj15B8Xu9ceWhLDTF9DpZ7EDAwCdvcfJ
5J+eaTwsLI6RxuME+ClO4fFu+vKtZYakrRjkbUvzV06460h2oAN6hM0duq7pqVZavsMjQxvKVEKn
sZO/I7bzIh794uM1UK8VmySy0vqNbNyHvScQfA81cWsYRj2CLkWhq9PQ+PNTNXxKjLS84Zwx0nL+
YLMXTasrCPYPjlY3K1e2moeaPVo4YNfPjH5/ZWRXC101xZYolkpVjG73hbfIFzlROfb87iCuZrLU
LGyrB9S2KGUgRquNuEieGN72ANI/UAn6Ro8a/F4zg6etC1joREw+OcD9mOCKDuesLN+/ZsaMnP1D
uqf9dDnZwhtckD22uzveTdAhFGziD7bmVKMfR2MCfzgZkbF1EKv1tXQjK+dsBh6tJ4Cn7zcyMFeG
aau/obFc/MYNPrZcetXTB3Su+8gxVbZgKi0NsSoUc3xrh5ofZySzfEN+zZxfw1gReP+engA0RpTv
qPoaYx9LNxiqJPbY0UxY8mf9jgL+o9/7gLcyodPatuzl7n7CB1a7zykUnhHSYW74KHk1pBRdltuL
7IhBpIk1aRQfbsGRYaMSgm/GXQSJG1EytG5hjzp8nVbyB8YSnd27vv9+N3OwbCHPqK92Y8JPYIsZ
Xvk/9vTjW6XkKLj+KIPaYAvaQm5JT7oc9TGU2O3dJBIshPdw4VNyQtSdQmRg+1fKwPyzEhy90Lkt
BMJtEm94V2j5eEfvfBgidAVi09zgwa+1aUVZFnt/mNKwsfL+m7+yN8cHmGiGg7WIo+EAG0+lfn/8
QsXw3spDBBgTkiaYvP0fqbE++dzrsC68QVsnlGHjinjsHYNgJFX6QCckIgvdjPZNo64zlUakhyYl
+CRFm0bI7k50bDEljvDbVZPtFVWcPPOEI8PNYqHKsNJaTdzkQvuwiP1oYKPk4Pf7R7dKQixr+Msg
Sqq8zYI6Zt14MMSv4cNb92eRcICv7eNfQjAUkjJGfj81jEumEgWFzGlWAXdTA/raVgIQKYLYn26N
M76oiKtWvC8WT6LTB7+myL+YuSJBaux+G3hpq4pvmW4subIqOwyeJs9M2AXjFiblUAM00hTqFKIc
G7dWRvPJlS4Zfj8Lhd8Mmwu4IL3m6beZdF7fDaXBoCAVMsWcNAmQvJWEZ/H3UsuGJQsFxsJbVnl0
EUCQ4sQGKIoxYbWEAdRy7HeKTm2kpbsE071OncrnhpjQPr/P8wBgTFlrudYQ79DvEHPI83GCQ4/d
lDNGZGOoQ82g8X2uFNPPGRMYHtHTXCztLww0WohA0W/SOCoWHnnQcLC+V1H0Ubc3ns7VuSsTwhQ7
yDmkUEQIUmC/Vbb2HtpJB5AgQYV2DOOKWJW8pxI+lxF0ACOmfovT/1zELbBEJ9tEFlQsNXw6gymr
7ndSgFP7H/beFYRznh0Ai8HboQPVFtuPN/3ausD7OE9LWptKKpMAr3iqlqzRtSAauxTs2JGXow+H
df87aQsFUXduQv3YuA1lczl0DAvMJleZGHUCoyXEpjuPjNINO5tJ3rJOPVYL1AhawkHJaqFN4yTT
3UKVCr0oxupCvOIOvNGKugPUioL1nASLt97GFvzTcr3eBicXEkmaQRzndMob5uDBu1BYnbKV0EWJ
WbiO6mDc70ymAK0Ox0n/5NO4y1gE9CP91e1TVJ5yThXHdrDdaCuca+H96gjCTsr/zMomJ6+74UFF
VxvUXmG6tdAzNuCxu0hXJQt39Bxs7FjSRwjATV1OkQVXawpn1JbpMzgk9Wg+8zgwHxFQPlZz/XzF
yWfTmnuJPf6kqTP7bCtcx7UH4uRbMm6JbGgRmZYXCZoKR2Vj4OIOS3mXv557Hma3cWmTfJffSSry
EJxfSbQ2icUnXod0tuIJHKXG7NDCZjt+bit+JCdCg3Epgf6VAKAtrUZZa6OGvrk+3odo/JootKX9
xp1PK4kj/tEi1uVa5nWgOk0aoYG5hhIXyWqbBXDrcPT0HAPCHH6WZ6J4tAp5IFZM9cgKCype5HlW
G3XBlGHHK7rY6+jejmTEXIydmDM+17QlRhGG6uVvU9LQ7iwDyK0QsQdb3yM1Eq5ywWUvpfh1Qcho
j7LQ1vwZ/9V/gk7353RpxiQtU7yR3RO9DRAw2TLsq7z1tzARLf001jAjv4NPmb6CMz7/W/g0Gomo
qhxGXEP8rYcEGRPss3m9p4s+TNlGqCFBDYdLEfg58npTkqEWyFxa4bbvAF24T2zl5MXjQ7i3BHaO
VzaeGxYNnY9Y+6gavqe0PDcLwRO2iIXTo0NcCD5Cj8cQlDu2vjXOTTaKZLCQCx3r5xQPSeKhEggv
AXd2cTihHbweF1mMWbLoHvBC8MGTFT43erY4QD0+7UYNWv1CqVaDqPUqvEVgqqsrZGTH9xLyZq0s
MfdqoGmJCKePPzfX5tMeKlj37rQOQ79w40KXaAX8D90dOqCKDA/9fbMY42ark3iOeYUJyiJH65jY
sbD6fN6NzuYukHEforYSwd53zE8UnjpaZnYRFr2wXCRZ4gJDUa1CKbKe2EHSXEVk6BpBSIJiz3P6
o9BZ9BZnhg9eJd1VTjJZL4mKZCrVsFZauvC5slmdbSL00AJJp4yomw5wklst7245jxhVPm2v1dXI
rnqwAOMFG953VriBNKrzdgkCI8GRdLkoIMuR7KNqwpZBoDx56goC1G6wyxh4hEOaR6jd4GaFTWi6
pWkuS5CgDly3LQy/qbzRl5WGd+t20aIBGcYOk/4BjzfTK2uuhMrOeQRyTeSSJGkEQ73q8qRsj1uT
blvtImXbd11yAIIeWGln2eao65U3Fb4NGIBkUH3rJ9omvtzLFaR678GJ9Rsq7+feLAfqQVbiCSy+
AYf8yRMtmKOgbbZIwtmHDrHpWf6BnlHz3+XlCXip8Z1YYMnE3DtgbzZRcVZ9QxWKzCX23gLa1HDO
0mMV/aE+LDYeI3tmIDMf+MTMPkMuvRUgFjrMO3TRIzEvtdG2Qcda6rABpMewGOLiedTuJLq8wJ+d
ErkcJJ+Z0+E/CqvrmeTxsZ87aY3/RCaqdbXMRUU91EvriVWOgKT8u5cQxlR0B7773/6jRZgn+qyb
qjZCsepiwdUhrgp+i/TGVTsaj9wL0kWP4ytFjAyq8VZrgHcLAOItFrbOj95UpjRGR7KzARFF+Oa7
f4Z6UsR9z+oiyN92uIXz+SJ1PuAFPaQYGGGfSijdpeiJMc0tgvM11QkxaBpeZ69AoWYU7Wq59tLX
DGft+srXBf8Ao+W/IxV3oxhH4v0seePN8NmM5LWxSViLY9N/Wc3rfSLEQAPpFQPma7ZAIVLkY8oT
s2JDOW3qS1kwRtpZ/f2sRvr692wyMk2yjn9+QGR8Rnmmalqb5+iM+rZXUMUx3zM43S7N0XLX/b0q
HyaL1OqNJRFMcbR6aENUKNwkzT59IiNs45I+YmwPTtZXF9p9LS6zUPu1kzdbaHY+PF5l8ScIU6G8
HejiKoczZcD+pcMy3jPVQY9v8zwNMLnFILtTBow7FibQ+mlVI/KnYvLs9oLsaMH91LbnUzsOT+5b
BS45B62DYLOXFF2r/GaiqDrAd1ogB+TwSyPHVt07+x6fWZ+tf71ySPYSpaB65Z+npF7qqBeGjJTx
BTf4q2dNCwMYkbKW5DrbewhsO/3Ee7hF9m8yRCp4M+AC4KQLQczo7ZMTziPHutDhzmUx2C7cUs7X
Cbr/TueMeyMVn1wZG2ww+MJhK+F3bxfjFGpiZWebxSMQBCJ/+1781mDEkEb9Xirwedox1rm8kw4P
5c5DsWBMWzxbtARnuNBjMVEr9Zhj/WVGKeL1w9KZq10Z7NEJWuQyNzyHEJFqUKJKBGq7cPBD8rg3
+intYuv9rN3Ob6v+pgtvBoAo2/r12ixrb8/C89hgFWrZkESDKewZRdHrGLaVkH4IK5KzuTt14NUT
Im/6nkKtuhA+8+TQJoqD2Y11g6CvepJQVW5WlvP2pEBpMgUFmNW7yMhXqXpYKs2PfBe5Nj28qXYq
WdBOCG8m+u80ZWXg6K6BCqDpNWPezBVeJ4nz3GMeEtuhYZ9mRS56OhQO9SAl7q+Mf1SFpkPb3QD/
gIpKz4Ki0M25YzdOLMTO+t4ovWGk9Kv0g9L2C9Ji9S7fD+mr1RkR6UtrG/THFpBBJOM8dtmsyLZ+
LCV0Z/OT0MDY13uSohw9ViaKYkM3xDKSYHI2CRNCQN7/BKjhiJ2tS4lAdwHuwvVAGZZfvKreON7J
rMVJ0BXO3SiOLLtSoLzVK9YysgHWwwqzACByQlnEMIRjLyOHzDUAzKMqjdmJJAn2qxIYHjC9JZxR
sg3DJaIAjo7ycYWSxWgFGqXpIy+aDXhYxkWrmKHaLBHSyPG+6YnNkavoeaeEnXFqUsJ9fkHj8ykF
XJdNuu9ZaCSKT6hGXNNmUnFCJmxzeD6HlsmeBgtj3hXgS1Hov9E8jbT/jv13qP5G4p4v4xvPoX9F
DYIscbUY/FWjqkEY/DGgTvKYP6cmH5d53XA0CRNpub79OK7u7HRPXfcJTQW5e5D25xdfX02e4qFb
FzAYkA5urIZZPMFbWqABhn8iCzB6eYToY96EbKapqExwToXjKPsUtivF35uioYyy3/WYsnd5C47/
wrAULUOa/VRFfwDzs91flaTL/iol/WdqV3vvX+dLe4jzYPBk/oo+0a8DP9gKjoxGsHsgeqwALVPw
d8umNBKUuVI2fMNsR16dbjPcW2vo35LoFx632moeUllPMVhcgfMfE7AhrlPgUSqZQ/uD6l+Gurz7
Jf1WWuAFY5FskuneoKs2dN0K6IVlgBBS+zRMMQLamXYZlIp3MqIRRYVR2itF1bWEI9tDJRuxGqM7
RtB90CL5KR/ZagwUeMgINxzieP0i8CoTz9HuhCQpK+swNiekcLMf2cpxCl+6O2hlP84h5e49W3lx
dTdZkXd5VSa3KkiaKkY3cwgk/xBdhP8XVhVneTwregdNZjVnPsS2bpDIonLPjXTWZ4hTwVwfO7fd
03QYi6/ogf72X3j2sGS/b36R5Fzzrcs/XhGLO0N3lxnCkVHZdgEczhxqBZyPCw1HyxSyy2/CfB7/
ipsmWFULpCIhgCs26LcFJYgpZm7i+d/FtcNx4sLhLwPqYH0JO3bq1FLr3s8oUUr7lX37WAv7aDjM
DRv/lF9JC40gLYabNa3dOZFs3+DwlJDr7Zwvxp11O1CqnPeobRbx5vpcxWye9/N/6JazPNgd+99M
3xCjGvdPSuVrdMhCxapIu0B9PaX9/d/6cILlv7tTTD7BGa9bJFHMhC9DTOfM5W/6pSrB+hlpOd0X
oGL8Igz7LrVspDxGOEU1lErseafxZ0vml15PWVNCJxIWnHe9ReSZFl6wK9jBibSbR57sCCB9mN/q
pZVBoJOSecj4lJnaqZuc4jQfRzHK1BGe3gRFV4iTblistM5OajDg8AmTonxHjwfOFlOqzhK5NDLM
/vgUv3mQC0ztc9nMuqLk3LhCEbd48NPyZ4qVcwdITLX9Gv91yuz1j2cKPOkeqOKbLYCeZQrJv8QU
aLLfJ7vZjtcgsZsDYakZVZu3CDGMJ4vdqdCujwe3ftiRp5vz1UQ9XSuI76HwoYTgcnTY/SaQKdaJ
sbQlO3QNCxHQ0VzNbLIufB58CXhnAOcW1uKFBUin1+7pG6WnZR5XqjW/CbrnRZDetqiAkwsIUp+F
+BGGlw2ei5VCG1VL1emGP6VUAmCaR6Wq7SNud+At3lBQ7V67AMUYztZ5ZywYhllR8tuiS+0DwhjB
iODSW5XKLvr3+0Dhy1J3MASc82pM52DpSyyak9oghYMg2NiOEzWURJmcZ9YkCo+tWEFjkNB5HaNV
XLDJiYU/S6S7eYqHYbeiTj/Hu5yGwGLF6EAZMgA9hNTVgKUQcFom/AfOqv9CwjxBGAybCsJkntYq
i/20GPj5SsJ45Lr32iMsGlUVm6aWg+r9Ck+DrZRg8R2IW0nI0d49TQ0AgqHQiZPPAu7EsGoPvly+
qlaX7TH+Oc37nJzWITXvYUnKu9oAsIwNBCftuQFdhtmUPSG4Cwx2tgxWd1NlW3jzKqBER7g1IbaD
2amCtIgZVsF7qlOZ2FdMQWW9aVvU5p/zFYg/9psZOREHv2zoZ2zZ4ER+4SK4GL+7xUh1HucN/+R0
swBx2YbZUw+HXtxb1u4rp0Kdn0B3Klvj7+yeyalqWWEqjVxAHxKYUT2t29KAbqNJb0HRK9kiXf6c
TU8IEbrd96FU6nJ6rQdBpj3/cxJmiKFtb4yVrJszOmffzTbCnrfSphRxc4sEsXmwlYACbWUqmKpD
JyPEUKHpiUEBx1T0+H+8Ro1e/Yvshz/bezeH0ydzVH0i1bd+xeUyobtugDuN7eL76MjMXtGL8e8I
fIbfXOd9x0Bt7HZfEQIBBxr/uOOUjryyadjKq2YDY71V2RM1ypBq+SiyI8h1Zc+znvCgZvx24P5V
SSelA7FgPfUEcs0BRaljIxE2IgChZ4SBGIdXu+OEl5dIt5G0iGYbhzB3rDFQ4ohl0pECr+Avu9nP
/QaOcSLSx7LcjqtsLbR6UGYgXgjy9BXy8IMw/U9A2hl+1met7vbTEFPilQtHW7/rWreVUBqEFmrJ
Y/HKoThiYDzhCNg/VuYaJZQTsZdON16l9of9vCH07HqQzRAi12UaQwx/EDW2to73qKMeqo9zQp3q
NNW2WF9wWpSzuqTumJrvvEOgNEm8rRHDIai2UnB2+PQ1iH1B59YGXZ/qQIJcy8x12bnSniMAyIi0
MDQYgQ+uB6spw5jgzV0TktugZzrqMcew4SnLEt3UmG5HDK2Rq45GK7Ehi2pQUDOC8ykXjxQj8Kji
XeAtQ4oH9SgwCZQ2R3D4DEwBpSzdZIa4CzQYGZzhKjIAqEJtJNQdLQ1CnrIZeTJhEFdA5A1aFYyj
f25YpdjjOrE/SqRDnzEIKS7Bb+hgefNK5pOKVjoCAFfgMInoksohazH41xug65vEN+rh56WstJoZ
TDKoi9izl/1T2VE+jXn5XmMmVQxLviiMz1NxSKWSL/tdOK16gY7a/GPMKydCRsePusugMGA9dU1i
0vPnEsYeM/WVve6x1r9IQGuF9drh2yOyniBpmIKvJAae5Ps/VYoeJXmj9pR39RDm9Sf7ye5gSXsI
GPwI0IRgQy6muMKPWeqGP9VjpOAfuTg2Yad5sG5MhBCkrD9/ZDuDXLBGIhnQ5T33Sfh5GqJ3nSO6
Ezgg5YO4BQnc/SDfB8PUNCj1v1CM793Ywj3fzoZx9/Mt8s8TEW3ZCGlq6meqbMR40A2j12Vpp4Mh
z4ihBjSNYXFQt8aOKCcdMgP/X5t+ZH3UOLuexcCWNRdEXC8RqVoT1aGb4PCzdOxO0HNqxyaqe3Pd
02fXoCh/4Ek/f8ak4vRKs0cobiM3/LywhtH7FW1qf82JG6ssAZPskw7j1EZT3RTqpLkLqLMJBqy2
cAM+Cdmn2adWz67iPH1vwnQWAuDp/QBkzjRGJ9EPadf5PmLTB1FRZT8TMeKER07+5HfD6hdzBtYi
VlbJWN/ld6TeBge9FaPVHrc8QNfHq3lod1ZZt3SG2LZhZx4gwcehY9FdOZsIbuO5Mx6mUGOOX9Cc
hwyRVpOZpvFfdPTm1HfYhtNjV2sf+H/rHkV3FXsTKtnC87ANwniTBeXw6CePrG8aI0uxwq1zW8bf
30PggNigezpVMfeAS8+ruenAKqRHZE3eCww2vxLIesj1sNZMHNjqz2Wt99EF2xjL+0kgF99Wwc0Y
4tdZhAPhz5HhgxmU0gmtkxOvkbKkdBiY7L99Li5ZFEeoJ0W3fRsZBJrwHGLIyXTimulvKOQPHVa2
JGig2qZjJJkXp3sCDCo6FpcG3vmmfSdl2zJVAsmKpi3uJ8RLQLNZOIaqfIk3W0d2q8EVZgmplNi+
GFttd4/06WzkC9YhyAnjIjsAw7UW1BOI4HkadN+gSzTANPdPjowj8MZF2PE2QEnYsBPaSv0RHVO9
C9P4WX0FRrUA+bBYPlsDfR4wzrZTxvZ87oo7eI7zkxQQ/M6++j2h8UE09PdoNIlgwhnp8zQfDq5s
OCnX0/SpKEQoyLjh1ETlBwKzIaTTS23qZu6O/vRtXat0NJ1yLfQJD2NjRfzGWmogA8i4tpK0ckSM
vdbmBFoiFZSeFW0dw+pMIsBGbWgESiq+6U321Gu9NmCJa+CPMp1c4HdhHnGikZGdfXaCgrWdTe+l
0jHGfUw972bgie+qYzs2bs/sz7lRBbTOi15+LuFBbUbGcOl+8h9V54BPGmWyGeTVAmuPjH1E7mG9
2daqs/qm9vU/9vsNdf0gQib8LN+BMCC3iDvCon+QA2vr2xDl4uQzBCGk8EmxENia4Npt2TsWiKJV
thudRUgtriQqrPoE4KUAxdqf0oxxf9vN0pztWEQg/5y0Ub+yNOKEP3+NhIKMpyBHK28F5z/+hnJi
M26jImqlyi9vHpxj5Bf8Jyc4yn1GeEYI/utDc/1BOQkyf0nKSAwk4LwINMe1GXbKwXpBRgU89sqF
MeXLwCjUQFY9YZK6EfLEVFxYJGUEqxH5IaHB9YZ7QhREl4aH5D+9IIrdltSlnAr+Q3Kd5+7k3TN1
K22PV1Fujsq7MriAGihDPFVBWydmGiM/342FhfRmSQZAdHuyi/8H2JEEx+RO9Z2T4L20ifVExKv8
AbdRCCVkuJXVvy2PxJfw9YS3y7hw2+eB8ikuGAdh29xSYD9YtNHcTPb53WZCguMOeUEFXKTcPsg0
hnSoi6B3QzZmk5kxYQWAaHblUHSW93sJ9VRV7qrLZFVfqdx/ys7iWMHgJzhDwOnfT5P7J3kmAA8w
CJFK9ceYdj5j+rhPF1UKUb+fP0xyakNsFXv7dYIVkrDOJNgIKohodvVd3BB+1GqUK0AbC3e9X3iX
a8hOIIq8xuwbnfOGMeAhBHQ5fvynKVegmfANIC402tNlsQD9YJCI/aIa5DmqTG+Y1XA/UYBdgyoV
gSqc35c0IAzPeR7Fbq7DsKoJxayCH3QN4uAYSfk+xqdg/SeTmzmmH4JvUqZbvDThs7OV6tHafus7
3dQosPMWqBi6o4zsW0TNM9M95WRWEoKelqqJvXDO692K1FvlfIrwY+kMwGtOhMFxnRbEj8wxelOF
806ervz0wQxdodpxDXkcUGSV+mLPpPYDrBEc1zZM3hKze99BXbO2s3e8XqeKpSGjXKr+gJ0rCpZ7
0aiQ3/Bhro8IhGMTTGRsBm3N93GPsfM0Cq5QJQ/vGeRl8UY94efAWB7zL4iGMHlcXxv/rJmQeS7l
bpnkRcSgpsjOiBolwwdZR41yVQ0Cq4hzIk75vCiRu8CG7o7cGuYg36fRe72NR87uqjVH78Bn/Vl+
+6YlMP/R5kyjfL2SHtVKWD2ytxPEl1NBp2H5bRkEESn/wzqOjUKxLxJlCnT3X93HlusPgTVhKOlt
7zCpwlrm2NeY2JJzBtURfW1NvvRV8ylloR/VODsrgddQA/Yqn/5fI1ybN3hAREW/2SIjWcZ0uAHa
qkaJ5erWgtFhD2cmjFa+AAr2QQgQMS7IMl/tmEPoI9rbzLKZDaigFN6ieoyYl9F8UPPw5qgnz6d4
sA6ODY0bDkC8dQ9x0HunUKTNNpTIWSz/3ZQePaXAc7m3WS98ChrcNi1zbCjJMeSjDPx4164ZIOvV
3S3/mCsahfnirG87t8rF4IqS5SmJw30LKje5BlYao5/FyINzpAdt/wMy2q69nCpgrEpv3pa3ea71
t4Qp7a03JnVzID+wd3pUmaIezNeSkxOtrN9v9gfQ36btja6WYVIFpaH76QVdgglUqbmPRn8GZTES
35eOxmY3yNa7B0n0H/Q+XzBCBIRb0o0OmqR9cFCVqypjwYikyKEvl1J5wQLCBAdP2QyUOmpwP0mM
jY4C+1Ay0IAiFwqddPBKobkCeEyFe7eXYlM0TnktzWknB5epFT64wS9d6YalzLvVy5U8yIIldTwu
MWf0aGpjU0etluChjQd2Qfwf1z78kZvc6rfVt4PU0kgvRz9xUhm3YBpvmH4l3UKBdpVH/mWYApD9
LLx0FvXPb4gSX7+2PkhXikUhoScW4jPhWLLvLMQpLnZLw+cecqm0NtMKJ+2KZLtaiXRDMsGrWBHN
wAOZbBmmUCmekygAodBdPk87X4RyIcFVKM8ZxZhyVWFbz9kBP7/8pKWoG/vSjj0XSC6lqvtpl6lS
1REy6MlH1J/VqBfoKZQZcG4Q0qElxc3mFJAxugtCH40rM+Np95IIoarWCZpqeLsIik+dr1bWy9vP
Btyt9jjh3SUOxslEiAUrhIR++XDf2uyljsreTq8N/jnDlDeARbc9bOfRzJLm7cOmre9lLh49gDAP
xxNyizR723eCiPo7sZ1uwx4QHJpGD7W0N+HOoalZp4Csdh9dgI9WhpT7E1SbNUgjHihhHPwbnd7z
bpAAFJpQzbBlBp2Ujmnh//O+ZZSGAn4EBIF7HXieqPe0d2lf1B9qj+BPlOrKA5H+jGeP0/nobc4H
vwjIWX/y/zV9OIGog0wFg/2wft5M929jfAVDAxHoVGDuDdqSs5FkczkDOEAFrRtxNGp85a5I0msI
jnECWQcfPJKRzrmf2heZtHOb+Kb1la8uJeucrBi186edRXAEbUfGmVdm2YSZZY9Z8UO4PT1Y9fUy
/wvm6OTJX2mVkFjcSNReNZZGG+Vc5xmY/IcBdutNefghXblNBhvsGg22l5rs7RzD/XE1MUtSShnE
4u5+5/cTu2lUcPJmP3HzOEYg/6HdL9Na8pHaf2H4aMUXjiebWTtG/9yuZw20SuIwbzZZ2lzwAmFv
EE8M8pwVE2LQgmjZoowAFzUemUSSYT4g85zHH/lA6Pt9fXT8Ok/7tbABfckEbbaKLspQHDQEHuP0
BdYahWY0Gtusrf1GdMF8YKXTdVy90IO6tWsdRL8vH6tjSpjO9r5eWOmZcKqQ22HJZny8B7x8nYG3
VMoJbZMkMZ6ZqlkPRE1xQM+9qgQEr3rIBCPiEFJ9BZhAK7Tp2o8vUX/Q8YnoBxLGVWvGZ5yI7n7z
NApGrUoUD3lAn8VqJ1C3foQewUChHckPNQ4c4nknhm5vObKJ7HmFW3HYDyaEPsJSYfuN9hs00Eom
befumF52Rj1/BtL722Mj3v4C/Btl3vyDSCfgfyviK5/p2Z8QxFt/dw4n5QNaAfMA5Pjyrm1Tnb1Y
mZMhnu3npOimGgtqe+zrZbPFHdYUNN6SqMtH4ns28jylW/4w2abDN5KlC8RKOhXcjUadFHK0VmyK
1Z7npl4zMZFITfKJttfZKJ628Fr3kLMoXhxjvLjvPObzBG99HFPhGgRRbD9aKNMXGX3WBjzxqyku
X6/zOLaDLPOJ4pxHDhNE9zvAHHCDn+90iUILJt1UGuxozEqOnOStiQyzVvACeqzPK9883e4p0IXv
qqb19hhy+jInKYp2uFysVeqnkF55Up+Txu87qfwGyMfH502s+TUkwr56aMyjuQM+koFH61qoIkY4
m6m3VswV6yZOpKP+aogs6CLo294sPVZQjXXQZOj3Nn9Whb5K2ECWIpLEjmoTWCEjheiElqLUOxpV
3mZ9TwGjPlnV3SSax8JMjLwITbiiwdeWeOr/i6spEUsEBiE8xOxposFtIHgfqprdBnYzCI9uaoAh
AOrg4tvkIVADpQMe0zdPBLc+eLmuZjYmJ5XYN+PrNfK80M4uCGWZCA7mmzIVoO3kIfF7KCGfIuLY
e4+tWz5GqxqRT1TbjYBJBU0JEH+nNSsOGBjyjjXJ5utWuBXETr8XHUyT1cZ534I8QsNRCECfEmjC
zvgJDy7YjMSk/blhLMKIYMrE8GdDc47pz227R/tz7kcf3+W3HkBy+BMAbbYQkBNuF+m80QQDucen
6JsZvEBdLaQ/i+3A5VWmpriuT8uLVSAAqN5xI0qN0wEEyh+yA6DzMsnNLqnHx/DH6EBMON/+uZLD
WuAx5ELV9i8MBRquAeUSDNzPYS1Dlz237mG7++PRx8dTMNolls1WtlDtC2kvew2ucfHTNU0jq2bO
XmuwohqnU72L9B2UWYTASTsi4WWXJewqd+M3z+L4XT+wDm8/opXRSvqRitMTlTsDN9alr+7eIiEc
kUZglDHFfWZ4ffdbK3rOCJHKF1JUI97vzl0vj9t2zwbJ7Hhs486mLK/AWwhb3LPXR9SfBWHhFpKi
UgTxif/oWDu5qRS7HKSx7JjGpuFXEJeYf8nvVFzXJv/V1GUjyif4eKaCAiabeddiHHM5YfSh+K3p
p06WiRTnryMwRfcFT9VBgRxWxqj5NFXxrSue04QBZaPn3RFsYgphrOP0wjAAbWRzhNj/YWzvtJJ9
I9IWLhVAedpuhsgjAkkgbG3l2iG0cYR8jVVzZlVKaIJtg5o5ZmsXMjf0xLGfl0L2R5YuycfpfMlz
6JFzBYpz1zunO2FSz/LZbeUfvvLKxkr38SjqGHaa26FkeIKatkU3Fm9MiCSEpIDNDnmQgpQLHz7b
N002gPP6OlENy1gIRLO4uMeANtP9WF85fIa+uCbf8Fj6dSmfsGREEc8XW57C33O/F0nzilk8iXAs
wbOwHvl/bAnDTKxSzENekaGwV/W2tBeiIDpPDtgo328VLICYSizYUZ7vkLqc3c0zzQ160FXavQUU
WAPEsWCEqEAP6iMFVir55ztf5PfTtlwcCnmqVO0Jcl/CSAx32jj/sFUN+unyffz020PnT1MGXh4U
ifuNutQC2fim0QXuHjItNivNco8bfAo8u0T24x8atN31sXpY5oc11O1Uhdb7gu1lA01djPipEM83
nntU2/ZhteJSZO+FLPiQYnyIhNjvRJbeuC21DCc63GLWoWZLfSkP9I9VsDRHSPghqu9yALZjXYfu
khZCGdVjVrBT+7vA85Y69QyBOeh6Ib1/f3jx92KSZWvB5ozFYgcMHcbV1HgyW/V+m0ZMGAhlE5hA
4CG8Hj+zwD+4UEnHJyG8LdZmg+iOaLmjw39S1UMMe/eA3VMxHXI1d0P9BtnsIGtKi3yVl4rmOicm
YeLE1281nek1Os+68xEgHH+irZFljaC+B0igA5mdxG+SufBuv26nA4BP8NpJYbmiCuQ7Wlk7R0jj
9rnwxkqqvgRxWDWSgHlIVTiqQlVVxkW3MmXxYjqEIphWKQnTmpbiUDMBoSUZzmFtwQ1F2lIFIl9j
M2Rk5hjNrWndpu+LMw/8zJRXr832JM5UNm1SqTuUo6MarGPazNIzxDFC1LHwOF1o/f+eSelUxE/1
L9NVwnuz4ExhDU3hHHXx1A5xBcZNN8sbIdQHVQsocfl7sswBJ9X/kvWBUJ4WIbvxO7KFINeA3lgG
anUI+46UUT8XvEOstsExIaOgC7rKYl82PN2HXFkPiYc619m7DkU1a4uFSiDqgoZYPE8/sb8gzc/M
Rk61GQJVwmE1mpelaWssjWH0IH9gIeEjOjR/LdCoL8GrOui7GuTLifhfnMac9pOTwd60npu1Nms5
RHSDMlNGtm+Apmt+QQBLwIucGXPyzE0MbCUoKFFiuqK3vBrYKsaWtf5KC8mGXXDy/5rliXkYx6gV
zdVdlLeKm6gXvc16scffphxBxLfN7NTrZd+ODKl5MzF+CmtUx7mIGIvYQP3bRt8zefaV249yRlnX
Ls6SpaPtwWycRAXjL5wAZZksNF9Lc8UcNGiKgECcEAfaoy7prAib2AZhWIOju85GINYR1XpPzH4W
j6HC2rK4A5fY/hR2SF6RHPz5LXwoKvs87hQ0lrZmic/+rhRAjkrfl8iu3iSO4j6Is4c4uPDqzM2q
cahs4KTu+pkdtCpPBmLs9hQ4uk77Fqb+FOSZBESSzBRQGTRWsHm0HzIQVytQad7Kq+2jo4c2jDdY
OScAChR2gOxdtKWEIClABfcxXL3Tek3lu0EkYnk5DZTDvZbiE7mMn+YowCHYydrgHeWj+kJtwmvC
McD/4lyU+iHPoJvmIfbMFzpCFgTANhxe4T6c+p27Kz86xNjvFNvkbABXrXtgzkvjToCzmG3Nveu+
u5OAEuVEY10rrwzMNahiBDgLBBnmb3Qrm56NGRz2DiU6z9Gnv/E67ddKWYCjBQCJ29iWwwxoLEEc
ha4Z7lb/hN7+6lOj6z2GeodhQzKod+U68it+pv5iGFiZ51BO+/sG5NfZp/LvAQlt6mdl/DClVwdy
uoQFRKapdLdBMIaO/KFZoGbp2XjW1uBDBM4DYDDwboMJsMhu+Vzh/0YYifwNcBstYrCzvTgDihYr
n5d9NuOCmFzS4iZOwPdM30pg5r9JhTU0P15x/oh5X2eQj22DnFb9KmOr4RbdMMoIVrvgsgERfJg6
YuRU0jtpnjNnNe9q3QjSi7d6/0vDcLkOwJgQ1YLtT7HHtPJYAtpMOO5FAFwdvy076T1kb4ufN8D1
fH5JVTItyIhBWP70JKAswy7hFLpnNEjR+0Jvn3lCmbr0lD+BDe+/M9wgVpYGy2PLdHV+ZtK3I+BK
5dxA6QObSaquBgmeZA++S4X2HKdZ2mc6bgifnpecuwG3qN3I1o2baxvYCtPFD0iO1VsepDxiaP6l
m8CKjVO19nP8nsrnhwn2B7Ih4u6phnBlm11/ivsOjmaEVmDPB2DPNUE4Ae1Fjy0qZCUhF9HwgbOr
BlWcl5lgoIvVqN4tSTlwxLANIlGKA2oDiXEoKSKIx/6MEm9I/RwFTl5Yz00VTpo01cZaG9/gw1HC
a6iP2PK4Dh+p2poUh+MFJS34qsns7BdUoC+YiOUfXk99fTHV1rQ7AYUcWBnF17agymaSG2jLBPA5
s4dOKjrgbk8pNRypkuaze/UCSYIS6/ELygi5DE42pOlFE3bwXhRLEFrMzOwPgMl8flNa68SjvgZn
VRkukCKNmfELxZJu25zVTkP/FcM/i/6mtpHrpRpA3z/jTvloM152pSbosP7nhktz+6xmxQ55AnDo
3vgiAt9c49ydbcaXAikO17uZJVc/EFTKZ78sancksL6GS9EBd5YMv0FkkL4u4BeReanmyuzA4XpO
j1/w60PHGQCKc8Z5Ys3uPwlc/TfXV9kA9guuQ0b94zpyfFbYxeUensn8HB3Bf05qZ51KXPVG7LFR
qsCXbJwG5k411743mV7TjytFv1jl7RsqKX2FzPT34W1eopE1R12htahnOjBtH9G+iF3HgB/By5EQ
JL53SpMVp32MqD/Ka7jDNzoHo4rwpODhrL7RwRqNgF7iTT7Vk3koHQVY7jgDzhYYu4Qsva3XfRnb
hZslwRMJtdKu4XRZko7wCVhUjF2+8xhcJjt+52q7tcp7mS6MhUP1DWpkp7NOyfpB/5lVKyz/ztga
bd6LZC8/EEFurBZLIG/d0dwlO3Q8hffh4PJG912PZdc70Ekdce7yeMM8YNf/qBrTsB38nfD2qoXL
iWDMTWPVpUCHXDlty6hU+tliu2kvUURPxRNZDyiQGtXvOlNXYuqYbdq97jbXCS5HDAMJ+rPDIZ/b
BHYFrA/Qus6pabXuPGU8zmNZpT9gSYLXgSZ+Ywb6/zfIv6+RHGb+ApiP9UvitDiGOfJNFJl6mqfr
9NiwAYYi5im3wNsDHCxjB3/Neqq28r5F2U9+p0kdROghepoOfiR+Moq8RpbRVP3ymcsXlVzdfI8z
WrVuhRz9ADJ9yTLAbU2NPDCcMxmsU2mbQl6mDz+NzMja/wWcDHEXTjBsAJ7mBw8QCv/ilHVq9Ttn
toO0cNxWHfBnVCksRLBTB7CatAtnVSgcHIBAcdOEsWFicHQ8RvqX4Dio090tcyUurSV43IocCJZm
1O0lGwsBWr5DfCKt1LuKZ2MwkXYsvZ5cnXRzZ1qXOV/+vS1yC9OwkKrEp7uW3Q3ZQ0NrSCGEuJ9X
RGXHwDcu7tsVEjXDkgQ+m5pBqR0FNynxLSZFWMokondR9goTQtS9aggJXq+qsH2tyvnUeF5pWKxM
zjWkMnXcko+njbQC9LhV5j0LxZYTxRk+e5R02psifR7e7UygMVdgZq+h29+1WHbGZ4w9SfAJJ/cn
mAIHep9n6yaMrxXb+bv59bNUGqey/sRoY+lAEIMdz/QlCphsruRuxUPjoVWGgP/jci8hIIhzFJz0
6m54izRSf4uGKJMcdxtPGgAZ8xOX6rlARlpEt0xJpPk83FuS3KJxl4ULW/DdMCIOg+101eXKELW9
UZK6azuQjNtEPTclsVceGShslsDzr4PnPGpeaJlc1w0oUZ2GPZcBdfhH65dAv/VTBtUHKkd6uLA4
IJBnofyWEXKTOBMGa2pFeUtZBAW2hJVlDSMzNincCur4TeuDxNOxz9G/lcn5/RHLqNcLvybz56LT
f1ojpwLhMVm5M4eDEtfYD9B07z07vNO7C0a8ZTx1LNRck48DHnjPXpyNBbrhGl9MkUpaLlo8B7Lf
ltqJyYG7ua7ZDaXTquLgIdczin0xignz2y6g8QVb2cKy2lkqe4HxsH8TgRWRCjTv0iKcui9iUGbG
0n3JzJUv/0aetGiq6ZV3GOMGuN95Q+g7PxKCg/+tZORHY+8SK6aTd+djG4u2WgRFa2Q54MCMfR4U
3g7HOoL6xOA2P9WIXzewI2m79AHtBxiUHYTHdcqQ32DuWrJykVfLQV6mOrLYfmK7WQbpBibV/exA
DppmxEu0s1XoCYBumPJOkjxR5qrYHPZR0Ai3yPUm8J/U2zwlo32qFEhl3783006+rpeJSu/yTiyJ
KfH9hgOhZeGHVfUD/0iQVd/Cqcj94oKdjvPrqsnsRZwwSE/hY/KjNx0C8+LOaWbSRvuMNhgr+yeD
si/rQj5tzcMT+fUM6e8r/9iWb0DvYqDR0zOFfkaMY+wiH1T00qNpubpkJgDQantvmE2+sCHifT9k
j3BeEqcZ5QzvhikHQbE1TgLn3tDMUWWs/HaC5J3nRWCKiFfuNWNMdTtV3oTe5tjMpgTw8+eaHSDt
yV+Ej0sJzBnGk14vDUKE1n55F96I5wHQFH1SnQFA7jbxtSzAkAXOqd6I/gq7hcw8j8wtC3kzBRgp
Y93N6ZmlHXGfxXUjRtBjktrOJnAZRAk6GMZ4e8zGTh6QcrEJE/+e+CXR9AdY66HpD8qFYV66Gcz7
kESasUtz9nDwl+li1uSmnOwXxOZwqoW64mDfTCqX348wOI1/JWFjtQNBw5CxTlAJZ5RVLIrPRqbf
AseaIQtoj+KmK/y2S/g5P7HZAdPDH/zzbZx74fUjapbq+FjmxCgFH1dP98l5empGKbaewW47rCuh
Rg1mMfioGGUyPCL+so99EV5JdcbE3oH0noeWAmblp7mXFD+gPVlCmkIBy940ZITpUOACZDkYhGr8
FYsYPKy9U7LGdB+GhnI6x5Q/cSrJQd0T5y23az7ZPJQPU9Chnh4wSvSPeoQytXGAOQ+xfN3oy++N
oTZGDHFfPNherR5iJPXvHQxGRfyoZZGGT2lZYUuYHIynWp+wmuyIrBl4HWsnHB+/i2bCfjrYw7EW
66NVGt2t991OLi0oMpc+G+kToSaC9e8Iswy52IsgIlQIL25mPMaTbBIr+56iDstc5xhLp8ppnCkC
xgtRemvQn9+GoZ2HxsS5TIiqoMnQ6qKHvPnfAyEpglUpdg0u8B9rHOHdfP1v8U9kySyQSPt//jdl
9DtBrmXnvjVwzZv82eBZtVWMDimeh/fmGBDtH7NRT9YB3Hgezceue53hXzF1Lvvl7FBeykhogw6F
Fr5Z7xk6oLprESMVPluDZNd5w25WAcJOhifJ2sAvzNiyFeDuuOIQQaBN5tUqHVdYAZBY4EbIGJwG
9gyZm9xT4PkJPs1CJk+OjG3CZuDpohc1druQFNmXHRTqFEvZXyKWw5IKvelofywHTx7Vd0M5m2ya
dVkoR3/lADLcJuRyKa7gp981xSiE1L/Bba9jN2Rk1USGZUYRKWh43zND7WAw5CdJhRNdBHZK2gVz
IVPXBeKWx83TZ0HjccNxmGklZFTyTOT9GvaxHwTAzAcO8r9jg0Ls4BvNNH4XZZD4Q5w7OmP+netT
fjD4ZW3pkGYyZoskgIs+5dWNM6QaXSir5qyOXourAGmyo8FdqioZlboFVpfOVzVopjr3HXSM/kgL
cA7KXakS0BOuTffykMNskMmKgtpUsZoOY66VI1r6udTstBYsB3eBQ/bSXcXw6RH+Z1rS9gSrXz4w
56xHq3eSlqSGnqwxPP893z95RY0Pnl2DvKyEUdCDWHhh8H6Wh6+MfW0E08DON1Sh+yJuPekE2RZ1
y3X2nf14w90DygDQ4BR4J+VHxHdnAdxk7kVlS+44ckHDTB/RMNgGxPcjHoVHkofInz34pCTBl+0Y
bPpCrEcjBdzZDbLLzQMfy2yemwyZeHhlDaKB6kKCbn2IpDo9yONDpcauUaeu8+nwolabrGXcnl4f
jfntXEjEkQBtrTbpLgh0Q2Q+Hh2x9Y6q9do1hijyG7aZskIqWgfuPy3SLSf9rhAENYx3IFoleSLV
3crp4PKhodj5FLA6c1mT6UADHZ62NmKS8lwogqPyyuikUv/FCg+1Hwi89P2fskTGs4E0yyGiOEr0
d7vV55q0ASHubnZ9pyefPrwtD78bIMxQRHOa0qvMfR4F2Axmy4EA26FblWIRUIC7SAf53KaTGqUJ
TIShxDqRg55anMX2aqiS1R+3zRuH3SjQBkB7nR4yqtOnmgdWY741cnuQV5lu2crsI9yjWLU9JKI6
Mul0V/FUhzBisV6D5d/yLzqLcmq/lHtCEjfYUEn5J+qSZ01GeenHxE2H3S1iIbM85jR6UryK0JwU
7DYr/nFPuyT3pIykLFD4J41U4yQ/ta8WDGFqmSaffZTPxuxc+f2x3DwZJwAiD6+sOPl6ALNeL5Qb
YOGkTGKQ7iBFAXpl0UC1cH6dY50Ve1uGVgfTbT8upvUc4FivCB2z/K96zSTDauxi1E6A5ya4hWsu
2+7wlwvqxWvBzQID3c2qPSldZ5wCF73LO3G4Q57/slBdU7E6gq0dLV42Zhw17pTSnSDB70uBwM7F
HotqzJvEYuKiqDdIAulyjeUFEm28ZS6vpLRVuJ9FNcMhq5IbG0rC+rPaHa9p8xNYqufYixSmBREi
S/7KUp8uXSX8xHaHdiK9Cj2sTEzlgUPPLvvYbWpzH3S98JXgS2N1chZPx2IzRkx6qYj9xoCn9C6t
wxMjLkNRd6eX6p1W2YNnamYjMo7XxJHg7c5wWX6HRd+YpJXDO/11N2ClpJ/1sx9l47rm9EfBb7/n
CYn9OMU/5gWw+ElU5cksbZZ3tCmGwpsshJGOo8wwTGKSZ0dlfHz9YKfttg2ebQkG0rT7T9B+SJS7
HwOcxW3n/y+SHuNXmy9kSpbgiW8tU6mOVd6DssaGbRRMq5FYxSQBMPHBcfPDvCXUh5+a9Eo4vBER
+tGjA8RCm5StwaKF7e0duYOSr9y+SiOHo+5S2ZWbMMTrZdwDOkqWIsP0crPgkLTWMlgaMdfcRjBO
bW5U/nCiU+FGluuLh0Rm5jOFgVagCTQkuoeWpDUVliN3pGiowLqJ0k80z/r/v2UW+t5Ndl8etQ8r
lD3EDnqWHdpP8yC6grFPLxU5ZIGwEIQnShPCGhTQjnV0HsqFpaDPToffjhn3gEyavNsUixJtwnol
Mx813kDe2r5SFeax0jSVZ0/MFELtv15JJhgAiVKaPyol58xo/fsof2QBUlO5VS2+6MaTygexYdfx
Dx/7T+58S+XWFJbL3ifIJ6nTbrpZUOHFOI3LWL6VpD/ryQx1t9EfIODDr0TlIzB3TkvTF3TpDswG
ltp+ArOgNAeculChTo+nt4bwb/8nUXOeji57D01Z9VUveQJlJ+JKM2Ho3vecgSxhiMzWfGw8L+LL
OmOedEH70rs4tlVVLeZ0WbhehmBhAPdjrWxQL5sECTJBvqSF13hLVRjmQTxZT379vQL9nDb70PSQ
vbG1wGKuTfm1HkOmkL20vA79gjqSatzeT6VdLRi3E6B7/9JMT2jrTLtzlgaMu8ZrN3w4hO05DgFp
Q68p7yEnSRj6HjGfHiaNXGDYhhJLloEIgykbyywJLKyuVs6McxYDLlqHaRjLOVJdUmThfw1D/aS1
me/R+1tCEx2NNFjQZDMQNKslQAHyCtl+u5xoRHSWsc3i7vy5/F+UdkcO+HZOGmndIqUDSBqq1SBe
BjECb9rzCpuDDbbBDmroqUACzV1wm+csfSJ4y/suhvOOH9GyehRyqF742rfVsFRto13cJipSnHXV
BVUwxyWDrI25qm1awJFdEAFcgFJdWK1STHmdPKWEY+jPGe1gdqxpgKIjiP0BCyE7gH48uGTBQvQA
WKUpIuXjx4SbqygxODiEtIXyPO/8ontLonPKNCOYF79ZrLqeVWwUiq3n91vIwDefVgwgwtpKXDTy
WUVGw3CmFBcKSer1Jc0u3CfKolq4qtC0pHXnF9AahQzhEXlyosaHdDc8CmsKUuUZlHZixWVNRPph
EwemgRrNELGP9UU9DQ4z9t2mJGltJ72Ni10bQEx1CrmNrVk+tw85unolESCiSfSZ0KBoeFNaRpAU
nKff68V2Z8J/a/kL33OYjLwRNCpsDREAbf4T0pvlSymm0M8NTCUOb0KS7rcaDDg/nE7Ez1py8hVL
8rEOGKQb7lOFuvpbp9FFg0kjrAjBU6mziiIFYkR7hHY3WPK0a/jBr1sAmbXRnhS9V5yn8whFPORU
1J62mnawHFnwT10oHOf3KaEBVKgbazhJxAhhpXTQX17TXeBInvKFBc1TzGAnhc6NHd7syI9QSwfX
cEPoRMksaAX9cx8cGaVlDUZJvFC6xJLDu9bRq89BflfAe0sIVhQ/CdFBI7+rlGuoLc5/PqZGIdU8
xdajbiygxTlEFLdydypVqqcE2KLxkAG5+KFx/YaWMWb3mJIlceFA0U/sK3TvEaBhC8QBiAwOoASL
AhCJiFZvumkkpKMYqAyKR5puZ4QQhLs8gHlQKP7vdqUcxJp80MGQin8xI6nqxfwi12xhcKFfvtML
GPx1x7jAwORGVKAYqN72mmMnd88P8GQOWA5S0tjnEBrR+Q//sAAOSmYi1xT7QDvwSMubyyqMjjri
VXamvLOEmXo7FKWK+e10+ChJPyltRZlBxU+olac7iimvNL33vyZWpdMrO0RehRNyQBLrG7Vd7DWq
eBbiFbRQTg7hEEG1bnJpydQazH+AU7tFs5Y3pXVsYkML4SK5Z9AYs4wzaMEqHqIgxV7KrXAn8I47
9nMK1SChgM2Mqm+gbWPD/cRRggrJjauUs+sMLxp7+kPPSawVNh/CB5V0oRb1Xu+d/ednA61XS4ex
bBmKzK37p2DpvhMJzQHYpAfnsQNP09fhWMgvkFi9/fPVAILlWNR4/87pe7Zy8gHsAvr+olBA/6xp
/sK2aabrkVeeodmgJzssmO35MpASq9p2Aw5s+bukhgTdCenLoaZbfSTo9K4fVIAe/0wDng2cS0/C
1gZ70k6ffnkKT1wbW36z2weNnLp7vUE5liuxgEU0ypk8XxyWOkeLbDj/tXt/V9GZGEmf7t1rkB9j
wqOTPamDYhcTBj4j8vjtue0thgbh1hyOBH5tPoiLNJfYvWsAM4HGqSwKufbY/7XXBUGl9t8Qgp5D
+t2sWU/Io3SJHrUKdRq82jeRVIxVLAn4SF9OkS0SxhOjDRzEO5pHIsFyOWVkCMT05J4aw1+9YEG4
sHmNUpVCyvDzcvgsZYlAXF4YPTm8tZlmI3RHKVmD9NiaHK511frW+kB1HYTdsrWEwPvnviLjBCat
OTPiZm700+rz2Yj+/IC56khROJNj1UNTmTSr7TcCBTs/owB2Za44yGZCfONP85RebhXntJ+nSOYz
DZY1xP+1fKT4sUFNmPFYTdom+tlCcbbA0maWwMdMfjND+I8NnRTdRAYIY2ABGrOngfeygp+86Rgc
dwK8hf6LC4G2aIBOvc5IdRgpngsMhXa+D9XpzT+nI3vjOkHpNSzXsqpBWrrUjeeFR+c1ZwohhZQq
hepoSU7FMjeUcNkL2jqvQ+tzDIrxgRvBddtdWLDtwfc8r+Uxlkyyj9kbtA5wgdUtUnGEa647ERXD
QQpI5e0Zq/NEE2UbCTfSRpLsJA0gu1SN0mJsBUqittu541VBrixYLgzwGVt3sKOFf8OKkN8KfMlA
6qYt6tIgpGdpc72yd9BAGzictqIqlHJJYRkiclSdNtd9UxyfbN+Lb44x3VtwzSe1Wzm7V4sasHD7
bK/eic1rNJW4BQvPDhjojG4AZKzJCCd/4U1AadNl9j0HeK6vbKqNEjs0lBGxuZeNyTyloyF5EWDs
nagGk6UYCYWohDcSFuYhtIM/1XKpEVzWjRE0Y4SZ5YvYrmdDyEp44Bh5oH31lfFnr8lSXPCDiT5X
brpqXUubY0gwtcD1iIyN6jZlGWTadiUYIjYIRTkVbnAPPDEx84FLagjyXhPc65DzF5U4UrMmrAtr
1Mb9fmvRDcBDaQWnrvXmjpOiGCRRMsCN6t8o7BRQvCvM1jJQbmmfaThOQcpXdRsBHOak7yICBS1S
L3f+3N0BaptTrKwIXvbyfyuVRPgtkBZgQo0SL+NryYaUhKgj2ADlKlO5sSiZkt6IcUdsAf1dET17
dUA/vXjX/Q8qvMrvbagyCoDnPzBzKxu1Xqzo8xss27iTkWAljyyhz6RMZHazRdHuo8GSbWt9eEYE
kmLeyfRD7o6fpYQf9CiiaX0DlWRs+DJlhMOccYn33/svapu9O4RAB7O6JlVmKO3MtAk4Iq9Ox2DH
5n/Glc5aCPGb4Yu07qcRVsKliZs9jNSXoIue+RMN7g07+5jW+qmdHpRue1pVLiCtTx18p/Iy3Xbb
EPJtQVb/QKK7dnIL1kAaeOWxWNo+mMni1TglMKzyQVtltaG0o1+HPHuaHtSMM8AADTyef60B0YBw
a21kxRJhRerPfFBxaJ5meadzhNfYshyauDPSxwK168p88p9aKaUlmruyeXPshssXSFX44E7WMlHx
TnSgz/hIJdUdvpmQQbTOKSdfc3nek+VQEnuwPEY/1wvDcockLfnGiVGqr/Dof0Du44a9db11nILp
uUt8nARyomooWtwPnsoGd2lMM+dERKqLaY3c0SogdQnXebnw/AIFildJIZy6N/2xbv/GMP5ZZi1u
w1G1QD8U8MtNoXX2kovMIPZX488i7LpoDtoWw/wB8+qWqf0Pa+kBM/+SprcenqG1ql4ffikGORQz
z98xf/lHeScTbduSUUo+rUXPunqoXtgghYQjdYTxXbScpsHd3lp10zrrUHIHultidcpj0gEHr3AC
Rg6ZFvAv8jrv2Fze8Fx8qZAnhlR2SFktpjfFdyw71SlZedZUSBbN9T10bN2aU938uDYPrh9VJiVJ
FNW/l45glO02u/oiVwpvLyfK6GQCGkS3c7RYM3WPl8eS9BpF7FPFIo7r2Us8gZcV4c0wIkob1/Rl
3TGHqrzuwK30QXwB/k1MWNJtTo9NjxspHNQx8y6N0BDOfr2Pr15n6w+rmhEuvS0RtDfUHT1pTkzn
1+uad5ktJEiIbZv8VxUE93yle1OjevezSORU4ewtw7IdxUXPzZI3voph5Ixfv6LX8FLQUHNYKnbA
yBRfKLI5xLxHFG0Ry62G7w6zIsRuDEaYCaDU2GaqoXfQIMQJMhoT5KLFwbR1V1m3dOZHjKOOfP97
+gp+wwA6OvQZTTq6dl5JGEB1lPQYW4IFuN7WfIGKZKJ240WONQVra9o16BqkLOpOFwgdQLqfYDJU
zPI61KE+q8xgS5pYb2zx/9weORECHH0YIvhLuxBzhOeeksuT5FecXCQnblxyQwl2gfHiQI0m4Cqb
hJ8HlUxk5lPm51BT2N5dGncmvJ5PmvVwwIqIVn2OOzD+yUvdRFvJY9Fh7TqqQ/vjzeR18gZTiN8l
A93My0JlAIucRKkedfyC4O9DE22nUo5UX115G7l4SIb1NoGHzfhEwG3IKqReGFPy9X8HDSXWExaC
Q9HchAOl4YWkJ2e0agB83eTVZL5cok/b7dnzK6URfMswYzcPC2e0FJ00+BKLwKTi2TRHlY19pPqO
rxQsGYD6J8sQ90wg4zaM+cUxGqOXxuueT2KA72uXe2mKIvKOOMxxNKQQJEQHHEtsemX9j6ObZ3Hb
WdrcySBzN+Xz7DBKLTicFII76iqI86YEhC17QBvSXBBkSYdudcaBStCgwVsXoAjA8G4GW6fqXFSx
bHD6sSNPaOjz6PwvyVDjlYGDa1wIJ28fRy1DWABm3JmqKDLffYn9Anb6EdXJHQOMAwOptYRzRBTe
gVvj1gjCXHnBWcT1RGt7Us7tYTSZo/ojPS6Nn7CBOt/eN1ILcdinmR9V7V/fOg1BvYWwsdwcGocV
65//62lzb89SJpIhYKNFYQNW53fS2zzSBpj+hwncHVPw/tCiyU7sVQO7U/45MbwLq9WsVFQnzTyo
Q5C/E5p9jrlLlVcamgVW6ZfwodMZ1LrhviRA5iE8x1UJySo64B9LwxqejRoU/wEumPC7Y4fiI+3R
TRGoXy4d9CG/g6NIEFXCca589BID1J7XQ8jldJDT3lCwcEgQwtnJIS+bbLl1YD+sLqqJSYYnFANG
Q8woiEzKl++I68G9Gle2Oqe9RpUSWub5mjHPJjvu/HlJBTMNH+fu5NFxmUmX7RidzPv+sMKjW/ut
ZW+8zFj/M5NADd5I4tYzYkKQxMzjAmoFlj+ecHNrnuxdDRHe2sPmMY9ombx2wDFG9xo7AZPypz6e
WmoLTlzIBASKMmR9bJEEyvMVSu4shr37TxlB8NHsDgZluCqKLHcnT3cSMnaN/2R+RvPmboiht/uV
97qGpDkKCTLi3jG86OcJ2v1zlebGNCAQGQ9doO7fT1K969bmoMbGk0+heNKwCnLcEM0F7eyy9Y5H
1n4EZVMQ/1Z369E6XEbvGWmbt35d+f38HbXWdXwoe39bXZ5WfAR4Wh/hoAFTUe62pWTWzDyN3c2d
rBtZQEtyom9YyDiEGWcvLWcWPRZ7CnOk3QyRT3sfahMGw5Nyu9mnrvvksf3TSIKCZ5vlNYpW/XHx
iKjmemMxa+cy3HpaXYrfhAdFvdS7EHHqQuIQbrZZFBHoHbmoTExl4a3FCoCaDnjqf2icpC3U6zcn
PCbIVPD8uoFP7++Kj4SEjpA4aoznTmkI7ZQd4rQBRwjwjqGnv/F2K7VrFFp4HR04Qyqf8xINsnCZ
FvQacJAcArgjn/6BpfxPdzeyUgUxI72irlVCyceKhu6YuKyMluoAK8MmcFacHkvMHKVFAk3TAr/o
sL0pMZiQd3vzp4Fc5Hu35K5jNRRAsMmRbbFQAJwF6yB2qSZq9IuMyKtFPQdvouLzlj1NgJHa2PEj
fkZIMqLd2CbAcioTPF/xa0YOitHqvhHgI+OlqG0kIPPtwS2ekAn6PI9l0rqqQvvpawsK+PhabqNy
6FqJM+mQFGHHuF4Vn1kdGTXPKHC1mtEI0dXRw0hjmy0B4Rf83WJt0l3SQ81+aoW5eDCB8G7t56oN
tZOmurbPZPk9cMs4spWfzDcQpXsG2jGHDtmmPUFI1F1fALVowjP1Tiy29TGYAzYcqAh36BOGBS8g
mMwV8WMNGFeQqOiTp8jDG1r7ZuoNvoQwtfD+vvWPkfAnlMCs/LopHaaaCXEkorFHSSoaRJFSK/Bs
9dTsaHo6j57vk8GuimFtInVhRB6KQfM4YxY84wtHxDDnEkwqJ8d9pg6/bu3W0v+k+xLc9ekokcoM
G5jOkNBm2nXaVOD8/NjbbNKGdPkzpEuEMi3tZnv46f1qzDBLD6N7EOU2D6gkNMDuInsrbg6qPuk+
UvIoj+ZmT0DiJ/cG4aDf5SelywjoZdE46uYkT4GjKKZLIL41cEPxN0t2KedBWGxBcs/tHuLff5ys
1NxIafp+ErEuBbUEwj2Nn1QDNsGBxHiOOhZYFGGeaVShefR+IOrcbZBcV4QGvuWqEk9jjvxfuLGi
bC8L25ju/HDl0BSqkmIOUZyY+4UCoyW8qxCDdsopBlrEhE0TBbEOs5ITI6Xc2BV3Yt3Jj/MyJuHe
siTfINHq2RDWNvL3Da8RWoMHQ2TGHKXJDAeoO7RkZZCw62moVgc2uPqQPwCH/OvCjNAB1/DGy/bP
ABz7Ni9ZSzqKgwz0WOfKJ6qdVlGzBpK46jDUCSwiv0c0FwWg2Idb4qq7otlZFaAUVZW7ktyyDtkF
CflG/DXyXZDJys/ht8zbZJu4ivdNCWDETHy8ydgvO2gyJB28YQssrw2jjamELLa56/mpshFifDty
tMv7GjclNcC4bz/JfCG+NvSoTGvrZNh2J9fTo+lPYq+s9WkPEnwTu95ncZOdkl+CTG23jw/j6178
6unbKDlEXUsfQV9kRoMowdt4a1taK6z62fY2iVvZKaKa/y8XV/lE2KUoTwVSb/PRGbq80cjF9Cq2
WSFfW4p8pOu/57JSQkaTlXdV1PcA4KECvRfLa5i4R5uzP9YtgcaJm9w33C8LSr2k45gmpADEl5vY
qdh/E1BSrcjnuw/mUi3E5T3qEAae3kNvB7gjqacNGn8vWHBZuij8jFKDJ/jDDPz6nOQvffzbLOD6
zM9uIIG7UWAFd0lrNQVLdd0G59H4HREJUWH6slHKsqvYTOVoT3nnGKj9D3013iTnFoBFItDx0t5C
qhwhwO0hp3prxCGWgkK8rXJkCpGAJeMMxK6OshcccAvyEDX2yj95ex5Sc3Fe/WJzKKb4YdFR3ujB
Zp2PWgumIZ3tFd2GiNOUnInwuwl/dDVN3jvdjAvIt8ILoT7iV+93H0AKXQ+0N3Q/sEgQ/CBZsnfg
iBwBP+Xy6HxaUfzEn6RI1FbsyM2jsGm3o+pW+c1gAELXJufvf0jAtfW0d93axX/+poApQYH0AN/W
GEdr+wnHCVXVaGVNnwcKAauoM+X3w4H8aTqshDUqffe0qhT/ukGKEZZ+XnxK30zyT2G8JkPxEZD5
j8tOwbs86u7MaFxHtRNo4uBBZmBi3M7SGoNhsKcCntb5FKpqQdTMwcIJ/m7C4gHs1WMRfcGTxWkh
1/TK+dDsznn8reup/UMkJnJb/BYnMqqImjShOKMkpdrPPDgVnnY/kkCp2WNebVbDyX+soRlzWfe2
pTI5nlXy1+xFb+tw58tT/Wgeju4pvf1oX2m/201CtOMN6gdRY4eZbjCzX9wd1xBHhohj7ndYp0Xw
jyCKGkBlsk4E3K0BrcyN/i5P6CYvQHesh1mZTpVSWUr1JWR6s6tWkkefJ1P6vVGX3xqbTiDVwpk3
ph8CJGFl4jRY4p8qbPI02HM8M9MwaIzE0M87Ql0711ynh4sNr/eTyPAtRqr2NvZPts58txzHzBvN
RHduIMMr+QuO6dBHXfI211eCzrBi1HbkmbzkcNT4aykUGiUyEk+Spgf+lIIbR0gi3FP27kuJ43J5
wfTsoN4w1O3tUKYDXiejFTP/pMXg2YbK6K3iSKft+1/CJXIbLMg3ri1wOrQIavqxsqbbbInCl0OY
UuxRYbEfpTwxn3k4BVZZ6pfhIOnkMkVJPrKQtD4nyoglNAXJ4G7GZMAEk2slmMpfgcF/EzuLY7El
GPgNjHTJNgaUFBaCoq6sqW602JvjP4Ka10LEf7kgQSOjJfdqvn6XtwxByt7b6jvRE5hH3M0PQVH2
UcK6zxE1cnCgFAqfwvsqAXOq8wQLucI9+hl3UCxB7vk5vVLYVydByd3wKQm1P3a+dQc0Q3J4ar0N
qy0q7WWdgC3fjEqYddauQrAwb85kBBW69ldodUigaPMvAEbeZ1AmqeOWX4ybAoQreJadDuwfDHtj
PVXfM8yNxzjVHjgasQoqmM4uLlGH4+PNwXoadIbCssXFl1ga3ci8fVti4qK7eSfzMCYIEZxJxj9b
wf+ZVy8n1xcZbxFlkQUx30wDO9DIfG2t7ISEuNWEWENEkoieZdrUG6Ndd2/qV2/xGVyACyxfIDHL
v3tbSo/sqBt+Co8XzeiYhaXhYblolGBd6F9FN8FXLr9+pZazgRqBq80OQxVr881iWTUa+NlhR/HM
646Nv4ki5CBOe7n0h0RUlaDlHJQrEgRGv0/Mdzx2Ry5ImErfjqD+zVnnkxFc2bnkL/AIDz7ApxoG
qnGhG5xbRR81ZJVaXwTw51exht9eIvVyR72PMhlbDTYx/o1QMfg/SIsnOId3ppuk+JgN2ajTrhfM
EEhZ0jm9epwRLLLzZSrSQ7IfT1YC8rAEYgrTFQiB4U+bYAQaUu+A0KvQBriRvMle15041FoBSf+l
YblTv0k7SWueRWaHPiyd59GPN6MDj/HBp0iypgb83niUvWBdZTZCXbO8fbajSfw5sBgZR02PO1Ny
aZA4UQLnLI8HXfizYI8OPWsNAvMpzYmH5SmhHzgXN8tyxZ0zps6d6ixJPSkg8xVPrUVB/yPanha8
GX1ZNofACyOwBU2HQp3d8+9VzQ1pQay3HCea0lb8iApI0N3JL+1lcvbf1yFPUZmZ3dpVpElV0OsY
YfUhuruSTiKklTqzJI0mdO3Oym/TV8Y2kHlkX+qH7pnpjP+wmyhLXyT5Rhk14VsDgFFywO7WZ0E+
m/bCj5iBZtH3AIppSWeXKYI61+eLdZh20uMY4xO7v2EfHndKr69JkP4B9QYgbLCGdJK68TUBGFzN
60SE74cfi3d57ZDIrWgBwyiDAt7jcnT1gXMEBT3n0iePMO681BFnZdsf2r/EwEaeFDHPre64qOsA
cwEsRn6gQ3a/4/Up7eDjO5k5ynltTJaOWDtGiflzNA2RSfdqfmrYyDehrzX02F52hBFcY37bXiXA
ll0lcaf8Qgbgc4lmFv70Vqh89zclosZDj2846LCGiaIcNkRP/PGhXC4eFwjc6iOeiXcQ3Fqmw3pq
jJli3jDpYyrqSGaryRtwNN9zo0ySwscpXE8OS2TZLhgsEOYvufkVEi9NlhRapu4dVYtYPFaiEyVB
f6OEljNUgGqLyk8C/oTiSxW6uUpiuQW3Aioq3rI+1xk7+DXfXE1CCxCLHHrf5YiWleAHSkUv4Xal
0/0URwh2NTMVrEtCKobmIGHHv8jowHyM+2ailC10544XbL83LOfG0hLVppJcGE9CveYBZs2UtvPI
eHlGpmfwnkDThMATrnae+VP/gbV/f2C17eeYZfPV+sFloGrzRrPeBkJpelBNQgEFER/9GP+oNtv5
i3MxuIGjC8fVpzJwEPbfQEoLAFOspIx8Su6j5tZ/YRJuQBIq4RsjA7EMN6RdceS8srzT5lc/7RKr
rEILBWeIhX2mQwfMeggkjzEPdfoAGx4Zvv/AAkyU9OImxEtzpm95gPgycr5/w3yMxy1NKa6WSf6h
gyw1FRDiQourZHJz9xYL3T4e07SUyYYWEPegHEfTrIqrQ0TIOcwX6HS8EUN07sRhDhVwoDnVOKor
zXgsX1GmALG7DFU6zatOzCX1QF49Qopm5SLT3vChjzGUL+mtgdad7aCxvmHimGWflYjVoKWVtsvV
nhu5HlBGkGArs8fTXcjBET6XG4T6YS6T+G4UjCe65d6+I/4D+z/7lFB9r4z9El5NPVeKD7K+MkbV
7HcoB6fi4tspkDR6x+L/py4K4Uo+eKpPRxjJxm9Pj2SUpjwBcjqfiDeX4c2wSsWNdDRDf61IGL9B
TRZBHbNYNVYcMdDnbHVQzFus9x3kSw/O4QzEZhrFkAcXfy42yWvG9BjzrBLoQ5ip3+qGWBjY/lyk
t36xELGgm13DpXomeAWprqDzjkwJCS8skP8FDKxx9E7yMNZ0CzdjuK/t90u8AT758pYBeopi25RG
+AkJ7YnthQ8/9YWs/KWn5YuuhStvCuwDGPvROksPIfKPorYOEq+Cq5H7TUV9oHCURso1rUuhjbDn
jX2Q5BGZGfa27vKMAh/kDa0Ir1Vl1TffAnBVn5ms66+sBHEEvsgSl896XpVHRw4kY+XMfBymKJQV
rAajTOU2OnNMNpArS9aoAsAE0YKkwM7ndJ3FtgOgVKpdDKW+1fkpJsGYTksiJ7bgp3A/APViG9ni
dmrDhV+q52NG5HFkXbJy9wd5a/mcfpgBjT8DO/C5B/y2y1Q+w2WMgBmhiUQ62rWX79/M1Q1PCKaL
21C5CE5Q125F9toIGs+HluckUlmePOTsegj5mBXCWHmmzBan2n9dmpFz4k14qLBYrIhX/3Eort0o
10sSV25/n2/NVyiHWACLnlAFIgEDcwIFCZvzqy4lzYsoGhlQtkA7Fd2z1eyQuyPeCGlIvz8umOJK
XJfGkhBLd4Nbe7vkl8wZS/Odm7FVRaGPikaJlf0MDiHB6TYa26RuJ4KbIUFpuisvnWGHx5FfFgpA
WrrrHUaoi8++eaqJqa0SZHnf0zBtkP0rpf+mGq2rbKmfCmidtth33mW/b9au0yYL00/z6PzMKDcL
qSTMjPznw7yL/1b+IY7VZYu2cCra5M+Cv51blhsvrIPeGc13TEp/iZo3/+HJd3jheAAgaZ24Am6N
Ylw5wZKADqUEQkXphJmoojGwHm0qPE37QeQApKKpY7WvJkNxCs9AAaxqVyMTZD/5j6ImiXFs6xve
g84b0HBKOLDktLRq37fy6KTungvxl3rZsGRE59+iKcs0N8AeHrDsSqfhKpnzMjK2/d7rrFw8mAsS
gwz8quko65NylQnjZ7o+tTIqt9URDQn1T1fM1B2g12/OVYjdWgbHwRxvLPNDvmBpjvl2+rBrlLGw
O04yVNumE7DdTX7aAJ8XWlyo9/XGGlGH2LekrT2utAs4kAvrq+OTbKqRSf0z+/9VcEL+hnbPzTyz
WjvhEZdVF8InOsAIe2l5kqXmmZRcRfdhd3lO6zWb8R84WwGpY8UzfV+Dswnl1BwTj1ClHYfs+hp2
lWZO3dzPdpAEi++XuKvz9Jvo+jPFCHWXudTVYHfLG1Kv0cFWPuoiC78Kr7ujl09xuZSe+lmPFkFs
a3gfWXVU3DnIxP8KgwSCccOm3kIMs5qU5eEEMhZotVsY1s0z2Nk25jeM7Bou4BFn7zr2AIpalDjw
I2uQ5hCvHIuoxL/lxeeVn39t07jxHDWQuHgKSZiFFCv2lr2NbjabHlCygYESMjbEBm2+wIyCPc3+
dQCKuN13Gx1yyKHWswmFqC9EwUq4kyjgYRNxBdB95EUBHcReRPrqXfuurHVcTX7sxoL6S1ZIJ17x
eyqtlsX+hSq87jH7eE1MWrzjosa+nB90qVp6OL6dPgmGo4wiNPucz6TOZHJMJBwL2HuAECQfxxOH
zf161eyrZ7Jt5GulVWW0o5ajFHTHpCJpx1Yo5C55rtCPed+zqvbloEVCeesl1ljymAWdomZGWrBP
8tA+w95AcEkP+KIlgXa8A2Jm4AwwiT71QFKtXDhXRin2uf9xLchu6jsc9fUisAhpUu260nQ8iq8W
EzwmEaCbXXQuCloiKUJqD+Br9MKcz9F0byEVFh8uOg1i1EsiBMfsEMjMWrUYm/zKBihttyXxhl/2
aaY4Nb9y452v1Bk1Zoj1ieWBFC7kPi+sdX9OTjCeGvojlLl+2OtDsJ98Oew3Q6S4DzgA7/5Nm/Fa
Wm4bkvyDVKWRB3PPMc5wYdyybj76k1QBQ4dYQqIELt9OXDODV8Y7xjcWriOtbPOejhEsIabAaJ6d
ofLNcJ2Rd+b7iEx5VadlYuMFU6CVRcOhHV5oQa0BJZsEfDMwQpMWUWT9IWd3xzKO41eILWycCBpy
qstkWZuRuxfsSj1RNaT9NLxFhy5VNphIDVIEtkzPo7m9Xgub1WPL9ZSm2VWBkTi4bqbrFN4AbkHE
ja05p2LfzpgB/qoa1r4kWRF5DKrOP0tQpeuToBD+++bt260jUf/e6Po83LsvlznvkOVHXAVMAxzX
jZadujIwe907cMFlrfmT3J2+dycSbBzlkqt6RX1wX7T0hkeDE8UvSE7JnEG3G9UDniQ5l+i/qEsK
V7wOgJDToyybU2LyrJ4Yh7OxhqZGeu/jhnMJ9jk+KRkk4xxVRW9nHJQurMgvl/KeOrBAafhp3o1b
atXvYLpQsm+2OgrSr58R8Aktvzqa5dIxhlS0lGX/ntuG+DxzWbcL0RKRuFsps3yqwrl/A8Emo8y8
/qpQzutTUnfZkDD34eBLMJkOFFScb+g5rnbmWVPSQInnBUAbtRHNwKcytMb1O39zC29xqR/ikFio
SsmFpbcf72QUQTaDxXykY1gX2d6BhYwIcM+sLFnj2G1r/aqTta04GAYwnOv296Tw/jeOKFaUPSQ1
+CMgNk+Kkn/O/P2KpRJ+LiM3Ur3kQslduqsyhQr3p5OszmHePh/seZivvwLKJFUGr5VYQhlBSin7
uyjRW2HjikR5JAX4J6i5ECXNGmKHYZdU16cJPH9cyMRFKBsvt5o3LjCaj/N5huseA6AxR3XaUsp4
9tjlDXvzZOi+a+bwxtQog+CYKZvVs7IYgnLy0XaKbwUgzSSnLKWLbR83u7KPHVOWMIgS5ypdJqga
OFK0dUXTb+YE7EqfYiRsnH9x0aPlg+F3EjHPbUNTYjD+MMfEcZ8OD/BMbhSYpFfRIsrCarh52BP0
2VNHi5HhlD9eZOF8ZA/8iQGYdfsSatVNA4+V9Mb9kQVyLOGSh8nvZKJS+qtxx0sgejr4s3PA0+zC
jNnBU7jtar0qe2FrZFIWQa5fQdXTLQ7I2fWMpz+L1ubV5OJiFEFbT/IE7Le9ccFYwh1VHd8oGB9l
PXaaxiDPAPEJyCDO18u+hmbdUBmGzWQqbb83cxIPh0NpwswnAx6bKbLPVajgVgVWkgJIq5pYDTme
v99zvI9IsvV+pzD5pM8DniW9B+PaU0xtKzRpQgP0h8626oyX/zmG4wxfwJoqfeYeXjR0wibktmgl
gXvq2Yk/7R2bbfIaHbAhl8bBdyzPiOhOQtmHcIHrHqwfSJ+g/fxHbs0rxABOhzmiwpsfYlrfA7Hp
N7y+yGKZOGxr7NYyAVEVVHr5xs6bA0nCCJzpHOOMWg67/CyR9J0Hh2dtl0uJga/J8avkyc0brdhO
gavDdFZTTzeCwZN3IDrFj1ilbMQTBiG/fkV0oo8gdFIxOXkvprfl5rXShTWiEqFwErCQe6DqlLQp
J7u4oQZIagFkPA0yIpsgwIFU8by4TERflDVwyT7ApxSaRhqwt91P7NwAHrUquM6J+08b7ELTN14Z
FioLSxwa37jZYH/iNcHPxmIRv/MQRwS/dkA8aT6dXI1763S8ZqG6a29nB1I/VqA18TCaH4aJU3zd
OBfPxQ+sxjWq2nFHVKJxANPIV7cc4Xj+OCmsOgILJcukzjwAHhJe/KYLJbm/F+/s9DI4XyuVpSIv
8G9AQrzJ1G5h0D5n/blXiHdV+p3kLTAd+2oyFE8+NJ9/hfzwqN8tyUSxrfZsm/dtHE99QwX5MoLa
m3aV6jzTWBBbfIUIUjxgKWTcVOCJ49biGxK9FRVpVf/du5whw0B73JG6fSXAHPmGn5DJ0jY9v9nR
1QkC/U/PZ862x+6tqN4w6HTqr4W9i7wOD/K2QEJ9UMLhyYeOIW8WuesfZDf6+/bJTFIUDIeOwwSx
pfW3wi/PYsb72BOMF1BfPF5QZlrfSTAr6u1UfdEY+YfiVzZkJ8Y3DUdmTyq+KMMyvauk77jb94Es
asghXn013sECL5wK44q4uybmPnr8V7rbT3CwvhjYIrRbiVY9y5tfATn3cgk+TTJBQ5RaxAQU3oNA
9D+6GR6ZzM6cAnaWOffUoYAgboqv40NG3CD3z3xgRV0TQphe6ldDR1IWvEiiaPzdF40nXnmI6RvU
dNJlqKX3UakUSeClpT6DBOZZ2c4Q+ge4GIEjQj653ncCB2XwvpNcxOnKuEWLdeP16DCuofNjaDHC
utGGV97mUtiHHiJ/yKwOvG+r95eiy+XzSE9WwSKu9gRE5/whY64dBMnv3XbJy9fyQiku4l13z2mv
VkfrL1kXMfIsGp3dzMx15fOA9xkzbdTs1T/+BGcKdWngok2t/AX1v+KzWNBONdrz3zhWRVH6fa6b
feAE2i7UsK77LKAekcn+0UQ9HWEczQecQzm9B2v9gomJyrsEKDdJ/hboQevgmw0kKaMXQNxNKLD5
ZCxDa1HU5CKXMQsVADuHof16OQnpqYGGJdmoz3iDPIPUHtmrjBykdz+8gQM/tgKClEo2+nq6oxkT
rL6wwnBbdiSCSwDvmnFZMU7eK49pBP7PNtStYV6VeU2o2sQmTfceBo6xvzxDFqHVhTcNEZPFJEWG
rJZIc/rZaSAOhAyb76m8KJMS9l07J8v5rEsTOY69EBKGpalYBuks1r06IQqM3CK3wV+RIdCQZiaF
xMgzlAit464k9fgXRxdq/OwBMILtEiovHZGGGW9LCUwU9UzAoUGsGtxhPMG7JwD+sXik4bPcazDx
M2aRPiww6q+0QC7WYbzvzQvl4bYgMezVu9GZXo8k5bcX6JJozi+e19Kjot67wxXYTbn+Uat/3S1J
fyZmBMbnri2aBx8pN/lp8bPHqVJf3X/eVjrQ9JCchRErPtfyNwwBqeGKCIH7Lm2YJn95UIuMcTlV
//xjeC6e76wAZnlQId/0jKjArNPGHMixLkePzWHm4mJaLCkQyVBvJSDLtst5fBrD2EkHvqSai3N7
UkZQ9Ee33ggjhgUUhNPy1GkGnA1I+tf389uPl1iXu6LuiyZlcEknk/TOanSkvrS5B7rMUH3p/Dm3
Ni8guPuNnES3lpoetW6o5bTxVwR7G7XHtTyIL58kGCxMuiJ2CsDBfk/68xq+hX++/TfAWPgUS69V
ir5ZEMchL8gjNhOKDwEi3FhFdVUTNcYLY70q8vhmA0hdt/tmHCr2GMij0Fxre6348aserSA59Nfw
0nk6w/ixRNPFRUWfw74A/K8+bVAASRgzOOjadWayvUlFB60kVaZjyyGJ0BoYpQb5JnLWO5hLxYrw
RuNzsW1ScEaFjytZiTRZ2YU4vcpHDvP9ODObc7mPnukpqY6lsqED8ab50p20BgvxO78vJ4LSX/On
PyQ+HMwJ69F/fat0CSXHbp/cw5myhtXjvkbU8cnKRsUtvJTIvDdaeW4Hqeewkfs7+OQb/14ss9pF
gLDI/4P03q4CDoHOIt9RmuPu+FO9hcMpGRHmpj4DsJ8FUcOvd9hPKiJtC4vMGMfITZg9A2sTVwnb
1OLhRY7POeFwuN3nj/gUp1i1sRr+/HJfJL4O79vmrjSb1r8THQJgPtMLrVvg8jcKeeR6f4PQqhhM
Ul/pFbZSDEkF96UFEpLFld++9g7+TEgwguKc24lEGreDXdcBB3PXn1ol3xZSWYw2LGteKjwVVuMr
eLv+bd4XbmsnCRiZ5SI6cZQEtLWQjMBmabyUtk2w9s402QINF5YzElwp99S9EziT1YA1iMpejeKE
sndqNbrJ+op0absk4ZYFtBPrw0us+vjqjz3DSReVP6GYAlFBF9yl3lJbwcm/6XOOUuqTT9W+gx+a
DRhhyJgrYt1pYwS+fPza/88RBUHHWNBP/+8yic2o2AVqd8OW2dKVhpOPp9BLLmMuNYzmlt3zgRtK
b32fVoVgSWBwklAxHyZo0XM72Lj3P56KmrJuswH6y5lexafhjv2/yn++1r9NaxA2UtRoUWWxuHen
oB16c7eBCa0PpLUeQgXd36LVbZD7Q/L8rVuQ0TTGeALl8sycs3pATy0j8psIAOPQxefH1T0x0pr1
5bfcsoxxxd6QRCJUZe+LMDBcFJoALKg2x1Itb/BahQnEzezGUnhCgxzvEYJVzmTXl3woQa2o5ybM
dJOfSlmX2/VGKoX7/4hWoDny1i4V0njpmG4k56sQpvGINRu/Q4AYN6hAHMvaZEbRMJRm/50qkjxX
1iqQ5o4IWHlj5bk1UrTSV97aEUaVvrIF5ofyffovtkr0g78nYaZlHTTBWC7aEBLXeJpOY6/Ar4zJ
H7F+MHBckKwx+7rcY96AvYz/adKj1X+HW+C+Uudtpz4HL5npxO5iOdbixM1DkIEVmDvysF4UcEKk
mMxw9M87gqmYdmII+NfjiRGzgBbr6TK9dJzbxPMJdaTkJ1LpIpNd2o4pSWJWwgGDd/jkphDysnvS
mnDH0bu1A6yTrR70hcCt6XyhOInCopVQqf/V2vwFajtQuWEfPBsH8i7y3h3AFAB1eZMnHIJatTrp
ApYWgLydOGqXyI1HSCnF29rOQB4pPer1/ifcevfuurC9T84ikN+j05ZP1I9hyItPlA4/jSl3WWEX
XWFnkfwguap/KnTDUxqfAGDLqJ0L1aPXMJIxvLQAzDIuSXoka/iE9sPBI9Drsfp5OedRW8Gm2Fqw
s3h5fsgLAXWR6un13zosn0LHiKMWxG1v9VlBSUa/FXx64v7ciLtSBNgWt4/wO+pp9VpN/tV64OKD
JVUmYfhypDhcpIprLZ57Dwcf2R0rhql42jgCz06jXvuKHudOkbAW1sValrEIHs2rpNLcPd+SOYbP
coAPX66DoqykKmFXPHFL3VuJblrYAD7hv87tMP32LsFshyrVvbos7W+kQnUE71+OTme7TcsipR0i
KUYRwnA5lLrlX+r5OwVq+xqZXNwDub7b/Uhhwh+eEQhQdFSnNwjmF/O+J9+uiIeW1n9uF7KH/ht6
F5MjFs28c9gGGn3HQZUIwrKjnVHLlu1xE4iVDOlxQQNDnhfm+yqjNADwBOLwfIoZHU/vhwXfZoJj
PFXppSHq4BjXkAXWHGYU3M0l4E1HrVXaBjJpJCpkTPfP8v8VC6LWXQ2ANYO7HWKrMC8HxEEdhMTl
Gsqk35QKrh92lZSbiWtn/D3q+cvCrkig2f6oz19441FZiIDmafAW7FhSWGX0mXvWnRcLdT5h4LJ7
yadFS6hrJ4xb+5RCY2cInBCbN+IJVdb6926Tv6gs+oFdem27wIvVFYIhIExfOnW6QMW5QywFTEi7
ruG4IlP/QoD6j6FGcp+3NW6yZObLLiMxSgOsYTcLoKonyGJvZGdNvXujRqtneFSaI8ONOfu5GBzk
CccATAaRWCBLFixmifqH7Qf1ayGBMC9knCQUcJ3V24UZ+c7MgB10dX7jqDKZ2GVT/DOrzkcUP9Rz
RyhxysO3WiaBxjVJ2kOAlVduNKxzp4n6C7AsULKE3hv4vi37QjM0gUy3MNqUbax6/sO048Q9J9q9
RLUxR56ke7+tj8ekgbtGB9NbchzGKypOlIxY/ERfjeyEUK2uaWYAD26og2mwyhQE1kvcOjNgkzSL
FwYw+lj81C+K8XvVcDwBi03r0xjmbnbp0OFkduo8ehRpU/49UNJrkoMRG72W5FMdyeXGibb+ElL6
qxoTb22VMnYo1LFbY4CzoOFL13534B9qoZSVoLhoq+nbi0ys5dQ5QkLlvn54i9pNQz+8aPUS+ILT
yU2Fybmt5FwuS7uvA2lRdJYf4tcTzWWOMeNApCu1MMYb1snj7oTbHnrkclnK6ACrxjMRmTO9Qevk
hWFjO8ARjewPQs0dPAwL5RsvwTeacQUg57/aBpnXWR5Vl1N0cmYcpA/pH6NbUf8QXGsXucf1TT1F
RIgVFj7fTSGqwO1dGF91nMo0CIry0quzO/PzjLtv1tr4T4EPd80J0Q4qOBCBId1P+/5+pu20iORa
ekLVQv/Go/RoO+HCzq+33IuUOcUlybgz87Ymasucz63JrtFkMye4VNNwpeiGjVxC06HTW+wMVL1E
83/EX+Mj6u6tXp8RF+bS3UYwHG6cNVwaAVl5f3WviDhhQBIatL2Qzg2RG+rN2uYBQ1rb3V6+cfAp
TzLL6Qw8gQ5AlzJZNhf2esINH5Eq8GgZ7ms0j+vaAHgfxSnNnPhrWGHu0PFfPvt3gOQlCvUZa6I8
WX/0JGrssugfhhHKhXTjNx7o+qgHoyI9VkP5eGfl+pWhf05PDz+/tkkaZVPzTsWmPVh6myU7MH+Y
ltUy2aeuNKXGvjkCJiV4x7maQROjN8ulgsvqDng9NsG1+5Mqd+ItiS/VQ8ACGrU5mKtJQr1eACeh
Ad2ObuT0zQ+93eKHwZ5FN78MknFE22tsbeuTM1PS6bPltQNkCIEVfFx2V170nvg+FDm8w9d9S6XZ
p44YomEdKz3W//nJ1IWNoy7QGRoprpupmmGCug8q0so85e3Zvyf0QLrvgZ+niF/5e91y0I9L/cHt
h2pX/jjOAxuuG3TJQ9dCntiRgqjPQSCgo+ztwL3NdXDK8RYPpfukD4Fm0ZWA8qfl0YvzPMciaHz6
gr8DGcLSBb6tWQkDA277vgscnvHo89OhREk+MxnGIsFItYr9nj6GtYZ8s5ZrlP6o1Zck+94GTCmi
rtlbrAPfFyohrAaV+S0VbycEILtAZG/0nBDGOsTNCPDVNa2+h6zc7mvc8QrK8h5lsVZitndKKolw
dBdok0Ynxbi5O8uI9tCnnWtHNTTpzYqR23tVX6bOp5r5VhJFjcSJSgLeDMLa3O3TaN+rD3/RLt5v
mO3GKC1wDbYdtPniVio/aWJ5MMFTYF3im/HdrDV6kXqVjosG0qca6udSmwvLP8VBV0uf3yKrDmxD
moVepGhDYNQPygTtM/9WJRDNv3jG8VAxNhEuQ671b0HmLwaQxhxvyX6N6sC+2TUTCbm9XFS5bnMF
MfJXGnx+tcay9H7OR0eRfho++qL9E5iosFKOf3ySoCF5i54/MEL/2VdAsjsMlgopmsyveEtosEir
MFTPz+HkrMmZRPHXnaEWTFr2ylQyf1m062vkpaPdEAuuV8rEBY09O1NOAK3L7JPOQiAFdDgD13QF
U/J+xlnRCqb7+RnwhusIyipcodEtWmlub66xHdSPTijBNNEWGbHevqPSNR7NPKwW1QDM3F2iDXyI
wGlBkhBESVnvcuo5fMLXHQs/WnEHyNCttG4khfbgwWt2BXVEvebTTANhkBFZvfuoYzkdeagqpxZS
ft+JMDd4Heo6+DOa0xJOhTyV1enh+9oyrpbSeHlLfSgIM85xntxrb0wspPoRxrizMWVp7Prfos3/
as267vkkkvm1ue1LCIKfiHfIE64ViKPY5O4ZfYgZ+hu28JaPVHK4WZ237r/7V3iwPKiKbzRVWJl1
FidMykdomFMbwkLP9zTM57aTe7Wm/FqVecQ9gDJkyeBgtLeg0MAlYjrL6qs6SkWwfn09bfn80z0A
hZ9MTpZPC4mSP0Pl2HNs+7fYSWt/qXydD3OHH/33qC7AAT6DUL+e8ulrSXSXbgn2/fvA/CTHXNgl
8kbH+3Zes9O0+9W1FXs8b3LTL1zjR0QMQPaW5+mdb8R6g0IowGE/+UPfNuu1vj0bpJbsmt1PtEgG
Iwww20Ctgs6SWD5dOi3Cd90m0XJ7mRn409iT8mdMDeQYwDGvaKiG7VkVcCYR5NJvchcoA1si0ZPU
c0w6ySr8KrOqnt8mckAz7ZzztTzzHBhNxGeSXjQ97Qljn4v/udVBg5xV/UhAN6wsDiDr+cPz4QBu
HaJdt2XUYb+Rm1nqiF66MDj41ohaM8O0rT8Fe8hPuytQ9ImcOVLpu8URfAeZ5J8X7lFCtu4Na75z
c6HHSUDcd3TegVie2JUBxFvoYUGANOTo2Yg94xuqYD9IKONWy9+6KlQFUo40LjFRGLYR2JKLa9SR
TZh3j+f3qRB0Jrx0Q3uOJJV7O93kR8+3Oto8qBHkdWvrbqyuXPQepdbpXpWqbFoibjNOsTLiwWPM
VhRTyEXgx3dziJujTprK7JkftE8FghzVaiYjmLfgMU3DcP3nr5NdAsE3R93JirK0ma61YpgUmxN/
ukhIbkNQL8TL5hVMYDn7NQ9Bg7TLQleaXcTpBazo6yfgxRReER5YnS7zrCc83fYOTmM98bbjpxtP
5SUfVBdxrCc+kah5V70U8OW5/gV40H1hCaZgjW3+67mxHrDgVEAlWKIJURH49ExKnaFOyEZxGeM2
9IoIOJT0MuM1lqAzyKyppUdodaPwaieGqAtQp/lIFZ+Ng7FOhZ+IISJi2Sz62iaff5caSvM2mOUD
jOrd/WTjisfFoin5P9CblK/JeJV/3ATBmRcInFqg6oxTKBPuQM+jIzcc4V74p9l01XIQlPzhB4+W
eUXAY0sR+FzVV36dYUO8Se+EUCh5GGtLR5axe3tQ8VV9l6fkJuL38heHwxqWjrAnR3JpxyefECt8
R3/7lZmbuTqSrxjhIsqKqXQKo//x+kprWs795x8yiwHrjHZseUSwT1Kr//lodGt8FK7VhJ+sk/Z7
2ERbghPnw9ntggMlGiES3cIAbfyQDP8mh6dH8BIsL6qMyx70VHUXkWpmacPBJ5qPIpUBFgLLei4x
5mj7k5fNFWDnmjNQAn5y3Yk/uRE4x0IC6wGhEU3nsqsvtg1Q/7gH3DjfcyEu0+Oc/5YVMBd660d9
NCjPeIlw+0tDfQnb27g5yGh4T9dlo6IBBqAYfyg5GDpv8dokgveo8ual+YkuWxqgP/CUufKy5bgj
xONMsWcRDtDqz0SNccS3clKgJ/QzN4F3BObK4s3N5i4LiCJ0WWYMB0Rkk9iM4sHXp6PmXri9/y9P
Z3UCYcutdiP7Fu3wMj5eYnBasdaf+zGdG5Es7KGtHsKud4miZiv/zAlXyOvSLQaHBiPLa35hQD+H
zSjLYzyRJ+3fCIrBmnPCcrHVcHtlExC/tFmEu/2ywyou85URNKBP/ud8NCtH3bqbVtWkYVGmsWRW
Dfo5eUc5SvZxp2GsUNhUvFGwWkIO3GOrqCIiImFoxbetbIk15t57sW9xIUzPGHUnRQd+P4ee7VMu
sxb/d0Szw++6ejI1kqZX/aQHFO4cd5BjBHzUSxgzyWIXdg/u0gqr/6uGTTvt1glhQ6R8vUAmV+IT
SCuFIwO1YJbfobfknQbWb885TJY4NfZqcDRZxFil7C99SGiGe/pPlK4abv1xiFaYOuZHkKruEKFX
NIAwwWHQgszIlr0bRSQa7SNhFmcbCF/olFAgFOuxt1w8Arim0a992zhtivyVlwRX39/jnd0YqDtw
6KZTjzbpHp8MNAisOWK1bj4ZGeanjZZj+R4vkcCEoTOloTOvwcDMHztl10P6T26Lutz1b5Z/7DEa
4sC5IfzdJ0kILSEeZZXwqATIOdfuT4YusBFEUAw3M/DYzi6gyzNuevEeJ5uAnHuETj/HYTGuF6ah
esW5Ax3VX37B2qIC2Ye3i8+Yz/h+3PZ6tvcceultyezIOcLwEdc5qpVusd3SCSNiR9QJOD9bm5QJ
8J/qonLKAoMrZA6wGSTRMY9PgQIR1N5ojDxXQrZ+MgDzaFt6JYluTZUloPhYKlEOPYXYdOOO9toY
QlXX9QPZ+aYxCKeXueit3t8qzIBUkSnjHAIcA3WFEixzX/ezaVioshmAab7xWlvJcHqa4/PCYZQw
ExHO1JwwfqL/xrj2x3nuUyvvIYKR8fsL98KsB8k5jWAAvsGzXPRP13oKBPPfU2KM50XNu6YEu4wl
LLcxrASVP8hswRhL0nQo6kKdfX7w4YJ3hMZegiAVFy/585G2qaU6cmlU0epKoObQBFovAiWebV/0
/nSO9WehADFOxUoHljYBTr7MfLoOz/UFqaLUVmT4LCUol7j8i+Osqd0VtjqR5dONzbDRY0zaW89B
x+R10TrpV48iyYKqn4fqKULc5PpA7wuNxR7xLxv3f1vLVG2kdvo1zoW5cEK4suMznZTYPGCGJrGd
OXgPkarQ0jKO/ajBk/+b4DDUxoQq5US4M7eEfIffcgPMZJUU3wvggUkw8kMnA8d5KFDmzj3h6Ru+
g8X6Mhe35hK6h8uqQPw+KNgiobaWldpmUWB8KSbWFLqSRDAsDomam1COVU7eFJeAXM8LAfi2i7zs
KF2ekM70oS4ubVfd548mroxAPj4rXiqQh8ISzsVm6YRtPx//T08rrMA8rJ0R8AmMFpTh/MlmnoUT
2zSbdzQUaGgOcRPRULcXeQ55Vsj90TRy5dLM5sXh2oXuu2y/9HuGy6tMTf/+PPAyYBK6E6XZUheu
D7GauyxXBDZ6IkJpoR1+uTnQhrsu6p1UZiZXTyGxghq3iD72S2S2Q/rMEcOX2HWat/o/OLD+xUA6
pjHU792LPgjruKPHE0LMUBvhROPfQva6SLAtU0juirH4YCk/rHooyNJoJXGvLdaFYARxrVQqQQlR
SllFvGX87okar6e44gQ6MdpXc9TLBQd5dYCow602NgFmv86WQykJDeroBHztOa2QEIAI5GlnEkH8
WVzkiTYovRU3TEFzXJqAclZue/VbZFFXkvo1A77JV0RU0hlm3IznAmfzJNqgYRBe9od7zZPu29K8
ydLWAEAWEddsX9mFiapBNw1uGcMBztz6DQd79OsTQnq5zqYgMr5ACX00IP1frNE0FLodhPjysmqK
/bjiTo+lc/JZAXiNDDjJNyrBHbSn369ZjYmC2vjQW7la5UuKpbKl3UcpWJ1M8aYPW2hym6zPDJ3u
lj0lz5JzRa2xFof6rx8gA1gO36w9r2Z4kFWhRj+rMubrSiGzdd+hvxwRC41omi+onlny71NGSFNC
YTxe4IXI80fffnwmGOgvRn+i3nRLia8xqQvhnDFiTTtS/b245IvKhkrYSQGc2k6CGxkeIcGC61Bl
gNAoV1dxQNxhSu+/FTiHIYXIIQNe59hRlpzzfmk5e0k93xR7PKrSgFH1mZxMcRQBQI+3PVEyu7Hh
lvdFfgx3wXUp3tEXXu4uKNgpT50iVPiDGngWQLXGTv5toOKr33U0GxOuclxwNSDR1J6cEIUw89z+
zLMglGoREWv44PSBOCg+e9GdqeaTR1vhdo1ppYXN+A7huILZ3D/1gVjyngvXj6w198vTpmFCHpsS
KdFqlg5Azu1v3WwqoZKV9IwYIgSEhHwjwcFbI+vCXutbQiMU1xYk8euruGzX8tWASlx/1MxeNwr9
bOnmJpbzN6S7pFaiBtEvCFkyweWJwYh4BlSv8wASKlvhBc+Oe6aRCiJe4iUbMi6ijlAz2Xer4gXR
nRuNf0ZchWQ/AEX1RWcUoTXjcL2JHgM94vVVmbwcBYyh4E2NRyP40OjjpzWJ5snA5NbXj8EBeNcv
u+IyywE7xU/aim4WVIfiLGy1Sv91V5q3fpku9XyFWBo/ZDVdCuu9hMbU0dhwc4W2m4WuQgc1scxo
Vzr7voR/8k8tY8bEYa9kf4hx029Hf6ULCb8odke4tpekQDHfI3dkpxrpLPTHsHRQHlMaCe+Fk+7t
OEkYVFeOD9RKgLoqkkFRmW6ElMAg9brEqamyCBkx05c8jBJdK8opVjr6tUhKTQR98tTs8OIlxskk
Bz/tcFVoZ1chLqHltOCKfp6lw637QBwdn5DqgwNRga6pw4JvjP1BZTOzXSaYvDs5kaRK46ik9Tew
g38y98LsJVKl5phoSjEGoTx2fCHCYpkM7QKYqacYIbwNjESk5CzBEu6GEYp2oHuTy9HW1vT5ySd2
Artc7FH+7H7+IJMqQZJLIsJ4DuxoKOKVKmpgGamxcs9iCHsBOhA0P8U/NU01xBB1er3iGcSUVtXa
V1HKIMg7ru0KnderCdvixN4DrpNzuv48o//usZGPIUZeKJ3E7NkpZ74319vSb0mIdtArC9mIyskO
JGD3u5u5RxWF7jMQ5KHXxry1yRYPKgWFReqnpzVqKfoRC8T4zj1d6AKJkSbN6LggbnT1w0ztmnvs
NY6InQvSk59GDGoxorpGmqfFTEcLKAEZcZdQMm5XAZUHDKYXyMsGRz1ZLYWSuzlylvPYQMOVns09
WUv7yBVpyYeY8KmnxJiqhitHGyGZEDYTeDY7L9sAAiZAp57kcvUAo1hl1YEPLQ+foUkv1VTR07cI
WQ255+WfNtgLu0Qq0RG6n6AKJrr4OPryGxH4+seeYgdwMtbzWyLydnlzPTAIGo/3zVAyz6j+tG2G
D1Yhm3jJn/gSztzn8GAIVox1omOLe+ceXTrysOpGRr9J8nb7qj1Gpe6ZDNzL92NXACPjYJWHeNp8
9WUpBvISCU3q5TaU64x2aZBkGKCiCkEH7t3S5vzyAR+u+Aeepnrpc9rI2mFuGp8h13hkjdDt4TIm
Vj43sNUpGblQ5Fk7PbPyReBcO6o7Uvau3GDwLLhCqMQFExSxvC66O3atyZfTJtMq4qcQK5iZCK1k
vtjbWmNOoeQVqIkQlo3D9tk61fa4nT6zmvhA52dcj15A1eOXYT1K0D+pvVXHktfhozPi03MD6Tvm
k/mC+IH3yweUOASBab8qrFBrEgWppUjXDIoS5cBZtK1yjxug/2CwIq1MWCy7ViZpdortwhpSncdn
7rGnFtEOFqbDPhvPlGh45QicNaQEtZVfUP+KU/uB4AeO8jfyyARTgXPkdZnoofRvCEFBDHzrmKic
mQLyZRzDMAXqSZhqBPEIvGqFQxzSkhvOoYcI69UD4MruhC6tbymGSMc5nsivYMWPbzJ73/xoYXd9
E8WuiCzGk71QiqEtTV0GqLB1KnglciyGVrKyawfk+JxXz/Su/rZ4L6jdDeM4x26+j/FEJZ+XnvOi
LAIzekkTnRnwJnTvKKjBemhKRRMCTOZgF1Njtygm7mx3esjYC99dstp0z/1Ydk80yoMSmIdmj+tj
kw66Ovi9pzKgrDEaHat2guy2CZS9Za4VES4ITekdNbaqI65WTmhUlDVNDojZ+d9XFYucL1igISmc
Y5I+ECgnzV2uVjMF6SfGbX6z/RWh+gUaaoJ91XlHx7Hw0E7wt6NQNBCXunLsc29L4WO25CkUUkN2
i5XVR/QXvFwn1o5gDDf3qhOZnJetuOBm3cIqYJUasSMfshMke4Y+b99SM+qTEQXGVHglmhG8rqKJ
D3Jz4YOnK9ILmn0PkpgypBt+/S8NBewbb3QvFiLS8KfGgm7kmWhBT+9pCfX38+/tqPjVJlpVH5hU
LmumW60rM9YlL265m4DJyz7BhCE+wbbcCwv1ve+ZEcGwNz/0qaG2lcO5Jhtpw5uBQgU9vkObh+kk
pOvsI533hcv1VD30l/gNRhz/sYDVorin8xT6Ce3Wz2xDRsFljt66YgCObgm8iVj6/1+Me2lvg+pw
Sm5224rCzoKT7DxaPTzAiHmn8X8nkuUi1ZXMEPrGRoTVE8gM5ilYzTpFncsNlqsedhafTaoXYqHj
vbwk33kpytQ3KDOcI6tGEvwfFzapDKgamKSYc3FALp6At0bLkXzANB5EIHeGokPRgxJWDfD0ZWUB
azLff5f6CGj2hOVXC3R6reGtW9SykYAQ1Z/cJT1K8Gev3DZSk22Ue9CPz8KotEXT1CIkm9mtlgwp
QJViZ0jQWxt4blhfZiyESgNPmjgzn3TSapzjViFI/0SwQQSHdRqM386QsCsq9+HChbBvFAMTIWVg
FtIVamxIRtudxHAoOL5tj3p2xineUe1KC9i7SUvMB/7vadXSeIZu5nNlc8ajo9yLCbg4BS7gcxzR
jZNoIO7oM0O7YIZ9mqfobu5ILtlaVJcZ00BYIyKbGfKk7lS0OiEbQFX3hlUcLrMVGp6PGwiChN8O
gEEIFgFNM6/V9Je5HS9HMxSPAAMf5mqzI1gCOC8hbmBKYWVXzi4pjAmrxdOQRdsRECAilM/BWgvP
sHLZ40/408FLDDqBY+DbSfJLudEoA8x7yxWogbZNUE3AFI0XnKi/aKVAuL2IfgljqlZllUjghBiK
dw6yoLgb82xX04JYMEw9lxk5jl7Yw1sPmzir+vhsrB2yUK5JU6JOvXJPb1SENy8ZXdrmQRN73P0k
bxjmzEByNqDSGhmuHbSNAWXGvY5ovxK/rAERUiTJudwpFxGiuURB2E3rxr1Td/oIIwtuPXTW5gV8
DQsRPkfNxwXNFdd9qBpVNgALsxOUc5QJc52YcuMiX0el2A3QX/zxnVfxDLTzNxQPHSouTfsW6IZs
HuonCDT4FXud27Jk39r+pjzkHo0hgY47DIXvM/uaCWuER+WpOZCrjUfdpQ0vzJ9fDzpnMoQByI4q
trM+hV/Be2tw7pVv8dNX5fF33kyrTYZWI3LwyMWB+7F5j0mExqMYfJdquPbfEnME6l4sO6Gjf6U4
kRtcPg2utjqRghN8UJxnjBQZ/KQ8WkciG3nLcBDEOREP1UWD3trguRjL4o1Zep4t1LwfNaqZt8a6
XhSySJnJ0/NRZ48sMNGB7qQqlZ+sI6JqRw+xuPZ2UvRW6NqdNB9ZB5TTFCiUGUqwZibzqYe5JH51
5Dq4L8E8yl7ZMBBUIKWmty68SlzS/TYU9cEm9GF0f25ia9Qd6WKIwGLgo8eJHw059+zHfO39C0dd
r9WOhHlqA8IvXiMF4Q5r75hUg2OYWQiqkG/v8ZYiYY+8PNSO6Rbfj2qBMSZ4sH2m6e23OXEnnYVi
ETyT+M2tsg6TNm5gO8yU8s/fPMaY58YS//6ot5b4bGC0Gb164OTzsWB/yH3L63HfHnLHVV7NsrZa
5MRrcX9icE6ocOBSAvgfTWPoj/ag2EKpKEkrk6AAHfgjnwueTWaqR5xY61hTGDr1VzP1EuKIhRv3
Axpr9f1hvUaSf2zTxXermKhz9vUqtF5UnZ+ztX2zbLIDBwr6zhoDXbSX4QAlU1EaEG2kZESbSJkq
K52IQlw7/+pusEu3b/+XOmKFrlJE9BDtHkA6c0C/ZrcnXMzImA34hV2ZcjKKX8oKH00/LoK2nUzq
FSEVdIcJvQ4wfW0zeSlSrEG1U0QbR8vw4d8rgleEisySdZFLYHf/kMgsBs2cHNdFX/ui07pgpSdW
mBHQtTEcBuIduEISaGBqXkNbJj+zAG6bO2H8l2/rhpFBxbTuK0GIUXtRNZP7JElRF5oWlzYG1Zva
QsimRDzFDm5PBJ7YtSw8MD/edPsDqPgZOj7eg8SMg30KnIJ7M8tfZWih+2YeBGARlKAIUB7rAhtr
oZIH0KQLfVdXdG3QEWyljcWTCUO/r8VTA4eQ305t/M52Wf+Te2ocfXazgcCGif0+12Iw4ogb1eoK
n2DAlDY85K19c/TENa18meEAHVfw8j/N9TqklW3AcGAj+8suVyR/wM/czvU6cHPZKq+wlv8gksFK
QqoE38pU+Npr1XWfT1vmLVCDY/JStQA1mffMPqGpBYR8v3rpguThIfpkhjwA/K0fgtBmkA3blYW0
CrM0QxcGXhqUiSNXfAb62d3wgvwWyLxPoD++jFsQMiYOTM2ylTVadzcVkueZimbHALU3DtaH/lXc
D+Vob2CjRF0VpkOMhiVI2cT4mMIa71ceoo/n72ILhFQhEKhn6bh8Vy/FvVmhc5Idxp9qMcK7G04z
CSPvcHJZ6nFwCM96Y7jf7IJgZCdA8EuJe+nezv0mrfTlt0Ec8uqtLDyVCPs/0sl/PjqSY6j+22bU
Jkniexc/bQVQqtj+udNcyqf8FlTSi/FfZ7jTfmVPTEPm5fqSRVX8AnubqzvrKkt0zzCa1pFKFZyt
Roxb4L/SfewBPiRtb9ImS1XzQLniLChTJU6hX/v0xwYqqYE+knlsd3H2SVIKtpuWUQyGNiWm437T
fQusrzNrzl4iXzbVhxr4PflAG1s7yU5YAKlx7dOFm9JrRkee5DEQbzKSGpX7nTtVN1eUi5mQc2eQ
TA2tcwPPYWBmp6fFpsyl0n0fjywCrxKUSSOfpp3rK3htRwkuYjG3phLEQvpS0rhA6TIrhsIbKrWk
jOqSwzE1NpJwQSkx6v8SpMzjhAVda7jEFsw3TStHW1xNK4b0FTaGo+ZuwVOS42V8Et+650ioPJF+
OxFSDa0TEGvJxVDGt63x5I77GPDQ9VW02OCmSR7X0sMYIvAQ14Tjl23NcA9JBoqZ+u3g0IDT7/w1
YeU5SyGgc9wq9Lf3FpTFpXox6/1ZsAipQcZgT/6hLo8nZcJWtDjCme72TBeOUYrU4USmoSuf/XLe
R9LiNrHc1eRKWtb2zXwUj/mpx2MM3dIJQ920Cc7cNDanl1KQVIb8Cw0MtucWFcC+2oeLn+HyZzWF
hjZvMjG4Gke1K5bPObLfKPHHDtegp9QgX2zLfdQBF6khf4HaHVwVLjc9XEv5BKVML7WsEMVclevJ
UkE4jeqv1669LRLsXZRM1pxwcm7A1LcM6j6R9YMhmeqVhFTks7A8q1iOGxUL8KHwFE2IeC1c9u/V
9fFi7c7djOoxF2rlVYwvIRWFd9ON5F04/uqlgzibT9ojnpRyk81+PyeDQ1dEtvBgtwpwG1lTSUu9
eNm3qiYWYgkknjj7ImcGSxfOmRZ1xL8+syLX+0cQ9ghOfYs11+M9kn5uWF7LHhGwdTVX27sDh9QY
F4xq6hlsgreYxi/cP/PSMRaVb0K6wENQXOUv8xHTZf3FkLhv9IX2sU9s+/wp5IJCIH2UJZGGoECt
DhPj0Bsfl5szILCbBQZR2UGl8vijcf/Eue7oDM54njyPsOLpvwqTfXb6GAglsOGaVAcQa+UzVfN8
NfO8hZDfr3jhJNmeDTFH1a66VPMkbfVfzQKaEzvtKgQKBOKu+hUtIFDg40yXkYH/fFqqkTMEKg1k
nRfchxJ+KbHerHdDg4kzQssbCbepU/edGQkUEQoNh71A0vd5ybZFc7FWT7F9CXFgPn4c5q8c3pu6
buvjedWasuGn1QLhZGfiiIHcnlxm9SrIHazbxGccdbZmiuBEgX1KI+t8OhiV4oBdl0F1MRleAumA
UoOGbUFrR3lpEf1iug1VbVZenvrtCIYGBVbnqNkC+tXkta9QQl7Jy2rw7Itj8+hB7w4H28Ge2gph
k+guzLRLni5SnldasyS+uwrXR8VYnQ6YUOE9O/tVHhVto+PJm+9BXkoR/6bRaMN3jvmHqHtw7DMY
2DKouRm94TIwmLVqrwldQ7wd7w490LYhCIxXOBnPEVkW64h0hB/lxsBFbP9fcCUMQmp61CXC0AKK
4kdeXQ+yNpVsbgwr1kMmPlgWW/B0b5QDnpgWLUZxaKQgjROpllHL8Wt4RlcyIJ9yPWQ7PLiS7Gro
17vN87n2oOBAAl71TnpB8+TUpDSdBWx2phclWhTQRX0SjmV5l+kQquBf/kib+KeH3ExZuoIOC44s
y97BkApXdOilJJF1JoB7P1hr71P6av+jQSTgvCV5q/mznD0j7j/IF+qCk3aK1V41/cGMi+TUVkut
EjklOceAVLn76h1MuFtKb0UcP2nZ2n6yUB1Qrsbyx6gquT+hcGthvhkXCrpY0wY2c6sKTH6Jrpkb
a7bvY/D7HAYh1Yf4zeapS6HC64LfFpBh0pk4RyIK6CAvFx+aJNK1XeQ8+mXmomUSftr1vmmx2ZOX
I2/gCVZV7K7SMvurPE7RMvhILkEsbE5akGn3lRE/pQCsHNF2ZDahvSw6cX8RIjitYxUL31558wS1
WZmEl4wvBzeesnhKW5IEaaiu127IQ8dE6EvsCh9Q18dUodJcdBNUuoMI8SEpzsuutk0PXnNkGpjY
N4s7bTmdkXtI2nvtEHKv/gvxQNlvUoCFCLD/fxUfZJJ19l+Icr4B7I0lcM34RwpIcRxFVeTIcfea
AKq3PS6kJ032CJsjjB7NnQEwayP44qBlnPdAcRBAiei/ges7WvHC8lJ3fjC+BEHuv9fTz9U2hruI
WYAka7SMX460C0Ya+vw7WDiXfFD12GTNmDgs4KTtTNz8tMvuETBlBqzReBgPbnFcrLhe3LSf3g0z
8mgUs37w37FcWnNLckP5hjjgZHiVFu5uW5U/nTIqAJICtgaKBZIpWEW/P2WCZBhgK+NmLj+zCi0q
wwVs3GSW0Z/plT6pFbiD6wU7gRaFFDU2htcuP54VeFiRw4BDePX6dulY29xzLpViuGgGKZkX6bPl
1dD/gJQ9HkxBkvq3DTsrJCNX/OBUafCgaj0Ts7/ybdlClEITlUIEeL0ZM6AYkhlSgjt25cepyyZi
SwZJKL6oQvHcproBbbht9qxnp7OWsRpg+3ccg9A9ejB66BfnRBdp0ahPfxoIHWv6ejtm1NPYBAav
vRbUvhUTatwF2x6HHx3jOnwihfHg8CDv1oOJdvfTPflE50xO3Cov6HbzVgzrn2GqBa4frLhIX40n
yx0xd4Wyk1Asroe5LiHnoVjU8oP7Ax9NvLSqwWPizFHnjklcSGrj/3YPiqmkqtSVCBXLFTQwE9z3
RuV322mAFedw78ZdyJy5pzKx4GSYm9v5hyaphEKLPnuY1WjWDjTaiJuirWXeSHTWSZXY8AeOZWxQ
JtWc1/QcY5L7pNZ7sP0YG1M/zVqcZ25+gscTZcX9ZVyw4/4rTixx4k0nDgFL/YR0qZkLT8Licchv
Qo/GX6CMIOvNRXuMFWtPnuf6NXZ/mNUHTeB2k1tRSw4f2xhRF45CjFm7yJXjLsFqtWBdNCdyALz+
WJ3j3EbbiAhbY6NaxHAxhTntiwVuMDJLiRhrvm/sXhyUXXTRXZ4X9EYqwmBIHf71o3CQwWf5dAEW
NlClO3cddo1qwtiA3znvj/r7srUTpmb2E86t+63VIJEuybkHTHq0VaROM1ra4LIWL93RKn1pp1Fy
cUY9d7/AtCPxR6GMxKUqZ1dHiviHFeDLfaG+HJJfMX69MXmx1wUtQ8n11V/Vo2gbOqrfqC5doNmW
ew+JVdQTG60HJEbQCGy2rpQCrp4XyUf+lD+7zrymut+KWURgsjf108pExTfImHJR4CkvKvPCkLQA
oZyz0jUNJ+M0hFTvuOZLtgTauoZIu410XMHUyGNCV5u4nCJtnzK6OtfB+CIK5QX5r5jbomMW8Ds+
y38oXS2U5N9f0RlyiC6zj+oNNhlDvmLNN30/OUHoE2mq58k6fWF+XrgQi3jrYu7Wsg9CW+2+GGqw
ygwzsdw3BWEcOS3zxG3OrllfGP1u19p0NMFg5neuXO8ggFTctAtPiOsLxvGySJfArMlwVTCwRi3H
xwfTpexxbCIhxOBKZEpFPL3rDDye7DQ4kRfZpWGvkdVHl7OCN8V5vSKXUJHXFL252SAWbt5HqacV
yba4fXgNXdKIszx++iy5PA7ZzDvPOPY+cQzpWE2P/TndPnNs4SsORZT3c5DbP8OV9169vvHk5pm8
8QBgemEBAZtif+4lRJpCMaYgvSr7JnWO11kkcf27w0A9TZjFzQ/w0w1MZD6YmYulNEAr183BrqJT
mYT3lNS7uXtxX8+pHNSlbBISkA1IV06jWMipStT5JUKygO714i8BNZDn0rOjgVa9nLELFP2h94am
pqwPLyjUsltxiepdL4JigHl0hsa4fU8M3aKp70DWvduJnHKWh5fe40MIp8DIwgJ4C12zrJNg9tIh
aBQipOxPAphPhA910BkHIr5WJox8VcbljabGVmQ6DFUbxGGuYHq6p5DLf/q/kpxATViuoKM6d/e7
Be/PeSOcq7CLT5vAi7glMjFvDiUqm7wzQ8nkVfxtP5mojecNL7znk5zBEN8aa2du+1FxS1OouwvK
efQ+/6uXQMr3QaRui6PAeCUWCOgnSrVIKOEXo6mOIYxfli3JV3nZHQazBNexNOf/8vc7X5P4Nz5N
76lT8bPnlDvQbNIABkp4Ue+MnXvBIhgpjro96fq3exGWO0HcQ9ZDVOCEnvpQkgl9gZLelWtIYgDg
0ep0OfgT0enIxnm6tAwhXi2DjKZzrvwa2mUoj0Vzxu6uarSrQcPsItW53Fbw+Zby16S5rc2iZlgk
JGLrHlzsRbXKk90GyLXeaPwQmmWvhe9Hws0HFUOt+TYbTGdHKHJPee29xFaD7bWCqsYH75JAQ8eP
O5vgyffCS8+FiXm3NG5erNyj8SBRPuCwVY1nZpg0NZ8rMifh1Py6/8SlyMJBVoe3Ks+eyJGNosH2
6gT7IzwY4sQwNNPNQQai0Eh3C7SM4m/m+tybzXPq6LSkOXYHOZ+yfzELPwllx/Stu1QD20ar0LrI
JY2sUqQ6aN0Mm9+rcB9vJaykuenjO9RlBBYRg4v1VDCziYZDHp37i+emIyvgM5s/5Mstr+m/mj0E
lUpqA2Vr28ABgARwu/csPyaQSsD+Uryv28ovQJ8+OPO38ivD0ruMnazcmZkxS4YgHmnA1fBiGtR1
N0T1AkvOQW1z07S9rurBuHGi9jvEL/xGCF8zl7bjWAyamK/xzCxX7aatTdumqKiAUtPx1y3V6dBe
JfNOJ4YJhHvsdJ2IscyCf1LoMyBgQ6RPt32tNxwwShkK7VXpHRMPwUw0WKFtq2Hrn3uZ/NpovK9v
IaKSYZW3l4kkmB2p+TdjuLii/vvtf1jdrGqeh8HTMeNgy29v/tcw5yHVtXH04razzKzykRVWhrTw
8uRVIsU1Z8D4aGnQTOLQP9O2ZKYQr3bkvo4WQDIi87Le7hw5fNf30sf8Uk+pVhH52fw8b7U12wwU
lwdhi+6NUKpDXq7D7vyY0aWjVhfSoQt5Hl0wQXjqvVF8avo83bTgM1tXVohVcBezfbJS3M1hvyeb
Q55sKnkJkRPhk5COj+BHGSd/joGqnDog14bHLGxOLBPLFpQ4/F+k4G0a1GpbMeT2tT30vOh+k3IB
qZ1gphIXVCl4KSJ2Vyof3vbh1NA5sCNIT2t1Y40Y2VeZOfGK4G+CjdxyUuVWo9l100Izhho+yIhT
WeD+S4Ahb6OEywyfJ6S3H/jAm5JeU7JSL5/iuo5EoAi+RvWbAcSRk4Oocov+Ny8Vw7UQLqAexBky
tSZ16Oz11MEpoxY+aYtUcyfp0LeMvK7H+IXAKywljS+2r+rpo/zT6/1N0t94/fASxu387AJvAKc9
H/Dl6rlXlNCiDnXrVfnjEFy7TpPz0Pnunc3Yc7pa8VYscrt7QhMcsDPMpTbkD784uHVEZ39D3JAP
gN6s2NizZiCqOZ70qkBIMqautL1eHtxqxcn4+QbgP7+HU+tgNKtnQEjJ18f84XhKOoCuwXklbcGk
dCsxbDsPpIusyIw/pKP0w2XeAzrt7/3yrYVxojKtHEF6doU82K5EhOIYLW/evvqT7DTy20YgU44i
JLcb62xendNad3XqnBaJ1zXbn7hbVjsiGDMviHeqhkB36ICZ0CJ9m3YXnnggDZXdv0meh079vMAN
e6NxrJzmvKui55mEzlBL/4/QNXCuWsIOCftx8LoE0eVspEY+meyYDD2MuSTFGKcGWGP5wiVFIoVw
PuCyzgaFIeDfRe6O7BaS3hArTbPnP4d6HI+7iXv+VWbxHul+stCv7U4Cfn3wjkCft7JrSO5l75vU
PzZQzt33ckXT0mvLpYGt0D99+bzu/wHx8CtBe9DF7DDpbvOM89HMLFr7LLFRtRNJ6bhngLUdmeCv
lGJFhxzI86N/a5YiRSpwqpFXMZ5T/eX69AqHrgKD0GR+uyAOGpu9kF+y6/BacoYmt7eGaIxKa2A6
T8alBXejj9RHuv9RwBf0ix7G+x7J5W1It00pnTHW3VTK1hRbPFw/ekhDCZ8U6qwsXtK13sgmo63Y
sgba1t3BnHx0XSjpd0wyUC1+8UzWM9dMQGYbCUgovw2FNFvPEmmZVYGKUgCK+M05Qa4wfaqvAPeJ
+uGjT0LoR0MKCbd6okmcxVx2QrAqKBpaPSFICyqXIOdyk3qdGp9YoE1KtZYCd7aYwZqygtJYM+ya
YTLlOSBObaq7hH7unbTvGIMl9OarelhfKOpSuZQiqeECD8i4PsU9tFpj9m+UyO9u6OpSSerjlx5w
VLhg81ytf7pW3ijt/U0B5mRitE5k8dg1VQlZtTlf0TpCBj5c5uJXrmHdLDv5jHaW5fSaNwkpkFEc
cN5UeuYmG8h35l6p2KZpF+syjbk76+9vwy+h+RMxTUSAkKbi6f2acaFl7xFZpu46CKqZa5PyobGM
gvIG/A3T3cLZ15/thXyChYm+pzUBae5ty34GRAKQwSUuvSHDv1kM1rhqSvypCIWKo+HtDnsJuPdo
WfW+fnNjW9xclFD/DEZd9gFHjCXK2WZNe3JNWyC6UiYKdx3CczqVxY8x9knTAnGuUnx41WrootsC
ZyOc9SZh+XV9MpIlzVLR94cvNI3lv2ltC3dLcKS10ohVjFIl8vYDGu/6LaVTtv/jE5p3ptijeGad
G5SuTL+2EgHpGdL2uDWdFCM6UjfvfOOk+wokoIyN63eXS0l2nQ3J0RwZp32qYvTea62Agh4qZ9k9
oiV7WpvhTnQVTzqYx0YnAoJKG8LbaUzFMS9Bc+24Gc6Tre+n+zt5SLySDg5Me7UeKcD9RhUuEL/L
ETp2vpFACTJ2aWJpnpYtr82XjF5DZAAJ99vmWbu/QeXCMCGbpmyGzAUFlzHay1lPtc+iGrB1OZ5R
DdPjZ3pnaUiziMuOu+XfNPeZuXRdXnCdfWIgcVqWT/9llafQKZBKr99ZhMdGC0KLzPFefnPkJsKk
ai6GLW/MLX3UEoYoI7bL0cOLZW7s/+KcJqdNmbSTm6qZIgqaG7sgEar8XteGg6HjOaIBqJzSFMzF
E3yxHSzQ1HfxHwfRbBBlW8GjjOqu2e3an9ly/DVGSENl8ihCb9Z20K7LyidwTAwGPafBw2eBO1h+
ohCAdJxTJT8/hGPPZgORNAah03T9+Wjjez3zwXq2p/us1GXyxq4P/rZuwp1cKb/ECEE4090wQbzy
+1Q4S7qxkIRBKgYW46haoZT5KcQWStxAvsZVBRo9KwiW76TuMHX2zVp8Ph/YTlxvKFtqaMy7uCne
vTCVJAkfHx9MpOG13Mf1D/baYPaZb1AJ85mduIP7kNOnRezS8VKY3pdeGZeMoeUpNQob2viO7/Jx
wmVnbMLbcUJ6C4LCVHzJYXttuXzcP1Wq2v1k2ngP+fFp5OP4ushVZ50Sqo++LXwnDOyeEGfcBHNu
f8Lp/xWLkPzImyfE0Yxg6UC0yEIYqAxFkvELsLHdZjq897WZ9ReKnVwRrsP2ua7czVOGb4O/spez
4AygBMcXsxA1/EDfg19t6fxSYiXee84LUizkYMXjKf5CFqqCBZqbbFQrVfR/2Svdf3qcXICAbnT1
Ws+ZmA3kYed3Dz6Q5N1GXAHPBEmHEA1LZpQH9WlaebH+9NmHQmxMIROPfOGGgIvLfhYPT9Xli50I
GlpnXPO4z99JuRUh0GKcTTS8IC21wKwtXSlM5ja6aZGPrekCcHyh86xsqwQYy/RbQhiJ3gAqUj+5
ST6ZKv8oDbXxdsqAAYWcY11dMroS/gLkfCznWdyB8T2aX3Fgm7yX4oFgzpl+GH6tuXEk0IS2bTwi
2HvnwCm3RZfpf+ezmXZdiCjVJPAS4rdVhQUk7WH8kw0swEzOtkWG2e5tNygVc/akx9e1hz7KuOvh
c8zbbzrEDhqEMOwYwxR7eDDaIyEb+t5/zSVHRqkjvQywcDCq5hayTg5Q8LL7H1myXoQZoIUV8rw3
GvqEUZwPN73lypZgTXxxBY/9tGqj8l7dIKVLTsJ97WIwyinuhcVuzu1S2c2sCR4bDOlfH/qq2YTG
MmEB1p4oM7DAxR+3pbfoemDdyH+0iADCyCHSbYCd7H91XJuK5ekVOHHJrmSetCv8RDAA+6Zap+Mh
B9kw7W3RLYLnp/2uTlliMtGWFmKeKbvQM43imvrEMfgGvbd5D2g2XF5VAOKEhyESmaOnkVeBLvlg
ZleiWP86Y4Kf5S/3Ej2ZYT0mXaektJaKG7zFAwR6iafW03Hs6UEazYaUEmwe6uJpY/Xol/iVXt6D
zlbvO93RYf1fRIWONl4GZhMueNaKFPBWXp+LTPfeJdEDSsjV3FRdTzlPvouKiym7zgWOsYPc8wcZ
JKXvAkalxNkyPM+FKXvl+1oMiicxAjuOZFDQnMyc7VAAXyqNTO2pBXWaJ3IWlQH7dD9Ur62D/Wz+
+1ZpHaBzYjkc7iWhbXRSZgDpaHrDD4Z79u8UukZ2y9e1rNPDeu1pjSQv8FrgkdIAvL6crJSdoUyf
kUF2DL7eD0jAhpGWcykkfSxqHnJaOrOGww75MarhrrLE61kGJITIHlKmmsR5Pv2NndSgpoGy4ieN
pVWTRbgZ4b5Q8E4L7m6YszeA1OohZ9ZTQkAYAIgTLAQ+FqpTT9OyMu1Vt70xAxth4gW3QIMGAwOP
00s7a47dWmtpjR6KxVulLGommLFMab9Nw+B9Zuf06GIwHiXHd/hsBhnQer0bsNCuW8ceOeaLDp+q
H0QIY2vUkZf79IYH7H7BOwRGELDNGZkSMHdmKxR1HHpdGX3PQsnj+KWLfNpNvlays0sMAOqtcu2p
pA3hqYENPgfroTi/KaSgdzTdudQfBSBQuCcOyCFNGBBKw1GnCxxflrPElM6Yei4PdV3jzaWJ1FM2
B6yQ80YF91gGt9oIeuPf7A1wLqZVtQp0RM7s7USLdvB0hKcV9tjnTqOcuX6j7YkYQUc+o/bq9lrn
MjDSMj1HrzGA78UJpPezEMdDBjf0tl+fc+Enhvrg5cTcLJGOCYeWRi1a8PzO7lxvh2wk0baCud2c
3v3cWtyA//jMmH/OemSapUWT8DjpphXfd7wXkmaRD3ITnqAYZCdu5oVB7xOaGUapOCl+PGleyugK
Iv1yW9CUva0HiAQwgkYAhrkjKEoIqSoKnXHnrFUjE+J9+T2Xwm2NaHhLabHkldai7yPxwHMDaEU2
aOxtJavmoFiDUEriLaTB8rKsDb7P0Jj69YYj8TEPI8TuTx8m7EeSlIyBBofVvdBHuz8wL45QDg4z
rsCJhXdPPoTt10ZAC7lDobb0BEc6nFKanMpKGWIDR/yQd0l9M1Hzvm+kXcej8jDk9ypnLF30TX5o
uz4p1NkmxzQnG/AiCrtnrrrtoHgJgFl0Z6tJxkVa+fa1DLbrYvgXspJYVnB+2k7IY7LOXCm09VB0
QUGxnD3O/o7dUWvCaXWo7h4Wy+NkDRu/986MyU4OGAC7mOAjofIH/3RG5iOPdueoz2s2uBWJml5g
a9BqwJwBVF6aqIy9pc15NWq8c5P715dm0RnmD1bVTK2HujVKlyN3KbEQjDpPdyDh8D1bQd3z7UAy
Iv2NMjFD371VatjixKaKxhM7BpOKG7zO/PKHKJNUfFzwGnbOgs1noVR6adxyHOajp/5b0YBdGbSr
W1PYxmQGo9jgYjhM/FcVUdp8h2h7LKKmMDJPpH7WkoHn8o1ZhjOZP/sKie/VrNtVpcC1smv3jFJW
gvBNEFaRqNbiKrUzNZu95LRBE35+Kg3dtEbA6rJor7PGbqN26cBlPVWgEmUjBJAHQVEnjeVGriUV
dlTuc5IWn6rCzyXmpnO859wcU3SudVKOnO/ALNJRyebqvzaZ5+UGiFnL83u6aWLfb7OO+SNYBoyJ
RzQTa98HedS8XYXSmmZ6MvUXSXgVNPPYHUH9AFLOUZMhyeZTrEqybiFyZt8YUJjauOWG9gHYJA1X
LnkfN5UPudaJ3k01zeoktucm/6rm/8/0AuHq6P1qxcNavQP1uT24i1HGFEsTWHbpz/um8i7bJ6DZ
zY69ytC22OztsnOnLTsTTC7I6wQEnVHd05RpOKkesp82+QsFyEKG7K1AK6bDzhX0cMCi5tw7DCAv
U80RmRZ/SC+eX7DcWXSbGrgyZn70JMzW6QZpxcOboGNk41/0nMu9gCIRj9weP1cfx0vzbrfdjs3s
d02F09/HeS7MuBSMMvm6vczacH8E5IoTmEWO/0ZNDkfdhDCBufSubjEQmrQdX/fSj8pG+KOWqNXe
lEj4L+G3ATmPv/3i+urMUvig9AxaINhy3Nb/k5zBrHHp9cDEko8Ea6EQ3U2kRztEnxffxCeeojcJ
ttRNPyHgZweoGH20UpM2pEi3DS/6w5nGDIx+/SsrQ0zKUB3Uqzgugb4unq7tHUwpf0Xeelcpwcl/
XX1bmAEge9YwTzrJB/Isq5gTEoLyrbQg95KVULyMogGejt5MwatSNtSVqQgpAOy0Aoocq4Vp8vL/
BNvczOYMYWluo1WOcrOew7IeeCUgjmduYMq1qgKLTtEC+SBUp4a2E//cXbCbx1UnSF6+vYjK5toe
g45ThQUbRkHyDdXGcKSBafIW9NmPendFS1xOUf5sFbt+8nZW74+GIteUWouCCUcs/AzxzGJ572kF
gcjoJUPLUScHVR+tRLJaHWbX7fIG7Mtzu+RQAusw67s0qq4EylrT6+DnnGeKclZxLcOakHbOc5l6
+yrRaz0ZUU/9XT0ZKXVJR1MqTsutRwd1265RGpQ4Plq3pcmzXGJVKUaoUiBJXWqufZCD3CDnQuvB
wafdaTqiEC+Vj6InSUPJiwp/BSeLy5Ri2n9UY5A7+ZEG0dvdwFArof894UQl7eZg3qST7svwCAkm
HJ0Afoa/EQp/oKWJsuiXSkIjDAwEGvSIDDtqHmfoLrqEXP8yBuvEw9rKbgches8MWEY8h11Invx0
yGLIRyiPf5uHt18l2wSLzmRG1n3ydLnqMFW3JzdmZ8WdfKo9Jgn1luO2U14GfWXOdPQxfLHAZb5V
YWTU22sAXv3WxcQbJCaQaMxQoR8sjPtH1h06cTz010yxuQ/CtpcBD1K6L0gWzGWJvmuyi+cC6uiW
4cQliypiahDZsLC0xwR329y48Lhv+k6B+cjEBAOJrFX8bXwarQOaZmrJRPXg7i2LRd3gp5oh1UIN
BkxiGUhcmSfo3Fy+ewGLysotCKVKog4VUgotim7B9tBqpysdLK+Bklv0726QEFq/eau6a4y34QzO
DpM+lyTbHLc29Q8430oIeE7h0QdLyzw2TZxNQNNjiR4eFuIMUT3qLgFgNfETsUeatym+aPicWFOI
WqGf2MRIBa0ybB2ilmWNaprWdztpQvUEAHdWLFJ1fucvjrTybaMJixYtK4jd3dfQXR+fcVFuzt8q
lCdp5qNWOCOfXaFgXjI5yXzD45yneTylhCzMFpRae3IWD+xOGAN53d0frrUiEfvZ+qtdEyCZDAZY
ZOmek3UzpNNkW5pOAKDfR5a7AwdXOAzzCnaxX5AkXZE7aHEODusidG62RgzxwN4J0R7xKIHDnxiv
+cs9+gxXfajqzOuBixI9f4G5ovIoOSVoTXlLEfmJfre70Gf+spwK8f3NN6h2/kWFXScKhdAppler
svbDmAOfiL/g/rduFIy++pboSnyEGQvda0vW0H6y+qd88PHBQc8BVuKloe4p/jeu/1aQIQHHHWFN
z9juWoc06Q9qNip3p+xKJwZje2Jr+rhAzslW/zFDkywGvd2gTsmoPGOOiyn5f0VhBVnb2XwqOAtG
kvz86s0/GhnFXWDVpRSupjy4F4zm8CNGtvtntiJffBWZB3OIoWBp4jaXo10L2qS1fWkCEuzydb80
THK2XIG8Lc0dy/JcCPQ216El0CN2kEjep3P8+UVpt4chUxUV+nEj1lpCDP5Enaz8ASaHw2hICnWg
kaQHJbGwpod1VJshEz6tDkFggrYCUlKObNLws8XMsdSn/oAdWBvz0us9GU220nNbO/r3qlX149rR
lO0Wz2r1dcQ0YAGGP64KQ5H4aDCwzRdslKscZ8uF9odwq9RBcOQTKJYmmONS0lwE2rd78KI3e/66
vfv9QiEgkZLbF5ZAB/Z1Tv3ASwc9qproNsyRIEhqCEwbel/+SaDzr0JnVqafO1A9YUC8yEt1wof+
QzWDtItN46Gyuj/6VwkxIMHYVxmoxbDrk9XngHTRgWHm5ibQ6bYpVc5faGH9JNt0t4Lhkl72KBc9
0vykRXUEruwZwMovIs3q8r8WFN33hdolFBJCC+05Vt0xkJkoKhmllV3rxeluRmFDoCEn4rsZ7Jnn
vGhwyjx/L01x2lpeBVWVyo4Zb1Muxo/xvX6UWJPJDNWMGXKBvcoP+4fkmbqrgvHJZoCVPRtYn1eB
9qS2xkLIoIErRXw3wHk26le/tWBd+hXiptH9JSugMzx7G7zc/hkHddjYkjUIqN9m1dZWToqdVCDc
SAIuUyO2iKChFeEExYFqCD6y+wb2cmdq3NQBV/ZA1fL/WT24qpOLBR2O0sKlyxJ09eDK7WDziXh/
V3HU76SiLhN8zHY+uU4ZfUI/8wLAcU7mJQlu68hqrV3u0besx6J/Wi+vmV1iyIHQuChGfZMqSiCe
M7j/20w54d+Y2HqC/9Qltmt7XS68CZiNr/D1KxdL/wZ7m4TKENYDGxWvMv57Y1gxvdaku9vi8nh6
2r6UikoLs+XX4iod9241uavKRpU7qAsEGuBSytVi+YEzR2lI4IHg/k6wxA9oGm8E3otZhLAiHieH
dhZTkueFoIxKyrHDbVaPjysTAXNUb62HWJkIi4JhdbKwPcZ8mnZcodJA6ZD3igEsCwqHkdLXb+Q7
2XonELIjiXgwQTz/plcKHm7sBsZnD/401yoSbyEICoWNkRq/seTS2vyMwWN9hIaHOolKiL77THCU
YJtw1UQ8Sgw+UHviwVVQaUmM/f/Fi34yLRVtWGjnwJxcl2L147T42phZjHb4KC+O24U5dJhKo1iW
MqQ4oMkEi+FcN4hfumVd9mx7OR84xuPKpBwv0oEWvHtxBrbRGUn3oUL/Hw6aqimxCNJqqHb/dKAr
Grx5bhfVel4qx1EQRqx2Rm5iIAgJMeJve4wlZ3EzH45bJh1LCMtxG6dirp3iW/pX4B65xYQQ7r3R
0dGeNSoUWSVOkHMO8uepl4iZ8KkTHB5ZEfgVW5VE1cnh8TTCWuQjO0QoUgyd2MXVKv30LEMWnxQy
gba4TfzRHJgvBXBgUnzSoHRfSNqEVuvNXZi7xoJfQ3ueTeXsX62gNfP10K54/0NQtXU/JfxUHTg6
dnL142mpu+5dsF32rMeWfQnJEC+4bInO/Ufsa3O6XZCjS9Mo2ncNO9J11rOjzfQpC86fchsajLOJ
rOQ9r4kR9TBkE21ScTXS5vpyk0s39vLnR/D8+ffGGuw+6+fqtiFKC5BrmttqnftMDCO2IXQAJr9a
D7GDF5HqQdsbdqs61IMi9QQlIGLqqII2aNG1RG9Hy2PhKo498JeeWoRvCMb5cS35Cjt5elB2h/Nt
hiN0Wc99xdNz5eXQB8BM4XyqFsWlPTzvRmU5eQ2cm2CmTy8y5X8lkKoXZd7KxVld7b+MW73qlA5L
+aVOQioMz/ygsGPbS6mCJ4GHGcRibn3x9GQ5bN7wtvBbD9DB2fttULlQ12Y8V6PpPuQCgzKpenMC
LeB2oL7Y22PWXEIpdvlb7DWWA8KGGEfF9zwpU0eyl9CEmu8oUjFaOf3fAo9sL2FS/JHShDDOLDnI
lH0ri2axqBIvc8YPRXhVEujDG7xz9Gmdb7O7mwShMPaP8r+yqekohr+XUwRHIplEtJ7sdzViWBKk
ZpdTJMDaKa7GYHOMLslQcCOdXP8+lk1Y8Hc8TTS1ev8M2xpGfbzuyD0She+Vzdd6ktxGpBtGucMa
SeQJHyYFa1+6irc/HvHsRmRF5FOYxEtNgH9IuHcBlp3pbM0KrUCnPVfCMF9sXIU6lwyChmEkJxsh
2ybxagPO8ty2zH8BMCdllhf14PBbzxHUbDFUZKQf+5NuHyCdXiqJqtkKSG//2gHov/nfpyug6SR5
k53iyMq2WWTEFoFbzsW6eZznV9OGJKl5jQGrtaRuQWBSqlS4pd0zNg+tT0sc5VYrAjneExykz5yU
a0svpLbGl6U29AS7+JFZNeFLbaiIS3thK4LT1Fz363SdP9nc0hWir+c7PNzinrI9+A2KytYFxdFF
9BetwPB1jEcQpXEWo74e8eSR1+r15u9RvqI23q7KSE1l1dsj3Gofq8atlmGMCfij+Q6uQE2ONyds
P6d44sdHwVSEJZ/mCzZB89eMlRk+2o8j8dozR6Dvjmi3qUAc9ipMwrM5MCqw8wQuF6kwwM1V5UwV
9vYi7AW71AhqpFM40T6pZVdTPFLdY/rkV83v0Z2RvR+bEX+VjR48h5qljxasBkhgG7eUEvF0LElY
7iSstxpgrW9E/Mmp+O4xNF+aSqyAqt117/Uk2wNbtKZCO0VkCUmEs3iGQDHw4RhnE/1ZrazAXscJ
pLIoEcRZhWGutpy4PprIWhqsmB7U4fcrBwr7gwt2FUY9Vfov0JY6tfKs6BKxzPzIqyiDWAPt+dKr
WQW6VMJsTmt65xocABWUDo859O8nhPO9HmVxIZF/QO/KkE1w62n5teQL3h8CM0HvIxzufrvLtRPp
I1J5EqYp2f56V1bXxApS+WM4lbIfsPJW6/vuxzhZjKPeIcttca6/Bt4/vQK+Omkng68c8QM7u2CY
gAbiSDdlZ7ygAg5xkD+c0WMHt2MA52DsmgzTHG3fowb6VV3FGi6WJGJaQrK5eQpu7Tg7VuMyqITb
o1Ud6ivA4RxkV2a995sctQggumW985YvhgYC6+FmWxcBGniNhgn0eBG6PLzo8YSBieHtiLd3MWZV
8Zw775/awmrAWim59P2OV0Ai8B8/1fcgUAnGKPNApVsPwCnGFhBtaDLl9ReJ4mP5aN98UWSiOG1D
m872Jz4VZUT07vnr7XWzuKngGX93grHfjY/S1spUy8FYy+MKDtrJoY+WDooGjIZTTrlOks7kCRy2
Q3r5KFQiXR+rHQVzIi718QTgUOrkYpGqFOs5DdK063ZkiUXVIRr7fG43sEcCH7dYfuwhgqoOfUmr
ZInb1luipomLDSU2i4wgjLu0ws+4cky5YDaTzOb2xSYa97LjKdcNp690zdlPmW+A8w020fgpbP4w
X0HPG5xGfCmHeZymjT5pJJ/iLs9PZMQ8GooBI6+b3dHSPBOfwCQvR1KLTy/+lnP0qRyFhP/l3/ol
mp+1E1kJe9hdXG8rf23MFn+5e+e/4UvLSSK8r+MKEYkJ3TPb/OYP+6ocWj/ymhz8rba0I++LyCs+
miU7RooEuTxq+3q+d/uymAYWePkcwKxImYbG2QiTMk5ObzWhpwpRLHj9Fcxpb4cQvhn/2dW84lgO
alAmLyIcw5sfw6w3UScDDPiaL32GC/NibfA0ZS3fzrU8hf25GTzj3AwWCG3WJR9MtFkAeuPXVVWi
hfuqzc57MjvUghmDRS/RBMbfhDyjNYXsMNMqtae/MhacT6Nha9jACWx7xcBNf4R/qq4AYaCKY6LC
o6mIwdb25w3/RfOImjvwi1zVjvQ9ZGEwWx13oUZa95rDVCkz7Qsn7iDW3rhFjGW7nLEEeVVBxKN3
q3Za0DOcZZP6rE0FezQuZSf5wP0LCceP+F6sfzFePHnsUXgO9AaI3+IBWMlKht8FVbHi66tczesP
dDz5l0ZMZB4Wft5jozSYHSEZOUL04EvktXUTx6iLqbQaDIIZF6j0HCIcnPG0QoEcff3wqc2fpb+K
GzW03fEGLkBdCITr+MtydSy8WzH5Q4RJdeOEg6Zv74GIxAns+B+dnA+sLs7MHpKJ/OgbohfC48q4
qPSof1VgQDja66Ajpy7tZLPSP3zoPSxbzy0zG/oUrOM+EZZKvmKCG00eurHITaQ/h0IcVmoL4sS7
BdtmywlflDn7UvI/REhERgDPQ9W58L1E2IwGlbDVXC7kvpJCmKvpbVBowLaAUsx2GCr1xAt+5UKS
NUCeiNUa4NKNdoRDvHNLG5wqA+0z0Kqrn1SU3j9dWq0q+QTgrLTEEL3xF11VRth5A4QG8xJTnVIP
d+pTKHk9qSZ05vPxLvW/ypHw8DlxHoY2oFDEx2jjv8QlfHZ/WimB+QUUW/GV7qxG9T+OySvbQwca
GGI7ldbUync5NwRmhsFy1bUJrt7l5zLvPbLgrME9eHKcW7FDKQq7F115V7IfS3WoXasTI5eDpynb
dc3S3TV4M4MmBTvCcwUahZoVmUi16ShFJEKNZljvnlFvIoVzWoguvQ6y43z+/BtNQXKV3HwVI1hB
mTtqz8SsURinHGHwBEqaQd+YBuu7uA91Pk7Zf6hDrxoXh7nmRgZyADPgCQlgvKtIqTdOAfXVo82v
N6a4zOAJDWPjKICTWvzXl/cnF8c3swhHIctHQSQv3djRmskrDl3K2fTDSFpcJ6QkXX4qYpRwAiQj
/o0T1v7SH4MaJplwwqfBIYuH3wNuKwhhaosExUpNsxpIAva2lM0ybxIhui78UB2MkgfCfQcqkaWV
TfRzdGOZgfjFwSBitmaz8Hs79jx1ltbHV+axZhAigxq8WC5Kziio1Q/eZX2s9GcHG4VdX6bCp6U3
MdievrzVOosULtTsS5jUkCaHwudVUClEnR7PTkB6nP0k6tWXGanUEsH4CvLcMZ1wgYSuoiyTGUC/
EQ0UoSM28OU/ekcfH3kgKTMoVaJYFTHEawG1e1I+nZPnCzNJ1l8a22hOkx9FJ3ylUAw2ba/gqzCo
+A4NJfXEqsP/05l8XZSG1Z/FwxObhFuPOmRMj64EpmwuXlNFMlaImyWJNFGdQgBgdDIM6D1f+FGt
Rcebh8NOqqAtoxha83fl7XPT0gsBs+5jIXi2TBgYBRkaS5MgzBrI60ScY5DbBph+eULsEvClXJyP
dEzAFUaJaaXY4j6EhWegP/6KBZmWJZbjexMyS/fZ1NoZuyBBe3aUblU9yk10xqjjHcnBrUwVGreI
3VKVCVGDscdxerT/w/500SJZh9YG874wlz4LVNCR0oPSrj9GL8UhGkw5zBY8KXDlb+IRkeGrJt8U
vsRVBTrnKenHh3PnvEDEVuMo5/weXO2FqguaQ6KS2v5IS5mcX2DnJ1mYs9lAXHrGLXjF1h0MjNM1
EbDkPWsoVOTeg/zRvcyQNMo3bJ5v0mfIz1HDsxFzhBOEe0yg0r1Md5IurABTsXAmceMQOV+tcQKM
fvIbf92omSfMKOC91R3J08bXiH0FyfiorizfijFfEODyfspn+x2sXWTARaoss67aLZCslaT1lsPG
dXQKsD1M0jtlHCwcOt5jrJ671CpiwZEW+cye5O/TYOHw6uQfME900d1ZCKXIRF5Peo+oiDl0UjS2
T7/juqOlqomu+IJBXOT5l1vm/NAkUIdFmpzqbQxoAjg6JV0jBODtZQiWY4J9599Smgk0ya0U8YsR
RZ6iQ+fL7mwiwA1wKKqdeIch0ieqRKI7/jFKgf6MPSWAzOdXwaP8Dor/MCTBeudxfcN4bBFSAG8r
/1O2tFCjhSzih6NUvDAOSsnh91MsFSayrVrG0QvXPHemgoKm/d6r5UNiyg9VAsrKFfB/uxhs5fEY
S9cGuA+LwyKeHXBQKToorA+7YecNAD312s/lpL4Os0LmnYQVz35MgavpS2YJXKl7BRwMteZ9H2c1
PtdnccnBGV5AtaU9fPE5vOJPvYHf1aou/1QXa4p4xn3566Uf8o36JRQvjOl1ucfNsoG0K5S7NJKo
vSGbJwR+cOsJGjCdgSX3jP4gFwvF7aRpUwNGqP/Is/Fz3+AtdTKT1m31mDfFypRcWMQ9+CEPHd3l
PUnhYlIZWO/FBzn2n9vnonw7xBs5e2XQccyLbiWSUuEP5Tlr6KydxtvGhYGJguqXlcpqFv3W68CQ
biaRGhxME4ywkpgcapMNNR2vGeIDpwqbgf08sLloR5fWaKAHPm4h8RNe53JyI7Vj1fQN5sgklnjH
mhtg11xghUijyjix2eiwqt1BQDmUrbLKYZn9kpnsrfILiTofPzCs9U27nGR7NXsYIdj2CKHUkq13
XUtA5J9zueq6CYMvla+2aq9nt/Pc85Fmhesanqv2AcZ7Flu9fBGqnoIiHkUxlWZvqDHem/IGfWJU
MBFhBpn4YiRqSg+dAaJ+J3IDUO3FtkeWpo92r83hhgNfs7sOvjK7MMwMuIZkppDNqS4D8utiJ7Lb
+qs9ZRjbXPGCUI2HMZ+gBKVy6JFhOF2exCzumLVHQ/LMQa+9F2e9YVxCnSy3NpKVkssLPu3SVMR2
gYTSIq0mi66RNk7G8h35XEH+fW9OcAJZucn5u/t8EcswFcepX+An8Zy04Vn/gcStkYVRhFLHwk/8
hSmZ5FmoRdsCLPoairVwDs0SEwaxIET4nvdajlPResn8TwYWGRipJ92J0EvflnVNHJAEbSz1EnaN
itbUPEsAQc3PZ7Nzvz+oGnsRvC9NLLBD9tlXb3giALCOZBkLPRuZomY6YWES2XR1Fg5x50Uq/pMD
ChGW0fFEC3gA5Q/kjKddrC2XR3XJ4tbv7TsbNB6goxpo/+HZTKpOq+8bFDD2aJGM2mdI6FnQVGMw
DqxK0yCJMi88MjzSI2xrEdTyH5YUJ+ZbR4bzQwfHI7FbJUTZSZn2vHOPnESsiOwWZIWAYNRdn6r6
hGfhyGltz4TCkvpKdpVYJFpsyFe5Wu+X3EttcVwXgnrk9RUytCsJdxDga4srir+jY5gRLWfzlR9m
2oxffaCHE3G8cHd7Z5DyCRIkn4q9a6hKvgp14VxBq7m0HJw5taY4Y93Xe8YtFA3aJOvyjcRK7ojA
F41g49+1QbgqwHd5/EvBUN2F8dGYbbAugVQK40L3zXYFQRiEM+s2p3zQaoFbnGfVzDGVm+6YUTQf
xni7D28vQ0tPyB5FkuSbkjdRt1wgoIighPv/nY78KN+/52twp4vKFSd2MYvz5ELnkMRyUX4lO3ld
btUuF3BdHZkCxmfLUgmv+uaalHxRUoWMFUz6E+9ob+OmByUpQbwf8TmU317vqB2LM74acfZDtYwu
cm9mGCj+MR3LoU8I0ZiKRKeScbbuflCmY/AAmzTTYnaSnj76d6x/hp8qN1v6YfDBAWiu8s3FdGAG
QcktEeUs3aeDHKOIeM4aLRzezKi3Siz6KntqxZgcFqyZA4zBWI27lN97RBl4746mI1IokJo+Vd72
pQJMk4a/mDBQA6WeIrP3KbYBHKEBFwmFngQ3aW7dwbu3+iNnfizq0rchUKPumiXUerCvUhMoW2m7
VFd9qUoUmPyxoEVF1WbBwGXzs1bzELUQahvhcYj+OFRz2OQL+wYlK8TqYzoHOMAecTtQ9cnV4a1K
Mbiz0qY3I5UgS9gLOkKr4PeUZrK+zspVqinJa3nCgNmvGI1EqZ9vTSE+F2Uti3/bXoFuANFKCgpb
OWh8gMI7RCjW2gFpFKzU7E4kLBvEQH72KzFidB3PwZ6H9VwSfDSFcXSTo/WObg58ebznXkI4aLnj
wkPrUkvL1Ulf1Oo/TH4b6Ugtkco4NVH6/cLOVfsjbff9oUT6kjnbArGjxhsFeacm/Ca+jabQdxYX
r9ILKpOkU4OWHZKawcQFH9m5Hd87n+ecUQZ5M4kWh5ITRSTyAkjHnfeZa9AuNLQsoEP6KBGwUoBJ
9M8eUgb5iabODiC1g8u3SQ+5KNLWuUkzHWKWxzUOt69YTsl+Xp/QKazxGPf1POwTEgWCsBgmfIg6
XAHUqsbwLZ3YCbJ/fv+/uECKNS3uAS9kP0pfK1WyXw4CxpAmhsrPEn9NbrmrxJ4TFoKngrMUjy1v
Hw942KGpxH6mefHyLgl3+qclmVlI3M0RtEWy7JKe9UJzv96s9fHctdiqq41CY5Aza8RZ8KPl1/x1
qKoVAtrtIYbrdzcUIIda3DOWLQ1QWci2ADd0OUE1p/mteUpeBKV4b+iNKTs9fw5V8BU7rhmQzd3E
az7fgQvzBLdE13YyAMkbodk3HlixdA5itqw2JRAtZ8xkVrQBqURXMemSvDD77Ip22M+f5CpiwSx/
NSIRd+zDLyaaDgZTo3WX3+nlaxFcIXDkAwwIdJynZ9H8RKYJOq/BENb0z+dgrbdkDS3Eon9vnhyS
yeKH5wJVb8NtBegW+FjyDMNvl9X8mM5JgShXdOQzxG4Xhe1QLdixY5Cjg7yJqg3uSPALLrRhPs2X
czLIIHsZuhkVRjF+pPTSQLoHjQbq+JHKiRNp7I1wVhIGXyGd0Fm10mkCblIZnp3ubFjsnxHAuwQr
T7Cz6A2jttrICP5OptkvocUcvYIegNiqh0dhyzqr4+iG4EqpEVZIaBbhqmzIlepDcmDcmckt3OPP
y05WrvPOYCgKAf7uGBc6k+HdNRs0cnb01fWvc3WRtcFr+cky7MeZHri9BWriggdWtzvRcQ8iqszX
jpNCSeOYqfvoFaYRkWIDwxCgjKFD2XwwzMXMefetlb98IRVChkVul60mI+oVJa+R6zMnIRb6tNyH
WJ9UcLDbtJFoh9Xs8NSncG/jiEP0g3/06MSUAaJo66NFFupOTgn9yJ5f7Clb3Ihfg9qH3T9jq1HE
hUp7n55qTZDL7DoSf6HEU+++vscspG/xkCQm+UpoMaftJ9m4lHM6hccTGYNX0QsOcb/WTDVHNZsz
kJzg2RbSu2Lr1wLHcwEd6LMClzQYg2ZaLt4xoYp1Ye76Ecc8jaK35/c1U7cQQCkgGItXCmceGVm+
zDmsw0bTMBlb4vMTkunVujviI4gDabtW8vyRICRq9UpAMRHxx+gjahDBLo0VaJbVGp3LrEnJaQXV
U3F/C1UhyvLdvGlbx4DCEnWw+p7iIy78ODLOYYyGMNvhg7nXJmGfErrAUY/LfyoTLuEeDjGNNbLY
4sDJqThMKSkuOXWAtu8xpdIvAokBzwFRVvvJr/b15JO7wjc8Cbq2H7bM1iF7Vhgh5cWpMMF9KMN7
79R6isH2up+t5lxHSoKALa7ZfD3MFOrJhStJdnfnsVbEJlUwZYF0NDyBOx+hBa1/CLUjk9boz2rt
C8YkJHja47Wpmr/2K69YTTf2Nft+6UKJITdQlnoyKnvt9J+L2BdEZsgSbQhuUl69l4djZseP4unB
+8gKWsYixO+ekQLKtcT4e/v/xl2VJnqgNliXcqcCbuE1AHWOx4beSkCnpi9mWin/iEnx2hfB4vva
4n6WlmMbwGw7I8mxg/EfdXQ4QjDt73d3CLSYi4UtZPlj4Br2KSPpj50q91GCRRYczUlEIeZR5P+X
sG8MZVeE8VllksjZnbf768AKoIIy0FBxAPTdExQpWjaNuOBJcBaOSzUqvWhJhjXmyBHnVWQ0LcmT
x3fkeTBfBlM0E1Nbs3gUCOMsL12h+guBeitg6EKbx1Yc15XNBLRnO3oeMU7rpS4RTfPByQGmahO3
l+8z/zi7Pz7KlFbUeOxVwg4KaqT6b24SQ+ECI3bqJUA7Xo3sV3HFDF3Yri5cE72X6gRCbwZBfLWH
Byt6zGiqFb8k4v/T4d4xUXQXTuMudNJoiKuP3DuZLQJPzTGl0gKDDpFokZ6CkSgzdTjW1t8wSJfE
DJtFodWj6DKRotzgejb07nj0WNycqR7kKF30kQ5VGrr+rf0mTde2m+kWPdWFyxytJCaBXrg8iAF3
KNb5AyHg1qKug1VjUUsY1oCwH/HLViVQ61IzQtvFBUzK1G5qrv5OD0whyOe6iyxlpuz9TGgb9x96
K+TbSgnvXzo2otfIZ25QoqBXOYsS5MCrXrF2sMeL/n/7isJ3DYFbT7k6sJ3xF2md+6THPAfq0m6z
P14XWuxDK4g0sgZn9tZ+iAEwz21wM2eCCcjIwEnU0RSXRftlDu/p+X4s0RbhK4mjYFBdvHGW5amS
GCL6LhrmzgY9cZ41j/99W76DGRmspB+yF8AS4dfgqZwztjuQrMn15htVE0LXRe7QD8sRkNIUhzj9
SUV0fp29/OgEcVaXmPghAhnjLY0614nIwSxXbfaBilMx1bMk1RgvnP+3t62vbz7Gcu6CAbWxeB3Q
aiQup43GBES8UPFxoR7wedlLf9B+RBAuRic14eC6rmC1OGZeXLo7/+B1zFCpver6aQaKsWBD1YpL
eqWqpoTdM/Klo2e2q8GEii49EbLSO/scpnaFbv3dHioZQPYACy1/JMALWJSqB9cqxKyeLX7Yj9e0
zwhgPVqrWXkSrYlJcLQGNwnDXEh3938GDvuVE4At9qkb29+xA+AwB4wmYyfKtlvzQD/4RsEwoe8v
Yi4n365TZ6wywoi2F9uyVNtpG7adICgRNWTJyDZvhi7Bv421FwUCFwpd6s3VCUlPCUbJ0z0aoPIW
DU3vxek0gHDAr9JY0FwjiSWQFlGk6/B+GJfWF/cLLFh+n5CuW4Kt9+AulppcrCmlsoJs97v/9542
HlwVuVOrYVq9dMNDHStlswP/285K8739OY58mxNgYhgNBKP05zdtzfmrHGUM/f2+aIAY5PZDvOAq
TQzk3Mh22LKP/3oQtnzvuLQ7brB2wVMQ2XZzq6RFbIaigqGXvc2l95WM9zyWJqlZcCFpEBEB/ZlJ
fhVnE9hbj4WKOyJVOtg4HFwe05trAjlwu3nntq5jb3K1wqEIYPeQ6jL3fL0pcOqPmJyzvRk1SBOD
EvDXCg46DNtLjnlR6gfBmuTuHK7Isa3A0EhXKqs4wAUSpntTuPyaoM1503DebmAIrhRge0ZhwCL5
NenTfUauZekoy8316sBD386Rra9k05/lk2amuEtKpGSvwwzAQgjr5vlayMLiBavowKHHhtyucT9b
tPw8LlLnIm17387wpzh4d6LqlV1xipFhoXU3W14OXtaX8kCdz0AnVAjVTNpCe0Se7kFHiNLSkPv7
6bapRJx904c4DJdgTXlLfJ6iWXf4EG+4/pdQAJGHiVBihIkPqtpSwYA7dGCMy4MlmqTrSaxeBD/H
aTcptUtKJugbSxkJzpidzDhyJCHsvCB9Jd78ExTJloq0M2vbSsFuq0Y8/BGwQTn/5685itCWU/pX
bDSQA2kVcW734ioIieIK2hmMLuGUVTV4Wcmb0+y9bhgSXRJ/oqBwXfQerlfMqnycDMxLWlwOC/ug
TI8HmVnOT7Oa8soDxvqYx8t/zRQ9om9jDGAT58IQnpETxuNUJo8kMD6QgrWSVYAi9aRGBQFMr+tb
KuqtNozzEZdH/BQ/sPQbJo2bjNp04HClXYc3Q6v56KVNlqUbvkDi8QD0QpQyeMlRVbIXz8M+Qm3s
TshpUC+QT7yuEy9AteGkS7CgHrP5/bOJvpKmlmyalod8pTd4URYz3nkf0bPBmSdDxREER2ThrkuR
g+CPyaE9wU/mQRKd5ArDb3J0i0H0gxByE1s5BgvMh6cpyhY3JPY/qHEm2tazJi1FO4schYDMzT8h
3XFzfXFuIVFL4SNx/MLagkh+GuQVKtxt5ipcIHot9bE01OKOepliclQYLVVif8ojx3W3ZAxyahL8
qJ8EV/zVc1L50tnjLYPD2P2HPuSpnnum3zDznr28gZsnNNAgFdZu0Wsv+KAZFrbzHIi7H8YoaQsj
hGCKr6dMgw6DdjsilWrVxeRbY4bAvULsGvRHWLidnnjOLI4P28KDYm4XjpkiRBhGEnp+UiGIW0rT
jw7Gu8wzdm4a+Qd52FdQ2xMz8ajSyjpYNmcln4p8g5CjoeEkl3ylojxxgmE3anIjhycZcwijtsSA
oG2o1Z+ivFd1js5JP7NADDRie6WrafIvT3RcYbIbZ0DL3+7UqE9XaFjcqTwr5Bu97OnPVc6OR0k8
ipbf2Y3LDRyX0x+dk7JiGZih7xjXPor0MgPINpo3R+bNf9Ol9RCId6Y2kVdh8wfonjc/zaH1v8aw
OV1xkAlWLuoqahtsJoVRRlk5kO2v1jcHWG1fBk6+FsdtC3FliG3gUZQtbIRV+vri/HHgHLLXVT6/
PS1RBUGMaonLa3prHtZHu8iyIJfOwpU1Xw7sZu1mefLNIS9I1esUsHlIc6C19dYAA+FWKmdIDJ3Y
TFNRcOpy5GOBzol3PfsrCtlCBEZBXhqQ/9wINh6aRU+Z+WkJxOwSdPXSw0WuIcMc+/HwUMYD48Tg
3b2tZOHG8LL1zaO+KCAA30fUq/aUaOH62Ig/ut4/8XWb5Ym6GSj41LSnapWB2X1PEb/N9HxPENk6
fUsZWulNudVx5oXftYAcNiixPk1wKeNHgpwcjonrHY3tW7TdDE3m2PGruP38A0mIUa1g6/5wzaqF
6cU/4bppIkf/GesUh6Wpn+qD+yOefjE+nvnUccmRC0Khpu96CqUOZ2Mc5XFfjiM56lzKaPpLou+y
itj4AOt4AI4LeL5B9F6tnOa88Qe0gR/N3eXtOfVrlERX9uoW8KL6oy00+FsGf/aYLTZ0Y1x0ttvx
g9c9/NUwlaJ39rNUai5YvjLCXwPWBO3pW0cTGxSQtf7rrDF3Ts4Hj37udxqw/2fnwhK5eGQOnfHE
tKoLhjpfkNke8tGr5VuQrGiMCXcIJWJ/zO4b0n27nyxym7ts7/nrAaNCAk9bh8iDlpodTUFupzMY
pH1l9AMHHxkGcGN97Y9aO/INqEFkOezbXJPMH5HtCNRgmVPHaTFMV01bB7ikTRGhN1rWTPwg4BN8
j7QEh40FvbV5ZWHHD9VGA8CxXTLzBMwcoWmfWFdFNcTp3gqhtvscahNfqzXYy56cRYGpRRqfnd6Y
Az6GUNZ4+sZ6eIT1OTZBBcqMBHYTyG1io99P+msMPmW4bsFhNuUlHlFZosz023GgC+cDaEWRS5WF
Jv6wQWGGttpuj5eb2gZ2yFRF2bjoktnnlgR8TrBGpbwFlti0/UeY0hB/C+ElY7jsVy+fQAjB9wTL
1wv5eFOgVAjt4X60Zx1+jT7pB+4QkaGJ3qLYd3l4TniHv6IV2PoWvPptR/v16ztlmt66krtIF+Ya
0y6u8Pybc7WPyy3NUYFH4LGPSgpeaxw8wZLUUUFl3IU1jQsiqAdWzTP7mSePkQ7kPrrTsfyiRUWW
5FvDHN+g+IghfufVLI6E3eYLiI73AnErUSEC+eXyv93WlzbG4mhR+oW7Ptflhv1elyESSHBNx/UZ
P7lgBvirI8k3PD3cS6YJTNUZjeJopzpeYcrl17uW7AtIwlbSoYKUS0yKkrhcd7rR80H3YEAgklj9
mCoNtuyDaRCRBpZ9ghnwHCnuTu6lCvF/7YeWSxnGOYgfkjNPcziDj1EFW77HeuCUN2PLA2SioZKU
rW4E/t9s83a+SrtQdua38CJc3L+vdCgSh8ZLSoVjBfScu4nNjlQxtXKPYGKKM5ad7lXgKBlxZqQu
1/ehgiYFldYDHn92uQalP58KpiAb9jf0FzTbk62CKu4zFr4eCAexQcG7zgynmjfQSFzl7TtlPuZ9
a3rz6tV4KjGVYxkKAHIzySvD5sMriRJf+e1w4LNGMCNtJYvMpT6jT2OmOA/VueAn0MN+ClPYIps6
be3J+zLwLG21HXGbm+EIp3iBSLTmIOOMjrIkGNHXUBVwpDwzEbOo4QoJx3Q29OodJ86lvBjx1x8O
x2pSEH5iwEEJmwFoaebiUDXfNlTSHaghgLbxBCdCCb0bc2CR8MQN0kqNsBvr0SnGr7cesJRHWBZb
+PbdQGo2FQdI1u2Umx2UJnGBf45ujfyKgyF2pQ4tqyjFT1SyJzt9BzQ58smNe2xu36ZY5F4JZRLM
FylwUflrdblWelv0zgQ9n4yzxF1G58B7sOvf1jqDRueBG+VBQeGe433eZStWYQ7i8ZFsGBTtUrmG
eFdMyFUhN1C50/I3qsxoeGB89EWG6Y3Be2m7mN6Q82aCMdXTVP17P5XlbEN9RBpQlLDbnTlfT43R
DPMX6d4uoLT8c4dgzj1+fOdTBKVcOCWrtapb5cJKS/RLc0XwexOLlDotX6Wadu2VHsls/cmgFAgX
M2xE5+sFURpKih+J+ly7ptcsXJ7AJDIeoELks/Cne1G9uNpf2WXh2HafCt62kZyWNEZjzz8cxekW
uAcE4/TDaCIzK0caqanqtE57zxywNFvcVnzyVSL/AsK6VbcWz6yhaSs1vOUhIHwhNYfHNDR5g0Gt
evqN8inxaZDHnd7/JNao7IRoOb08dHboVCvlk0GR8p/mB8XHZ2PaZM9cD/6FwGwLRrd19fWDUbR1
PJrR1oHwHovTSdS1Zb0AdE8iJY1qxLxGYLJm7WIfS4p6fd8P/HD39LKkkYxWI549A8Pqkwo8WHxW
twlALjCztkda6kmNyFYEz+8SkcgBMDsCP93+25C0obBt2/mYyEZS6iKQxR+H3KQj7eidOfRcIBqg
3JhXHWv1LGQgWp6wb/EdA2d1vy5f43hJpC/OG16p6pV5iTbwe+MTQxRmvZyE0O+RnvN0mwca5Av8
t8qIWnnS6mBfwNmaLalZE+MKPSVxwu7agd8/yD1MfWsC7r3hO3mfd0G3X1SRa4Gi0s5J80CiDnPv
4imWWGMZ0iYildhTWFIOwSDjSjdozDqWDnexgEuPm5Oq3Owu8vQ+Z0iEvWzerIA/LGCs3ouQiE6r
+ZsppTYPM4B5vsEMZu/OZHcUaZN1XRDDQoRV6Do+fdw6zwNh/TbJazFCiZsoZxwhzLxQbA7acyrm
6da8ZTG1Z5UUoa7fFeaVsTPBXRZHhbMikcEDCJ6FMsXhv9r7OSzLq6kjpZEMDLDwk56mZ3Hu9cDV
62ZG8IaQ/YddiAaU65YCLFM0WD0psiDvGHOyBw8g04AqMno+tAYJGQyxRVv5EofIlsn+KwODK42H
7ze1s437F34QzjBBelVPnstneRP6NGUWCwOe7NjqlsM+eiAhEbrQVvDt6zhBqvfqBhhwkwVZsj2H
DNuYN/y3844vHtT+cxOExVjW4GlTX51W8JaVy3wsFquPmVg8UOCBU4XjI4AxybECyvqSYpOpVxmB
CVsTxCfzwboJCn905FEcVQJ4SMm+VoddWqdUyAmUp5wiSwh4w4adcMEwUofA/RyOmRntLNw3OwL6
dJwrCHNKBxSZrRw6rU76PsUMvTQYflPAleQUOs1gEucnNd6lQ9Li7zPOjRmaJ1bKSSM977Jp173A
B+WJmE5NEhbKRG2alozmE4L3oHLJL/Sm5CrllYIV5ucQEj6hiC6SGznqSf+MOejUABv1YGJYkREW
fV3Ye4yWc0fZ9xbkMGXaF+3I0eTLxcUBgsjiGUaHyG+dCpbvZNxMVlJ65qaFt1nfhjpDWxPUVzPS
GWGMinonq7kZFOWPqu5ZeaXse6hKOSc377iGRAQZ64yxrpIahey2RSrJwz9ff7YoFJf4slh2nFAj
rZPtanIotE132tNibocmM3NVlmc/BOoblw6fHFjs44oxE3+RZ1VmGCJaUtNpScm5r0z7z4y/KQYy
d5jq67KAG2lw2DbOmv9JFExgAOd2fWOQflUlRZgIYgWAMfZcf7JvauGdphfG4BUaHDYSqb1ZS9/0
pFYeYk2VUUKVje1EUQgsAvpnQSW0TkKo3zkEOpB5Z2ODHnk5rMbwNb0Y5Yog7ctfMEHX6mFdIFJg
6NPuceVuYZGP6EH6Y1BWSgxUWjoBcBUFo9GubBbNUrsJZ7wesYdsN3adnMjuXP8XENu3aFhAcz6g
NYh0tG7suyNYgWzQHVnlRmQkcML6vvL6uSbbbpW/quEDhjwdxHC4ot89LsRuM9EfRoVUbwHVlvBV
7GrExpFlCpc72poYC85i4qSZxD6B+i9Ud60JZmzQm1fJtLf6QpRvZqnotq4BQ2hzhu8gNitibsGN
TQmRsAkW9FFBvzO/KH/ZP6TlcW8x75/ik0/rAu76LSesfbUawL2o9QKwom7GJQjc7Wg+iFZrcV/i
fN89YGUzu9QzlT8BwMMPGujsOFumFgkW7o8hKgcTqpRKz/54CXJamtryA8VG3vfeHdLiPrcngy9p
M5QsVOuDScOEm6Y/zqA2Wix0BTREnzBeb+XPqKDJfv9PkxCmPDTl//pPD27oYC06OKhBvsaqnaDx
F5NCdyfsWzhdm6X3QYnjqLbO4HMmhP+WBcXbjq6rMAss4wOrykVVxIhAbbZSy1f8IWkQx1EibvOm
saElFgsRICZF1+PzFpfauHdQ7EwcC7q59efleq1mTpFS8hiY45PuCWu+jta++/b3afJKEY5M1q51
rQZOuhRiJ1u+6+e0FUwlvUyYnNu0aRSY34z3wT4r93shigmj8p0jH13HsrLykIBERuHYrevGCclS
rFpwh87JvBEpkYEaY73BMzgCQ6r13EkmAoq+euW5J7WNixLzDFuGv6IsYI74NUBO1gDnpLQRpuT3
bUwBRSec7JDgqvMz11prG9WFofJSsQA6MLNk6Ac1awisRlKcrNIVoz2Nqv94sm1hys7sugjjQrXD
6wXyOFtx8EFaztTk2rrlMMht03sHCKR22MkPIopeF5rMOws003vT0oLJMCE777BU1Gh9RMO29Rc7
2iA6lZ9HMYoEBIviURaegEfWkyfsgEqqhMQrF9+8K29CSIfNU5MEd0EKEIfVxFZtNvPjuzH2W1il
2BNxcsCiyXX3xsy6rT4yM8ZW3CArOehcThxHhaUOq/TMrFwjnZulHdGRbKQe8CtxdGYEHv3i2raZ
Y1lzH9jd0jheES6woimNTHcsZpjRmVge0+Uw8+6bybSGO6woML2EBYRGcVum7AZvV+y2WKSaDwHf
PK6gkebsVceg+U1bToHofsOqo0TPjPnIPEe1T83cgKZTynF+jgQ3PoSCpa66M8zoBolamYguIfb6
wpV/5INdNDoMRoOF79PNq8QOYbFdwYusc7sOxiiEDKZpg8DlJTaKudvUktplcoWezdgSpHl/YCwx
QFFoWHiBpgIwhSRCXzCWUjwI6Akv4ynlaj5jI61pVkGiCgV0mhH8GfletYj+MChxd7EQKRdMBioS
BHqua1OQxZTF50iCCgrSvEnRsyKssVpkIXDqyaoRUJjooJPtv5vswPsN40sxeTfTdluM16gULplP
6NQh0WLzmGCb7w/F7SVbZ98L0V2vxx+TK4mbJoZELG7Iq9oSMYstIdKuTN700n5EkOqpvmBn+WDg
4KkWzaPFLrESy+bfWJO1/LpKj3ZX9zWnYhmsXLIMJgJ1Zs1vVf4oMy7bjGFWGpzN51rhIDWdBTli
lzE4mh9phAlUIJmCF5B5ZO77wx2OOsmxiHRir0c43n92cJuQvDPW3G/jlmhi2bV1v6NDty7zeq/G
4Ai3jW14IIeS7f3WnXhcHV5C/5PMZSdK4ZMwe0T13BvXijKxplshxQOD5ZPRxUFEdvPhRRVobIFt
J2itZB1Ped99hD74LPae4Ttac066L+xMfx7aoroyNf8GnNqxn9cgfKtPEFaYTbJ9DmgF0Y6oevA/
c6I0pBJ9T+A3vnPq2/M9M+fNSmqfnOTw8qqfrhrL7Pe02nT3ycYXxe3Dj16uqWBEiWNA2dHNktWF
RiPwv1GqFWq5RrodqRW+DmgnG04GWHSD2xTAwqBV8heBEVO6ULkYKPMNxNw+bW4kq8LYF95kR69A
eDUnp0rUTCcdqyJjH6CWlncTHQ2O72sowqx0sAuN3+9P531BbkR1VTYGNOBKLItmWdRcRMeYBb1e
rj6mHgGpFXEGPtNSxbCi5pGQNwjQ3iAYrF6E7kikmQ2WpkyjLpp/Jp+MFM090eM/XUJGHdVveLqG
1vTAPW+yZkYQD1U1osDMRCppVgyy7b3T1N2b1o4YVrxA5KybSg5ejOGPtdrXWtDS+EprAIZsKkDK
Ux1cuTtxJS4b7zcOkrPxSOgC4TEbefIlCoo9dV3gOewDKOpRgWxR6NREiD+JP13kYCz2AoCr+cod
cYX5XL3Lon90IggwMIOUbCGv5p53FPFcRm3raxn8ZMm5hu0EHHBtdsbc4BaSi4NodjStmU/oZGGY
7SfQB3MqL8TmqD1ybVUcGl82VA8jdV8IqiOkURsoun/9DqkMmztgkeFCi0Rk2qTm7z/8J25S5X2e
UhIFXGp05xQqYzBQa3c0EUViBInjTi2z7dd7INJSZ6M60FbTloYXk+EWS/ayRuDasGRz2KntrSQn
YgQwTlf7XNDme/nZ1SSnSn4qXLGBX5kNxuUE3hfGZRXBOxp4rRoUWK61vrES5u9QV4VdoY3YHF3J
7t5D4kjFAy+WSssiQYEWPnB2utCFm/klp2lPHVK/H0Ci9v9yL3MAUEwU1edylpPB+JRcHu2kSJxK
nVuKFEGtYEHqFUdYtsskdBKMGf/9nCaOshJUag7k4VzKG8IZQH+uFoYSjyp3BERvXJakEMYI2dfJ
kRbsmsw/STXTRPcvfBQS26agIZtDYU0xNcAfvRHaaYedTnSVOjMa75ZzivBwQ0gfki6DWbCAPjyK
FrpPQEdGSljlzy3ezQ1RXeamd6Rrfr73em5O/4N5ZxKnmTReQPaubQJsJahrOSWPb9+Fc7CBRXA2
swvEyszsf/Zse8yeEhjDM83YJsOvkfVXg02Jpo4iL3VxwirYGy+Y6TWXN1uSfTd8Zilv+YVAonKw
zFta7mZ1yveXnL4qugd6m1k0fJ1mkBXfHe4foJjlLu1PkVFA77fy30+3jLmArtyYvdpZ4pDbPAaa
l4bBs4C1HC0hnHUAQrjjPqr/0eh/UjMt/09fT1WlZAK/iBpi/fnkQAZHFMMaxrW9clr11SLL8edR
95FrFcDq/AWmMJIMUhA1ZHw+FT2jhm8udlA3wEucbSUh6pLBOxPyzoc9nY1zHZplKPotg5cmpjfc
ReIB9r5Bph2CpG6fsZ9csuxLrNJXRZYDPloHypm1iwGalrHl3nl9ap5nh9K4TNY1XKCJhTU6S2/s
DUtY997vMd4bwyNqb9iqTnQ8BHvv0fYuiwqouEJy/Lqh39BCHGycs5PuTbWGGLWxczbypcJzA5p3
+ktaJ+EwZn1Mh6bUgQXU3M+DecXYVrbiHWWoCp59hv7w4ZYcFTHVNk3lHWtUGmVHKdYVePGyXb8Y
YsV/DjvCzqdiqPj34yRYVT5UQryqB2AF9z4ijDeJJZGa5kDSHaVaHLkE3fF3btlL4AoouYaqpCxw
Q27PgWOgJr/52CcLXxreeMKgAZAFXj8NvotKdk+6pIPgmwUA3eoFO6zyO695pfX4ZskBn1ncQEum
BB3mvPkl1kJzcMNNCITubosUMjjppovkSxNLVQTvtJppoU6WqjIx0CihiunJlEMSzamJRxOHZxtk
QW2X2av6vHtGCv3HvrDSeOpzvbzHnVb2SquI0H9VWWHfr2g96T9jFk6f1LUnPqd9VKlOFW27JTfj
vHnAMGlAv80WMch6ShwagabgGNqjFFHifoTA/CF8oR+dOtT7Z3Ifxqnd/2lyH9qllFPQL0+jCcEq
0WiXayPTFn3YV0/wnDwJQ/bQij+k9E1r8TDtWzb/c+r6q+VTn1zeah96p1bra7RqATqrUgqs98ba
d0nc04kiKGOD81WGMByXeZWvm5eckZEbFFk/U9kny/tcGgDAvxs326aDTMr5SwvkNEDjLrI3iVxP
A3XtlSXoiuAwLK7otIhF9elYZkl3dkCYz4eWshhXnnzabPkZiCHmTqP5LuzJIbL5GNsHWNxe7rCZ
RTk8hSOrgCqoAHbFX06QlWT2iJwArrVCsg5PWUlOCKWUK4EcWF+ekZN8kF//MR0gmkQfusfDhP30
NO5+EcN5z2z2IwuDxhdbsOS4hDSrqbHG0tCviQ22UHq0DSVvHLUzUQybTTQN9PDA/863BrMbw21F
NWPclJIcwdFNr5VScJNZfW7DIdT4j+1c8P+ZQOSWYOVxonuCpVzpwyUQw10V5Jo2602JErxb/S2b
yjhitDfqUa4RXXbE9aEZ2tYAI45z8Q5gIz+zJQs0maCOx+A+vbEvTSxvgCCS7IwmJxdLg5NvMJSf
ANPA/VsEtSqrpOvrYHqY20ogiPei7WjapO2DADpgAuOvTXn9pG0p+y/WBdFgKV5hinGpkH6OZjpc
cQt3hUZIKD3tPHVVDTbH4bklqhFeaTvCUly6kI5wU4MSbjdZ9D15ymAOPFdBDoT73TRcjarTGnEW
AHTbKEe1sEex9y1jXEenKihNl2759duALsfhyyTyMkaxpgBnoZkSVg9ztJBl6ega0bRVN9cWIoqK
TipJYQv37D+aN/AoYHwSLSkUyN3hrZ3AxsXRfDA/6UlytC3rqUXYJu3Afhkm1EsCeNHDJA8PmLAs
dRlpebzKqNztpvqTBfezd1XItXI8d+UdbCdibeU/V8LZ+xLy48a+CHYKTX0HsIzxqSAaRze3Klek
f2Zmu1/YIgN6XaIfNPrrx4g7HbtDUNDKM8t+0exnU3rT827JnDF5i7nHVtgYzAU7+5kC27RaNCBz
+YM+bjm39mcmgJcgH0xHkQhG50D3HuQOn44XcHXPEoWEP05596thIoHR/uK9X7YTLTGUcRDCh0kS
ImVyTOkyfO5MaotMX2CVXrAcfZLi6Qbn5WfKz1lGPfZc+TAlgFNJSSIdHJRpWGhJ7RfsTAgTdbL2
eOYQ2ZquPDMG+IUPDgbLfjL3VfR2eI6QqckSkdZWhJuwyytFBDM9LkrU6g1AGGMjPnmIYHdNfHLR
wUOyMfQw0MuNziAG5j5+65vBqRGp96a9pTbi2dO3zSATuxWK/gtvsIo7paA7PdvOjLutSA94lxzF
HVM6D/1z1a776vMkUq+Fmskm6DwSmZID2+bd/t58zly0w0VDos8TwAfJ0ZYzJ6v4SROuoi/OoV7q
R9Yd0Dl7OnYNbQ1wLXKXzJiREiRpOTnTWv8KL7M24XIa2Ni27zL/ZG4bx6Pg0g1tv+uRCkQy+qJs
ASblhZ6iNL+ZD6xOFCrPXX/AIAWUbgUtO6VTRwDYGjbNhqiA3wujkFG8AJw3VgRmLciozRVg6zaA
UiOyQV80TyMlFovlxBMV0o5ID8lvdV2BhdCsiMZY3sTV0nRJwxSeacivtHNE79KETJarig6dcF3m
vDWwNiSTC4WjfQ1NIVvImy1RTTX5+FmJGMwQ0OxTvvPiwfodLiDOSiOOFJ/XKAY8pWy5Q0oppJ6A
tZUEhdilgDi/1/8kPJYJpGdmrnGXiSTYd2NdoMeCVHcpWEbNOxdWXqZxuyDKs+UTUn4W2UMU/+OU
9rY8CJ4WP7Lu9Tj2XGNf5Vjy97su/Fg8f6kw2cpJQiBN9shaVELMrOGoMwCINpK7CavRl7a7N0O3
IvmNFJnxnBF2H4BpSwMFxsQmHKc3uQPRKAqU8HPCLZ/XnLRUAZ5MFr/LuV43J23WM7A7gKLp0O8P
zrDyIaBQijeiTdYho2qFmpguOYa0XAfjbfwblvGnnZX9yogx2YJsg6oYH1o2y42aGHPCK/rG3NaQ
K1aofSxW8FNqfRwxecFygj/WUVgS8bCwBY5Y0OnlSt3iMF8lGTsgrGVw7t7qeI4DT8UvlQoliWTo
s3A2NwwQowQJEVwjB/QPXNNsjwiiZecJvsvXthjynFmABWMdwuBI5tf9A/27rAL/f1YrvldKdAkh
KdihIIa4RFgl3zhaznhGcCqcydz5nvCP2nMAdU7QUsXTX1+NS0dtNwyEGda7nZSfKn4dB1llWxB3
cuoVdiOB6Rm5BaCKz7l/cxdppJEMdJfBD+hxcOwLItbXWUsWyULDl52Epz2FKFm7keCZ+LLZerSX
35PicoCQ/4rrknwpV1h2WA0b1BIAAJaOPLhkxn8VG9Nz7pJRGuCEmZpeNyyPq3VCDMqgGr2vo2cg
2D9PJET/RDwLKpj22oa8Erv5ILRuBZqGMx4SeVdU3WV79JcCPrpY+HyNm6rFCqh7MLR4Ps47JFeX
Og6pH54CP+ydvyVe9tKQ9Gn8owx/Vt5ALjAxFV7W8jq5qtjMLfTgpWFGw3tGD2h22eKl8kM2rsFj
DYKt7cV8qszcTkSgU3mY2tOjk/irMHWcRWd6NyulVbBSkF+RHnVGEBNUm36z/E1xPd46ajiI3lSs
e08Qdc8O3gpCG3pC7/wBxpZWPvlGuwxGIn8dAxhNluPVu8UN6cqGBWD0m1aGH1ZH1HXjBEyi7C4e
aHmJ/TO559GaRBq6tLWVHd6AhCvIzLRECx1eS1CeTB5/ind2g162qi+2wpbeIjM9/oSjUQbuprx9
6i1QjBSDapx82LQ5Kxr60GAIl7HwkFb8PQB9Ou4mazU8Gr/O2zm+0vSWe5SYyGi8q1UNlfd16pRM
ux64AqDEV2XQ+uNYvf/xdDM0VVJcjgCbYQiyExGhlfzk/BI77KsUQodyz/02awMPdBSplfz0Hr87
IeMGZEHDhqpF+e0eQ3yP6MSwiY2W4hop7AUUAhAPK3DC4uin5eKpu1w6oFXeSRoPyzsmAjYv57kP
Y4g6TyP5Gr9d3CGzhXWdr6Z23RWuRfGWr3I4DCv3XOyZoMLAvqdpjtzBL1PeDNXYK587uSE0A1+I
mhm3jU52+I/uriSJQ8dINT0FvecHpqjmVkiKIT7htK1NGQ4qh4nY7EfrCiQrHaZl1Oo0peFvV61u
8IxLWudYHtQS/TN4CCQOBXzAJWqpccY5V5mtENCKkO70QDHWeiydbdsODO/xgAuIhLa5nREKGH+Z
aLfOpRdwtVI0mBcX5ENuHqfxpRzg+YpsmW0Xk3y0FWIlUXWUaAWS7/voJ+2KTMzncnAmey5LDh+G
72cCF6OIgiQA4yck38oXJxswTuwXgxtW/E86cUTFEi2Tfw1NPUAsoDVNmWyUeq3H1oPjScWL9f2h
UtFbNML8K9Le4r2T/bbHvyC49rAjV7woHnj7YvWULJpJsw/lyspbutJKjrh2cbSdAt+kitTuHSSc
JE1kIX9wS7ibMRikJmm8pFuGWSdi4dozkXBYNrb0TI2RkOjaSpWocG00yNnN+LAkExci/yzAbIhw
z0pgXX4l4ePJTVD9eu5m4l0zuZ8rGCwr0R2MT2JK/bjCrdu10dHbI45b+W22CAm1ruKPW6FMVxej
S9VvXlR2EamWKHrDEh6oem+auLirf4UOC1NMhxOsbJLoKcd73T/DSI/BS31T8I3/5a8kG4B1yv9j
/tlFlFKrhThVt4f1Yxc132DkV9XPKDd2B+InTUs4x0QgnLwLczc5xNfFVcM6XFGA1tyYDi3Nb5wg
wzWLIfjIAGfJHpcLEP6eita3b2J+Ny4ALwvej+WkAil2KuvKkvKdaKjxk6HTXRA4bTSoGszlssxF
1Ap34qv41BdTZ5Ys/TvGGhN3eXmL0fiarhqJFNGbwzg8J03nhhzJUQ2Dc6JXuu+4BOz6PfMZRG5z
Pd3Zf/W84Dq+uiJYbZmrw59GPThhYmvTFJsY/wcJUoSqckm2A6Zo2YslQfvCJu8dZJ5DFP2dUP+1
sPcQWD1hKbKN59hsSnvHpSrP6ZUFmPhCGIUGuEoTjksiYwiOM8P1GK9SEpPG3AVjH9sgdOhqmPD4
IBXJ4CG6ONKn4WQJwJs/UDAPwWxfxOI/lbjAqwdbOyASRNwYqvsNKM4rPPxct3YONwDLH7udoXn7
vHmnM1mkVjt0nkeAZ8Hdj+OuBQtTMe8E7jH01Qcx9iX4G3CGT7Yt4tKYmR3Ig3DaOd4Rjbm66qAB
jTpJrcNNfh/ZXKBpH1gPoT3kJg8W0n7FkP/L53uwiA3twaBiCdiwsFEKrkVyRP2AZImkvSsRAgKt
hog0hzC/gAoQENaZJ4zywyGNVpitZH/pUN2hsdCcOKWVGQkeCz249hFSZ6npp9GdnQrc+qIULVvd
ft1DSW5LO9I7RC5K6UetQtXJQkBZM3mVEWV3TryUWAbFkR9NZlBrQTY1ZzrZ18i1O8Ceml6oAARu
pwVeL+xGrr46J5rQ9AbB9mFXdQge69yX4VX3E9EyF0cJzqS5mbahT1WO4yDPx/Ew9xb2cSaWFFHT
A65ejBSHE7qwJEaJkp+PmsqXebs0F8Yo0DYZNk/TaBl/QRtNVJS0Nn4RNcCoVzsDyo3mQI3VW3B5
bcURibf+i7az+tfaAE61CWjnFEUuleRbgaPniFCrmEs7YiR6YUS53oGn4pEL1YHnmQnXsw+gY/8E
0bbCC8WH4nOt+SvyYfsVdyRfU90ou2nftxCbdnTpYSAsIvpITALs0Ykpy8I/zlKU62d1wPY4iIVA
gzXiiiMgHNL0HbyHx/TCsTfjuMBKcf1pwaDahb0vuNEeJ+1JfCcIJ/0poCH7hS1nwI3v+H16hzY6
ow3xMczNP+chnTZ9o3ysDf+dw8UzxHZG0a3bMHWdY5FcV5ah+1F05Jev73r3ANy8XLexDuSjAeEt
PK5EaJYmc7YyYeP4K308RDtHFtwW1MqS6WQjCVL9daj79Hzv6ePA0VrZK/qQ9RjwMDnssWqv6gJk
hH5mcDEOvTh/KRTIRMioV0RSxxs96Xj8kaLlDCjwZ7vFQJxjt2vh2ry+75caBU1wtQ3lf5fUNh7+
q08/MXm3MwGkBFfqQ2OLkwlA/KhAwT02tRx8nU3QKdlMqmUgdDltFhzrpRn4w4jKapwOhL1EsWCr
vvhmrMJacTr2LFpbBewBFRj8ITzY2vqyUv+Oe1qJIuBAZHuZ0KimHwy6bqIYZBiernChhbC+kSIn
qPdoe4jkuz5rRlJQMiR5qu2r9lqWmlx9V7aHG+yuzUJQrzA1r3HZuRIhHsphKnQbAgXeHhGyF0ZD
lsyJdLHq0JA32e1pzONj8rfdQylq7eNzaWSImFVEC2q+K7ZhHs8Rbtm9QvgwbxACNTCJEcJpOyqj
rVCvGDJHgYfhVKqMeANOLQqEdWguIWNxDF5AR3qYDFY7U4oLoBILfpSlp7KQxlZVAQMOWXUUJ+fO
ERUwxdOsv6iwaWHwatUXy03mxywnZEfcZ2AXaf4HdMDeiDRhirqnLfnB37WgEVRgatqmwsWDTjFF
8XGAwBlRqWLnLMSOrzJr4NbmSxaQT5sn3ytqri8I6UDg4qKrxuPkMPQFEpOBCl5YK/zd0sr+n9OD
lSUtvK/cDRC6sqPVwRz936pEjipN65cxz8EFOtlFKAlTYBoUGs2XJ39DV+tdHAoB7HpShMRU2RRB
e97ClmwYOIMMoJKmZmdMMg1idnETYRwY2OJh0HcT9el8IN62StU4G8Bm2EHEl8EDDJBYuEDemAxM
U6xl/O4qW1hHN1B/IHpfgcbszxDi2qHxGX0dVNXG0caTRog3DULoQRFhnS5APNwNzDL37YMG9EFD
v5mDMRkHtdMSc548o1fzIdCrdDpR4N/imixd9gc+gEJRQ8TaTDRWJdHw4kHPee/MKA/N9stg2/jU
4seU8gRjRWDNbG8GQ82rtDDtdO6Juw74u588zzK14P3qQM1J/QHIOXxFTFsCe1XW10cT7wNJVnfw
QITKQSmfp2GxrZCjgzs8kZPz5RyAJtVBdefaLiU+z1Z+/L5csKRVNcdWRDj0UJNVj50WFgmOwxC5
BMFJWr6ecHgP7tkmh1D+q4XJGsseyfT54w2IwzSVekKI+z3+vuH3yhozKC5cDy/cQi1F+SxNi8s2
29DVJXbXh1F1R2dNiSduKO9UgxwcLONxmY7K5ZcGPSSO/MlPiL2BAOIbesXUluvNSIs0fkIH2E6n
obaWEPAiS+utK2avigwHiG0HF7hrKSkbMvvW1VboIPrplr9UjDkhr8bzBGtgOi+SIgPJgQHeQxFd
AjW7x+hCBw7z1QogljWe72wWfOh51a6gKbDbxmuJ2pAnX6kjS6Y0rUrtzHEn+Hg2WZt6dXLglbzy
t3ELMPfMsb8XYYhVXS+ko2SZRAH4EHj7/wA5mucM6+2Oycjxqd5rU/PT43hlXZDHKijzfZb3PkbH
1nsWyQ72wHIsorBC1wuP2F+sZXh90EjbVB30AzpCWeRwwYK+xMduEU5IF68DVVLYKQ2B8askpb9e
GC8qRupCTa4LNVEzJk9z+CqFiR/Vq98CjjYKJhbO5lIlIi6Vh7nnAxvva/q1VCxAOGQ6iYJsBw4E
q6pYruk4O5DKVEgbzPlIqxTD6FdojJpJeFuKhf1oKEjTOlZ6LwqKe2e+AWrP3eJwGsWhxkJwN33z
TRLEI54yHSmeJx4IVvYo1ZFaguux930aKp7+r2m97KLCSIS9ZYbgbT3CILdsEKWTYUxrtRrjK2au
iQ1BGyf+p/Zhtk2jBfSSu0aJ/ZMxSEYs2ThjglIr1keVbtFPv0gDC0ABq9X0iyPI33ekwjl4qwr5
YVZDiYSFzfIpnIp7yCXwNwat74r++SldUfWleS6l/pVuZyjG8fJ7rH9QPsqwC5FbPo4QjyV4zgTW
v0X19ZdWXNOp0UVFTGKSAINyw9vQvNU51euoTVMPj81MW/tn6dA6va04HPT7VI8mwAsO1kOD5qBO
cG/5xYt5InmNOx7ODeJ6NBTQrz8G+UW56xOOh9o6F5swwi3jdVSWFkqS4pfkGl6a0ddpCb2dUPLq
vUMJXT/ShDZUY0d2ZKP31Tx5lARslhgZT6iWPVJxfZkivDLeRBEcsQCIkCgBaL4e42QchyFl8bVb
xwyGcU8QlWi0FfxxwlSPsuhH+YiXvx2XhmaoLxc83L2GeGwFwDWZo8u4cJ8ogAzIxSaypgJH9vvT
aSRH5EptyWxjNm50bFRLwYiwI5omx/40EJf2Yml11Bv42RXrXifEwdipHleNesI0c8fo86i+P9cn
5T2BtI8Uye2OR+SVPIOUDPGzkRq/ZkWAHVrpkybeKDwEOSiV+34sP7eE8nlCspxnyfW146vjxsrY
ON2DzShF2tCYE+nbnE/s6PD7SVPhVV9XuMUIRv7FdZOVoqrOczPzviM3CR00iRyiBQVNaAC9qVF3
8W/gYrTPyGEDpUPcy6TlI08I1eE+fF8glIo9cWH1Pjb263IEU1WtFnqtxeob23hpPRPUpGnud39m
BnsusasWp62YfkEaHdJ5Mc8dUypuKzWw6PtMe5oM47gYLofznZuFm3kr0L3fRM/Tdv9w0orCtUxA
3kXGO631TbM9xBsaeqIyuFJTFbyCGjS2FkGxUkpZpOgoqBb2JYKtAySU8szolZb1M2UscOVWFTmW
IHSVLa2sRpRCXEWk2/QyQ7Rg7xZMKAIX7MkVCms7sujzf6Xre9yyiT+13wAHCLXE8Xfj/p6LWhhE
eXdp2FXUerYlHAM6NvTELhu4goAfXolSCsEdwIEbZ/R+WiGJ7Xb17Om4KmIoCrpwxgh7u2JRlcwu
4yZDO9lmKn2I2jC+YBWLu8IekQNIQkffCx1lwXwTx9UWjB/S3Us8JfhXyDfnxnp8KbvJ3W5syzk3
Eg4XTNExibxcPXlT6lD/djih//xlHmO+m+nncNdQfFNbK6CKxcU7XEzBApYQBsGwq/J76dNn0STp
UWcJgl3oMsmiYU31mc5D0CYcLprOtnBs7Q8QMsUoWxVvVyLCL1z+bG4A5YFB+E6Ga789bIhHCyMG
RS6dyQEvqbREMdYxJypqF7TSplfFwROy33u7BOVRtdGp40QS1sYhNBT4bLlc85xSTviXFeO0zLIM
cLIu7WPuU2rS2YLPdPbnKt1k3JOJmmqYK+KEeBMXIvNwMUUyhhlJ/zBw5m+xtW3F2+5w7DjBaQ0h
rU/34b9FfL9ksewOV7ZjyoFkUc7QNAtPxAfpYZidztrEhmUvXQv/PyV4eXE8bBGJokKU1PH32s5G
QGizEELMOjxNmnIPmTrdm6z8A/q/Bpfj8jF3+J7IwUkVWzAYyLddbN9t2yRRCeccPcCqd5FEzUVE
UZAqKCmLmxz7T16RrsSTuYsoSKO098KydoG7jvh2q7pVzZ3jkFpVdBWTbyKuMNiubFFGfwnI/ODC
xZEx+SdxBp6bo9qFMo80MhGlLeUgydoMQYZthFTzTH7aK2BiS3aCH5qbbVmaG2Z+djal/FfOZTKZ
E3T+08+gxyfjSStUw5tQwKjRERiMOpZk+G6zD39cC4xeI986/UeuQIblAWtdrUxGlGBi32MLxSkr
ZlVj4y3N308H6dNDPaSLcgujPulkUWqVP9H41ZFwcTIBooGs4Ifq8I7HaeiWov9huEf9xWRBanEP
V0kYIYaPNJtaA1Q4CKRhEWAEP9W6TS32JTxcC2+fFuBsIWae/6eRPeIGrSjmOs2OYe9O4Wwq4XBY
gxKYGKpKL3sYqz3MmcY+jmajaR3Ws33WP8P0AjFOWr/45odOqDjuv7r9QpiSnU0tqna/OTqCEs7X
zuhisDnrOhHd4yrgHPgvPDMVtXIn3vY5C45qCLW4mAp42Q2z3Thgzci0lVL3IfYjT8Q1/JvUEvDl
kAkFJqD8zY81M0+NXc8ZqUxIKS16lyHampe6ceNl2rH6c8sD3TyiwFRUWqTRwFXEQ8Abqrg9+W3Q
kbIZxGggwDaZd/Lg6jciyxTXCcIUAmcrLS4ufadTonHl6LiKD6SIyn8YdJSzqod8rPkvKPTqsKZP
D9Myj4Noc4dZe3LB43FlfB/FGpHJvEfl2WJhVrKsv6O24AMrHgCEdJ/qgJRtekGJQ1HlPdbpt4BF
LV8CPgPnuQx6X/1biqzxURQp/MXBSAorRwZmd52qJT1juaawVtX1Jl57mhQ5D+z6L1c0sPQv58tX
DkEfvraZRMCfW5R2lHpRyGnMh6pVdJjx1pDhtzfanFPBnMpWhxv++vIry8/1UjwXA/PtTD0XSMAe
XBMJ3XpFFppJPIJmvUGIe9wmG/axDg9D1H+73N/mxuDJYk4C5vl2pAK15NM5iZqH+eSoTLbtTJfT
PpoG/IMniG7twSU/tFXAaQyJ8dQuCM5yuIjN6zG+WrGMM7n2xmCd1NFNSsXlSrv3HI8vQCFcA7b0
XQBeXmeJ35H8jXkFlj7LwLspfFC220hVRFfVmHA3+fr9X+kihmMueqGiKTKHd0Lpf1FuOQIY2kqi
YgisvyHdn7hbNCQvuL7m7Cz1yP7NfG2AEus4dq4/Lsv0exiWTBCIZil0udMEFPQvToFLtMG/pvki
aINTCX0d4Q0ynwLmZMcZePpA12eBOfcncY/qyZ79K+/qjQ7ZKYhaF6MLCaR8L/zRjTUGrey5mSue
nb5l87fIbbMdDWS/HiDYNdNkUNXqS+VvDrFNKOOIUWtQaY0QaFbnltTIAWuXXqKMn6ahS0MmSjo0
qZezyt7Kr0AGsVKVjpGIef3vBSpz/FKCMo0ARdBSrndFnYI4i/rit/1kC82pkx6VsRGn1SUQEZmu
bXW8BcFgABZzDHKOutGHLMnOeAjUvSZsriLGqCgcN0XAfKZwgMAy8qKyhwYMNeaotTotkrI1HSUU
VLetFEzUv4j3GrNbXpCllwoT0F7Ob0HM6xk22OrkOrsFOaDMwRdcgMYt7riv8B8oRxJlR0L9JP2F
Khg1no1Z4lQdlIpwOmLUvmy9GPk9Wa9jYiHS/WeyPjcvmF2hqSgVcssJm9S4HIdH3a/9XGQqbtjP
rBXmE5IF/fKmKCwglBHShsZOJKrxZZbf7LvoaxddjP/eUbNeglYCZtG9bZoll9RRuhSC6ygSMmZf
9Gy+lJNFvjIozvJ6j09cnnBjohHFRHJVZKQ4NCxJMRmFyzKK+rk/DAXUIYNm4Q5Ncw8FWahxCPfY
bYPxjyGZKWvD6dR62XekSoTacq79bpunmHgdtZfxi5VPp3z0tfNLBVdRYhip2VLTK9wHSkRSNLZJ
LC1P5yYG6RhQPAOf7s/pV9Eq/tUnBLbhI38/8Z8YX6YbaLhn6LEJbs8wHHsI6gicjPS61olFLdk3
7/kyeKfNjJo+RQsqNf6iR92xn7MBzJVaVVPoz4TxsSTUT4+3DZ8gTklqrVuYTtsu8a7S8vNDM6ar
F1+jtfHAujjimXA/qWV7+x0x+DdgVGputiIfwYvlUY/1QuqIvkcPDtTwKp686eXx00cy8feGaCZK
KwLrjzmT/gFD2cdqZCKl9Ryy6Ow5FvRLfevREzSh8k159EA5FpbIrrp7Q7sS7+cu3tH+VoYlLS15
NjUo1SqAU2jLmQ2h2i8tK3ynjgNz3xWqTA2G/NTWnPqIBHrRUILZwzpwHrTAcWfONipc4v7A6zJc
cF2WYKnBgtk9zehLyRUKpcl+SBuchTWqjXjurEaPUDH2uvB1+WUZoFVVXt4l7iVjl42iMXJ+9Kd1
+Jgg9/jeHsMNbVEJ8LZii8cNgkIL9Ag3cVa1rDt/zKm9iBbKvUyMEyja2Y6qVUTsbO6j4L1dzsZx
2AxCHEUVFlkQRa5+JOw5HVoLpqSen/US/IJx5ciqnUp94Bmgl/vAi2tU/sh2cPxFN65nXKuywkTy
mnCXyrFsNmD93+M9lDQTM38nXZS0W3u4a5fdY6bhmwhhv+H7c6eE0aYhG9ZqnoHaLtg7RuH1lsPJ
VXrz/vxSsgHxlGpX2Wo9+D4O0WoYWq7feExzhk1BvpfhdxKOdfTj5CCkiuZCBKa+M8L4W/5iog3T
S1LnJtboJCYF9RTEINQiuOVB5asjQ91KoVh6BVZWY4N+K0kjqp1GwNz+x+hFx2alO3FXM7QTSvEt
hRZaQERZBEkYlNzJ32imlpK1Ct+VUpXkcMDq5Drfpf6pgBAQTKcHvsbPhZJk4w0PIXg8XAofIo1a
3OO6dKl0eZnfYDTgJDCNZE4C0TMfEcV6uurCPWgVCAR/6BryxN+GF05R7MR9sEMxLKAzXzHjl1bC
cWRps04WuCncJ2Jpkbcrf1+nPtrpGWR5P3Hh77YoNn6VyL9Y4JQhQA5IvMv2MbexFCOkrLU8zesX
L/UTPIQooNgWyRIqm5tj+N2U5Q98+FcgcnhpK9vOt9anFgX6PL+L/KpIA+XVdJpPuuLzkHoaNTbo
ja6bOzAdcM/DfqMkdB+OBkEciS8woSyPKlhZP/HWIbTgfN/sjZFRG8Uk472clVginge6ukpucQ8T
obpa8jWQf9kWprXj7KJs5zmmGdcvLVWdRagJjz9v2kDjXi4tD9nWpaNOudYvWgG7PAlt+K82ypaP
ehmgdnODA1obRSvz1kvdb+1mFG3WBvwMu/gzF9aFf6j0bQYOS74FGVD5TaYQa8i3tH1lHIrFlnWR
vgK9C4/vw7KvQP/LkXYc/sKVpOAt4d535lSgFNiFN0YrGGTsmxIcXVD5B2ga4kL/uKrT/PIx1deg
5ZdpCT7Zl4cbYdSsagu2x8boXX/MOXXn6Go2cdz0qbIvsrqyyhIX8UlW1a1ty94VBONLvq/kH5+j
iEyGYIrgTDV22L/QDSQfgDyNlejun00+Jc/+V06ptLJ/XMzTztgm2XNqpFGmnoK+JNbSVsz48YoZ
CVdjgwu35JTdQGGTH36pvoRVFWwlYU+eDngNTGx46ghD4LSRTc6xGLI7I1TUQ8Q4Y+QQYxWnqih4
dK2M5MW7MIlXY5yXVIqL80m8cwAH6MHpdCBzgFx5w/5YTrAwQUuoI1Lm2PyLTKsk5AfCmNEB6dxl
tqSei9sW43ICCGLlx3CkNfrUqWP/BIdS60CSWLX9oL0N+EP0/Cvyk+ngRAb5ikKNtLuYMiO1Fz6B
SL6AMVIwIUljdWnaZueUF8zM+57tRtVJ+Zdn/C8BE4TV6cChTrib1ohH7rI/yOlkBB0/sK+ZC7Ed
x9PDQ+VrBs+277gtLVM6r8U/vbpSMC5swPmN0E+3+VdXKNYVypLeiJh1d1M/MoESEb42h4kxhV2r
ipndGvEp7rIOExGIRszx2TsMpmCVvuCBfe0fbZ4BhYEq/eMKqFpyapXwhlZoJLIUZKHmKk3ReEuO
CIAH14sMNkYzl87IIzBh0GZlQf66gx/4bXi/9OOwt7igs1FYgdX1sp4loqEUi7GSkiwMZcRx77SW
/kEWspzthRNdHhwZ3/IMEeZsj3mD95PEl/1qi3Z4xTs86shrkintKVEdBna+/Hg2iT4HDMYxxAhP
2psKxvub6iQN1e2gPlwJ3AhVMBIB6Q53n2F2vueajWVXHz4gP3WgKSaP84c65ONpzumVGdfHT4NY
ysINK/7ZyATb5JEEfExpLhyuoPFD0ETiRon/Y7Dpv166Lg8dLsI5k8+4Z+k1rdDBIJMEKG/szy9V
8dYpf1BPZkb0Z9JOqPnp+caCa2OFIwxQJEEmBJ1YyY0aC8b5kGYm1CHE3ubtyANiC7vAvwrJ+XXV
5IrmzeSeosE4wrG8sUFJ6MXWDRTBr7Es4zl16J5YFfG1C88ot9iC+jSjpM9vUt+g2h0dUkkRY1dx
KRjEjI2gF83Qfh6zZRh32Z1RsNHyfw+CDXYG1jbpJ0kHxFB+rPB3O4jNhyrP0ZOyXzcGHEy8ZPbn
v1RiGX2Udcx64iigDKN0TyJaZaQnTa+ZJnxN2N5YKMn/2y4L4wkJ5vEucW1GmeHGfS3oO9kuWKiL
2eU0c3FGjEAB/fOtYogPAneCehdfxSsECU5kxDBGGwuLuYi0HS1s1diDBoQ9lxYjbGd8/CguMXFH
keZFN8P7VD6CtUlIATc8v+8lfSoab0bioNAWL7rZ3J6qUFz7unruf9xD21jM1pwsTINllViHS7U0
tVDF1Tg1C5GNHolsMrWKuGZ8Cp86Yn3pgJSDdwh6rmDmUMhPvDthTdsT2Y62y0C7X364CTT3lW21
EJ1TrTFuzymczj81XtIJGEInfF9sTTmaA5BI6XfGiOAsxQTx7kDxfYCqEFneefWR063u/rdPlOg1
pmIyPaRMiP4qMtxXG8O078o5avB4aHRpYaJ2gIPbJt7slE99Z+MdzyO+rEZ8q9bBMMq1qPDF4Xj2
A4mBTkgb7YvL04zJzVp3+GNEjPTO+6T6Scez9xXrkNv5mEFjGEIztvOnT7mQI5mX3aY1SE53+3aI
wdDpPkMnyl+PBPn8zAMM//GDIY4nhGZQZri06a9cnEwshfNvbo+5dNNVSg4zmofumaqhNezUQ99M
fbtIsK2nDVceZturzTOuIKdeVX5uMDBc29Uiny9cB1T2DDFKhBWUuHCbOt4cdc3OPf+gay6suUxm
hYj1bkbD6F9OPGHAvN07dh4dpmBGB5NOnJSi0POf5ZtrybMHoVWLgiqsJApwG0QIArSknuFvziPk
7tnyDCZLqf4esa/2QqR2dUxQn8ztbOt1N8B7qYTmDOgLR9m5AkMMDRqXFAb/j2wrfMxcXm2lGJ3w
M2vkXto5xf3OytUsDVxU5Gk4ZWOGT0gqNyL/o7/DE70IboVMoXF9MoLjZ29JlN5BNd3v5NKvCWMk
3h/4kEho2WCUIDxmmErPkMg9nTSf6+A/SA0rVlmhrPkDpim+w5v/kczbt7hAqnxksuxIjN+tbodG
rIAzvva+E+e6ST7TRci/riAys19CuKuuDwwoP4x2Ufjo7MPqWp0T4Cg15GvxAKxdQ97pm/G07gEt
tAawVSL0FM1oG+uBZINd9JSWVnx7+TwNN6jYVJ8tObS77B1zSIqXh5KumliT11SZajlDClxi8ZSe
BssHkhEpcFhSfYeasVUDbZOU0DCi6s4n6cgXjxtQCPXQvS0lDFCNi/WCmSriWHSMvLh1ucR+BYT4
4KdHOneHpIVRWdlLBbs+8+RzTWL06h27TShnWlTx4QpEmLWd8FxapMtcnUyHMXpz7jpOlqeaNk8U
I5OuvYaqJqeNuvM2GXyAQEGcrLYvaKTtQ8ZRtzxGs33FKmLK6BgZzPHv+raBFwwnaEzMY/BBweP/
iN5nG6B0JjlPTz975dQ56JCTaMHKQwhvBMlYeIRpu3mARu/UeYCC3CV2PEu5N4gBpyue5NVHgbV9
0JHlosq+fK9GWo6f8i9kNoZ6JvOJc7nIa9iMN2cv0qd5WjHiEfQQGnGu/wZl0qBJFh6EFtmezdLt
2FMxREhKK6kO3zIfaBqceAwhBfwceapS63W4VMIJJOFI1mq+7Y1Wxzlm3uSxmFIM8ug9aCSur9cO
kovStC46/5y5/bR0QfRJmdfP6NxXtd7t28M0byN2M5m9pMVP/TL1rZeUgzFP90gKgmztg9NpOFfo
odt588AoCYmTy4ZYRgSCCNEybqmH/3qEKRp1KdCE3jkPpPY7x1ivC/hs3IAsHfk5Ha2FzIo5oUAw
xotYIXOrmJ6hHvFWS1VzFe8Yke3MNPTIlpXAOcr+zVPWgQa0jSRCLBiAPv+UCJyPLa1dSrHdQ8rn
x2bi050ThkRqF7mX3ObaeBQ8LpBUMl5i4ezxY/IHDegUSMj0P4SqbF+aaLexIigcVlaZenlm2vyU
zSKlUoz6Qy/Lv5tjcSmnMWeEpZ2mBwyOEc+Bry+htZ7dYhaos8S145qxnZVtTwOWH05ACPIQHzAP
ycoHMvUZ9UsaEnbjYdJMu3XNMw7drtnYwpdG+/8yO2AZRJbCH035YxFKSq+9vpfUqxDVoSprSuyC
y+y3JWMVuTjqNii3X74OhzYX56976AS+SAsjoE/EV78gEuRTpJns+/poIAIYmfcLTZotJDf88T55
iaUdRqweGLh/ltGL+j1Wgjw1KVgwdndJq/kVolcSWqJHNGbiivSuKW1xmR7YN4I92LmWhMZpvxNj
1moiT7qeyvFBmel36qtifhpNdZY26POgk2XOntSWwGpuQvV+5aIH1whF2i+fEcY5ZyRNz1rL6dbz
Nozhz6O07RHxzY7FnaudEesiHC0QSuxiHEWRzo12rSEczGVT40MocEFarUOq3QaXZdeS/fTAndVe
U0R02IKM9KiwmVtkWYnsqhnODfKuqWMvNjdVT8ZIEfky+31qawWs8qdZaADaIpfaREjVhy1+z4Yc
qIcos8C9mVbJcwCoLhbzzm9Z0/8FqBXWajPLjHevwE1SK8fkCFPE04F7+tL715mpv+mGNQqjZS3f
hZir43FOM9HjUoO1xEW+uhn+DsI9jU4V7VLEuBd3CCwE0/KSZ1SmPUlxfi9u8wwACoUf2NDTvMnc
inDKZwWaq1VchRSalmEqN/N9EXTrh/JlhikfBUKeidUwklfdHtpRF4pt1OIeMXAPIMjuIJ0RysxB
vrzCECyBgm3Umeo3UCgZEsPJ0SYo5uAnbPc8HWU9qjKnbiDnUZdZwWHx1AWcy8ty5godxWAwUgkJ
X6AzweeDW+cxG23cGrPcqW1AkEJqWTOXs9z2b4wBA2qvjjznF5dOB16X1kBtK0ig4waEQ872e2br
gH5cHBPygyz6B1KuFE9viShyoU+xJIREdaURGZWzFsPMz1CMOe501B69/IKxF2xVOIQIPaNPYhRd
gpBe0loInQSSgvSboxePMg6h9i5LZauCaNmHbBgKTnPuP/LCaz/pEAg3hkt1S9J0Aq42fU2psIwA
EWkV/MeOIVp/bze9HqRvj1MVOAjJzd+tl0qAqqmgL1TEd6Oiz1HxJCMMFcfKFJ+0PPqPN0CcWxj3
rqWOv14wbZLqaQptCr7o7WOotulIXBA/8Pv9/CSxIivQYkttEJYzZRDfeVYJKl0MCJApLRc5W8oA
QMNVZq7oUai9ME3yW/KndxE2gQra2cgOsLvn6LYmNLB30dBQQ3yfc2WNKI3AfymydaRLmijf3EHy
aqQD1KODCtFkES4TxuTvGwSCcFUXGutlcoNu8ok3rHvjzB613jSqeIcYCtdvDO6lUuotgCO0kMGj
xzrctNqWD7SlGjzNHWXIuKCFyFlmR+UGKxW0AZZXjl34Dvk0EoRhjptATlbdUroxv1lr/RrwpSN+
EY22fD9qMJNbuvEgxqowXLpaHSUYc8kIcGtmJCpQgKBGmIRwD/ndVMgYE7H0WOZ2rOtKIS0Yj2XS
IRUbObACfjBkdiWDm0zfYW4OqScjiQJvK1xxMXzvOU+KXGIiFfwp7QQbhSvmeZ7GTa4xzTBJGPSQ
3PcE6MoVJk3NWWUNem6AAfjwBpzh2SIwpidRyWCmXNGOHMGaZGpIdhTF96E0XEuEX5TLH6VTySJ9
3uptxtkyNRSRuWV7nfpmlRtJDOHD0PHBIb0ZaFQJau/pqZ7+G0P+7V5LMd8Tba3weVRN47kx/uHd
QdsQr1HIHF/f7fvnjKcHsAXcs+z3nFftwF50VzwygHTtsCOVmfug7LXCjxQ1mUJ61MCT4uIH9aPP
MCYzB/N1YrgCnFDOG9+iCSoaQGo/IFRR3u0mNVZyGFhTIAA1tYKY6LbFIf+NzChfHL7Qf+wDvOkT
IAumZ8iQhRslX4BpgcYQNPh2MT47/rgcXX1UohdfvdzGzKeB65EzQyIIFcMBLyt1tgEt9AWoKV/r
M2/Uz2RGG7XWgou3LGaezGQmEPGXKtiZTob8ooblt56v+Q3iQn8wuntS7nCy8ljReP9m9PwdZju0
NR7VkHtHt65gdT0tJxZYPMf3Fw3KP1WoqgL9H7aMIQOTl9zgw1eX/q5sazJWEU2Wfuqh6Q73fHyZ
3GtpZvP8TicEdtO1OGkml9AvaH2khV7irZYzL3QcYvKDmOKNA6MsQFl6ZDysijZFiUIUdai+FHsT
0R/C57m6RBxb8b8atcq2PMjSEKOB15asouHgZby8kDq2T2lXsPOGQOBF8dPJR4XX36BfYC+fPpTy
fGEGgnhg4WIg30R6soYPGAtsglLvYUfGvH+xDOoPfhZKnuq7iA1Y0tvFXjQCRduzknVPy4eMUs4q
nfanmVBZf+y5e/jjGX8AFk4TdI1aEBqcvBOVVa9Yurmtan7IR7oRj3x/ktEDPaP+FBzCxL0vj8Ry
Ne0yw8bUm45pRDnWDJ7FNJtf6xZHJVrMvD6R6jy4QtQjnC/MKhHACo4yDHXD/g2biR0Lltjr8gGX
BwChxxAGV1+MLZVPI6kt2y+naCIURKtasBuDv97U9VFeMnFnKzYhdBj5mqmWPpJA4Ezeb+YJ2zDI
NtBU5UolvBTRtd7gd9++6KAiXj6kxMSehi1Sam4nj4+yQGsDTGY6gZde5GCrwuWU4IchdQnAUGcv
iw+rIQEvACxnb4BFOqrmJxG9mRE8nqG7M6j/qIkmFYTHr8UiTLBBQ5qSOQa84ZK9m0uU2PAwHWcF
I0YwZ2GcEOug207nUM1pDvEaoWCh5uThvxC2C+Vb4qJ9U9iPfH2EluhjyjQhXERn82K6j5vDrcLv
3rhOMH13E6dve26jPSxAJbXDJWxboHusJRJqo9crQVzRI3ZIX3qcrSkSo6WQP7RAqJsay/f0cuYG
44Y0jmpae71WX8U+tUgJruda0xPKnACJB53zqsh09FGP4NUclV+G4wIm0DCed249i7qu3ZSX+Snx
XpccPIDmVHp7h40K3ZyK0x218mjnS4IOJiv1ZbIDRnEzUtnURM2fosuoN7E1LyTx++nWGOBAkqQC
H0ipK3eZfY0+kuBtZOKNrJwoSVATLxfJ4M+B94c3aNgwN9Lz2mYoG05celt7cvdoid03ntMAVTyS
RV+aXf8HK7oXWhY/vJvJj8+1QMK9isGlu2Q6K9s7JgTSGHIa3KpEvxFJunCwRySa2c6a1aF+pXW7
4cOrpp1C5ybUMRydidJzhOQt/K/ZXVd07hESXm8DhUvO15IwKgScdd5FWk0e3VfBkWZXCtEZMTf8
lFmCWeYgUd+gcJvuUj+5ewZWX7PK4ayMlYKfOMQpr1Ot+4/qtlMQFLf84UH64mXkgHe9RoY2lScc
ZcCDJh0K9RKZaLjQHjE9LIP02KyKpG2NoC6Lb93BgGpy9QdcAxfnu/F/MgePmkVQXXQH8h42wtso
u6Z9XNlG1cIPxIgnqNrfdkjNwWXFmNIXob5ghgzXoCIrTgYv5d3XH5p52VT/5G9k20OsdTA6FEA9
Ttgw+2LvGOdUjYa3LChgwiKG3IpBb3KkyU9xHLEaJdnGHWjWSPGj1karY34QgfbHuhFBWtqWlYgQ
aTPTXbp44KpDSKDplMxhY0Wj4cW5yXGALnR4BL72Sl5hZ4TGpUiKfXCgvyM0bbW/egX0VK17+W/p
+DfqFxhErrZ8pN+Gc5W/lGLvPNvMj/wiSyxBRvbyXh/K/9SW67eVdBq/nX5Agkmur1wTNtxKbneU
gB6ufQbbDVJS18IqUr1NPJeWs5oAC9Wob0NTRXTvNJt7DXvwA1QzJW3vGF+ltmbUx3aunUAOG1kj
WT72DFncZfhaZwJ/UoMWKJwUy23AKqH0xEYs++iVne8BbZVw7Bmz5iDZjoAfFuHEMG/aESJPygku
EfiT4ycES6o0FFdRhgT+FB9S6kaGrL2KhP356mk1EJtOg1tHeC7aWnNvv/BoL9Y0DDZAiMmS/jgJ
B++t+KaJYOHsqoBDqG6mGaiYqL5aTXY+krwjK+OkHSmnynykrhdZEFqTk+Uat4+48J+uIIjeAYck
hT+uQ9jdVziqfnJK1SfLJEgSbJCXi1Nbj7DHW/RJKdFazGO+x1Vyv3QFWlF9BXRMXULxMUESdJvA
zq5GqVEn0Q2R2NlC2YHgfw7z60Kn+TgQ/dWqGi3If3s+5iPFvrTChTTNLPxBfv81pxP/UIK5P9Qj
s2WJzubqEyU6ZVMLMbz1oGiI41qsqi+Js3Qh2b1E5GOpYteMGeab4si62FFWNfwcmqzUN4pKZ7ln
Yp+a/4ls9thYEzadz83lruhWMi4EGDPaxRhIC79Xg/hzmmG06cmAMbpoLegLuo98lmOcMuL5eYB+
WF7UyoaEDMwsFk6ZgwYT4XSkCfOEAESM7QNdwFw//juR1y4IqqtCls7PFQNn/lBU6u8z8EEOo9Qj
KqeTgWnvtB/Jx6J/PX/uTPufZW3r2r86m+vtP+i+dFmxiOkqQ3aEfW7dqf6K8L6aEnXJAtq6xVSw
V9w9zF8jyUt5Y/c8rcUyYUPCAawGPjQOojO36ZvuobH0KDigpL7A2VZyJyr19pGd/Cbv2bZqiHoR
f7g40V4O3jf4tmY136h8TuLTGhUGF4wmhZWBYFhSlka+aLDX0P9dLULvMBxq+ZBS3ELIilaX3JyF
VWMaj5fnWl2M8GB5SIibABc7/acWIL0q68fjQCIPNS3zKagtyu7uPwdtv+AkTfZxodj2NMF66yYP
gFIQBIKyxEtX9JYK5YLcOJEPfNMw/Ql+sSwFH0NZJq7FwI+93idf2WI+e+Ttvyy+1P3PZL7L5QC+
94nz03i7bZ8DXlxpRfYxFnfszAtyt5r8D9pi82FZ0OPN6Q8bS/EO6efkNF1x1ZibEEwWvJxruYIp
UItqejuZCz1mKvpsXHkK5GkEws9iSKtABCf8mqnqQxihj/s3IGc81usSGXZK74qqmkmfZt9JKEYv
hcuZfr36VuuVNsr62aJrXzBjNg0b2X2ANGzTHm2XQaw+UuKuSCMz8VzLS+BWrmirZEjrGjERrabQ
1biB2BpQU1p9IG3fnBSVm7ovhzUz1hSYt2ogGw0TW2a3VBbkg8DdTVJrgSmPpXZlrxLOjTLfSPoH
u3rv2h5AtcgVeCpEyUcS8BRVrl5xCEqKiM8W2Iwf7/K00NC+2i/3Xa2IfTE/JR0t680NSfqBfzPt
NJkiB+o1f7A5B1vd3dWlaoyoM3JaKaAEYYLtUwwCopxb4TU/+8AfJYwkTzjB5IYfnLNyh6Cmp27P
ZBQ0oNaz2d7F2fAP3ASgV20fk+ZA1/D0bWIDEM/93zDyYd3ek9XtmwT6FPL8WJB4RKD9T1qBfcsj
pZ/aQIjV2GNJ6cdT8fwIE82rIsW2d4tksZZuWAtpN3a30Cjm7GKP/koZgn9NPf34qdi/RhfIN7qy
gdT6haJieA6TX4hE3Ikiq2F0RNbSv/WUe1Uej2GFugKoRRAcoToWjcIfHM/CrL5TCjrWdn22ro+M
77o7L9mBOfQ9d+8VRPOw560vnfE8v2tkAFHrcRxMmb7A1syILa9AuP6a6RjD3fGOCADSqfm9ubVx
ebhhRaQhTlSIDh8kxKh1/nsuFtHeszVsFi2f/5nGPjxzvDV4/iZ/OY/5Odt6oGx0dOOfq/2iHG0b
XkHKdU+XWlZwA2Jr0MUYfn2YU7iNs1tCITzGNuteoNpQ1HiLQQlLivsiPdjoqoCu9EjrpwK6DUqL
aDFmSsY3yId5hNRFBqMwZQa0ROnZwoorwU2e/yUmTJcpj+dDfgyWeawBcqKmRsdyEuqglacKkzSH
ocAv66Ova/x9+cyQ5sI+crnaUjI2MMHGeypAV2v5lEBjBiwXzQWHKwWGw2Tc2uGWGZAYwMaoEBvs
D+d6+Kcvyw3XN5tcKh+roiJLjTnsvxo/YmrNaUZUQkZX5yKEeQtRZOzb64r9Zu6VQunZCNoqcLVr
v00a3KmOhJfQ/Qb38hBefJYw3Gkx/VVGI5Atp+3x6pGz4YeVS13rEOVez2JWMaQ4HF9eaXEYOiXx
kUvdZBcMxZ339mBWKgcAZZtYUQtzjosiqkWoZOZnp1b6/Ktv4sEL+e+8Zuu0YS0SJLeZ5cj5a6Ws
xMz6yeDzZk5I/ZyMbWktp9yD/Ze/G6mMpgArftwiETFpbGtTqExJFNyGFQRUXndgO+qzZqK8/1oN
1kO/2Y9bJGuwuaOgIyU56WxYd2G6gLftYsNx5nIPNW3QJDh9rg2gXhlWHCq9a4QfTykSX7BEtzNJ
CiYLsR+N4GWqKnr6WBjVwFuo7WT85Gj7VxPLKf5UR4OXP9rG74mIixPcEJVZ/2nI5GB99zbzPlfc
Fo/2aCrxAMWEjWFehzhd1smpAPktRdeJNGolZIvnlQR9c7ga+5MPtB44Oz+Cu+hejKOuj9mwUZ7j
896P5Bq2tv8NHYW0+wFeal0F5La1kJgn/o5TW/B5f49EwStoyWSQl1pUN77cKJsNH0mtNtffZ/tr
EaPk7g2BxL7qXBaXmSCiMCUoO+zwYkbQF5tqC6Iyd+QOulVv1gGJ0UK5ttMsL3W1khSvLNicVaZf
64i/AWTMlII/bcIPi6pRft1HqP5l/cRpq7mvS+rofLpS3HDWkS/Ue3UvGrHYbAKNheUqnuBfsbOT
/EbTJLaejo5ZEu6kGCqoVv0ItnrcwC735sPwTdJrZfUXU/oamabiOBTqNvF/WYrlEhvnJyH3raC9
pYQGa3MVGzwM+UWrwBNwUclEBir/eo8Q0RvkgZ3QlZ4lEuZ3MrKhIaM2/VzH8MnHFdI3OfdvMEDo
OjLZL0YnZ2L1qzguhcjBJSa5hyVCICwgpRWveAay4cSdttV6ywdCVuAffKU8LxfF2uNoJUMaPBQI
30FqkAwapYrhTfL5okWkL1diWVg1fcgqn3i4rluPSDHnyEMSGKESGLQDhRGzB5OcsHdiN8i2dXSX
NAfWe8LQTI/i2nsn+Msf8mb/XrlluIlc/SX1tD0qE/JQoswD0AEswNs+6E6Bp0i+RNGcU10TD813
cWqILXMKg8n5a5BPFHPfiYKU6PDpN2b4/xq+RJRt4I8eFWlu0MzUUOUsZaosHYbaKb4C9ou2Me+f
Du1J4nRZx1fSyN7re4e+NY8blBfDnSWLfAgw9BylIMI318fPCf3B7gh/niR/pYq87OGr1hBLb384
imcxxPT6VNNd64/+HGRp7SmqQlh+9S1yTtQ8nF+E0kd+qjkFaXV8oQuXTWzgCKiIYvwkPP4Fh6af
J0B2qjPKmshYTgjyfNt4n5PL8bl6AgCVmaHiEG5rIu0RvUamE5Vgxja/l92VrS1/pDKGqeH5Rajx
O4VFZBu2Uj5oAiRl4etvPmLl6Ev4sOf/bV3eAVk9cycf9HfTGaP3iPIig0fuVN1EvWu+pxCwZiqq
kIhn7gKF0Xj8JWktyqRv5kX610T0o8VH1i0ip99WES0Gf7pB4CPJxM9ufRcqMMVu5JxCvrcH74aN
hF4P6n/zXqq19Xvg+M+iacZcQbnTpSQ5wrbLH5iSurkrwp5ik4VFxx/WNxEoPU53fSx22KvuIRmM
9GpZZqJZ2QJpvdC2onQhfmZWrYmfWe4e80pejTvpfYoM5TUlskTa+Rz5XaWJbNdIj03BruZPbq4p
MzKNWowbTF4VWULXxhUY4S3usXEFw3/LQ360ap07ISbd/UQ++pXlbRMfAV9c/OxvtMxau0dstQYP
/at7DWmbrUSM7gAcP3aUBTxOhP7rxMmeTQlKR2ib1O0I1dwa8HESKT6k4A9qFXnsQvRkeeCeh+yA
3SefaMMCkMSDx+RBDrE2wd4/sWxFXiYykPB19PqQRhZJGYD6L8NJGSXg8nAIc6GIbpPY93MI2nbf
gTFKxMSGzYt5l2p3/3rCmaR5g6XL/oHQwsuPRXrJpVnF24gnMv+MRl1OvShxDPQrA7KR5Ufq1NtQ
pcENoDQFXhWDIXU6/kyBSoJ+iRztm0hLmEl2nC+JNGuwjNRkwgPiqJ6npO5ytMVWJq9NWxX8EhiN
j432Om16EpYgPRrWeaMFfP8Y0UJXK/jMW9PcfoZcCtqEBRlqmwSQzTNedw3PssY0yNq/48RAM0iR
v+Yqlrkc7osKszye8lS+8RrgQ6GjYzop9Q2JHZfMaQNvIVi5ATmT+dYhTYN5Go9WZIzCoEr0bftd
LoRVjQz1iaLDhytIZLpHzt8zk3lsDU4ufbAvulLguzQUvO3b05CN43kxrNsQDQtd8GfNy0xIdlzZ
bri2UiU5O0qe9475FUnnoqlmPruQsFuJMfJkDb8oOvEl7/a55ak+p/xjIEbtVsskymX+CAGDCUJ4
Qxfsyuwc7F8jOYS+U6DTABGX+VcmMkMPS3kCNZBWKJFPEVYegAg879hBf43TjRlR/VpBBs2wX30j
mfQECeSfmN33EqcfnwkXqKuNiN6sbd3caw2C/3izRW4nyF0qcq68jQOT12QuklGDH2+4tTmnFn37
aFH2p1FRDWUPe5oMU+KGyE8b0k4+qC+C+uuZ71pA2OlHCTkYmqv2Gn92Py+Q+bmbAhgoqLMVVvxd
egcS6XUVv540MdnrySiCvev/7/qTmLgbYCaRJzUDYe0yA8lFcQPVCdnVlSMqN5d2mkMT6Az7/YMY
3wrwJiHcS5x7nU9xJFQlGZNMUGHEu3BiYSvYgtfL8RZ2YoIaEpYdXrpyNYCudt4DtmDMga+wpGUl
E9iHLAIqJle8zor37diq2mpetQkD7HR7MdesyLlLYBtk+bYn621nAdx281FMt6qftVJlpdhjhXgV
bqWG8QgThU2gO96uAP9lDnRtUR2oUjs3If8ZumJtjelKx83Ffgx02LkYWD+0tzHuzrcXeR0PU8+M
y1v9XCFahTbbBT9m6igetwaeVCugP+oVQ4ItTbb07LQBc63RSZqwR0CKlBspiGPKSIzr/ZtCo9IE
BW7IbjfZMR7K939gi9Vz1Xs41sfAd26gCXccbnIylSKACiPOu/giyRqzFc20sO5BYc5VEmzjaahO
ac9T+kRBjzl1k8GRDMhGx6oUUmXUt7OJTwqidigsoQEj86Ilp+ByUXzT37TnJmABoMM3cTuJ3v9C
+fLbe3Sjb8k6Mq4w6MCmU9jwzI8S76mVv/E9fHAnXZKpvlIG4bRL0XR0JBubIER7GAngpEI5Gsuw
/hhFDBG+A4h6H7vqWZ+O7YgjYHoQYXtwC2d0db3yiBrsZeNQn72EHgzIy1RUGZeyzXtORshDBOF8
tX6SkyeRp2FqAQgyZLPUMQU1GyCUDy/2de9+c5bP8qYLcfLpjz8RgEbikbPruan0he7USog5i7lD
iN41gD4x40YYiGQYGUE1MlI0mUKFSlhvS+OZHXuozX+8AJwhhO4f6PUbREo9kt3TFF6V5SMtQFc0
DSuTkmUTtfEIIb5mJ+XFBsuRAmyzagHkzfylNoqog/iwIzlziCCKZGwrmwkLtDBdt7P7hDnpUF8K
lMYTPyrbtPQAZEGP6mXi7WFgzYOz4Z0zpncqfLK/jljMKMP9F7LoEm7iw5LEO/5plcp+2WVQxtJb
Yo1l/nmD8SgCKfEXn6unXNiBoXpUvsLE+48yABDXVtaSaQmBV10p2Z0pusgwBRWcvrtjaAixz3OL
j43dRp+KNNv91TCSWsxWgB8ezXhJJ6tGs9ggip+tRlvrYeqG6gu/K262eugg/GL6d+BgQsSWWOXs
zymDcNKM+J44zWWkFQBf62mfQaLe/A0gls8XCgRutmgwVWjwTU0DOHuyL7mf2e5PaqUAl7L9A2If
BZOwCxe3IJguRBtwmWfCBxumAV/mOy33yNkPtFctFNfT62z8/9G/33Gsd7rZSAQfuDbGXzoRChsW
0dXrT+3fbAegr1KxLsyHD2NYChBuJsO0smCwDzyGJrV+RgTXfS8cVd61CBaCmGkvk0/AZ2vYLJ08
Nuugrd/OCMWwHGuuDquw4BIgnr3jDWJtkOGgJBTfTdDc+m0q+8AF9aDbiEktM3JSd2Vu1Ka7Os//
40e/WR/uvMhqkMtdk0c5MszFt0spBr0qN1Vlh+LN8BjHRFsSh/HcuEPI46y8D64LK6xelkf58Gm2
tlmiqspp3YRKfK0tP4hUyS/pWtG+FebDUD2b5vFEL3HRBA4alX+++/eh0/ULqXpS3pUmhgRpKJNn
5LCtDaLzTfjSFvDTWqQi6aoN98ZJ/D50dn7OxpINDpLLrlnjhTaEP+N5M4G6hhlnd5sl9CcO1Pgk
MY6f9cr7IHHdFy3Fe79dlaoTIjgUU3nfPt4YDrxUu+RqraTAwXm94PgX2PtKQ45rBJUKKwccqVJ6
6DinxTjGEhAFKqPWtIf3oX4AO6vz925RPzS2/oX34WTZibLUKzxclvZbOu6GSc+o0ucFvI7Eh8WH
qw07x6n5PLHSlLlFYu7i6JtuNPFFDVQ5bGUrpEtBKtGi38+uUNzCJI46Fe6Ab8EJ+ScrNvmKTDQe
Ahgrvn84dho2YNZaEJWwsr5L/hPzfbXpXJwcT+eLAN7ElsvHfcb8fUFlSHPs3dM93AS+VJiQXhkh
U1a85GcEhv3fUtCgAdknj2Gtun8UCaYnq27VfwUnaudzqskvu5gXpgpXdipVHdau0/oO/xcjflKo
L5ITVnuGonG1s7bytKEiPQG6bAZF6xrqTBsFFIm2DBgG+K0N+xn5zGylAOW1AnhZU7oKw3pXBak4
UuDjeQFZyDpvCP97w9nAzeb4ld43ukEIgno2u73mcQpWeAU/C+HVxpZvG9n9GEtzuRc3muyhzSGr
b2/WfwfcwIdznacpb2tZ3DVJiapBlJS76BtDbTX8CFRfv1ftlLzs461YT4XYoKMRBt7lr2SbXRRO
Vjo8YjXTv3ZXUHlUiPHQBS8aAgsDlgtV9HqNk3WIV/HnT7ruIUJkLHzj4nC8+Jw2bu9ogHrDP7Fw
osae9l7nm15EYZU7kYZrUAFy/Bh2mSRNjd/qreY60aiFOuqv/bjeU0CpzvFF8HskB52ggxeIivOJ
ljlRm+vKoEpFG04uEETKL/w/va63/oBBvFw5z+mzRgRwCN205xNui7c0Gf0ySvFgHbFTtrtAEqp2
ZjCr2QDzSqUg1S2FbV9WRtudaphBgCbItQabUGqO9L8AQZDoCI5LDwHdAIXZaNJzqilBPBnBoz1H
6onaYzdBFY3fVYQl63FGUvWZo2d4SXub1nozt/v4V0pRuYooIAmN/Ay3+6hLHA6HUCt2bPoZsQIs
N2/ge4vmSgj0/ct7UEZ/jwZ4IcEFAr0WAttYoGzHyaig5PTmxfk1gOZFTfTSuSFpZdc9Odrr1HA+
k3Y+ubArF8EaXt9PdYnLsxuRUNQm0qio1A42+N4vbLB+KvsVVvSv2exT8WOSudI+ku61mfZhTfnQ
YYCO1tQcFRfeGtfv9jJPul06RVVr2IgaOBPsWRoFF8KMXu7KXezf0QPZj/Tbm5YSfYCP4Y5YWg9i
/ie9XX0WdcIbXAbkxkE5l0iexDmIt1ru1uc2YiSoGwnOnDLIPRqBMKnMF5WSUcp1bYB9BF6G44wz
sL8NzfwpXQWLEz12jL9H0DWxHtwkGCau9q0QbpL5CkgQ4w2oY+NhFlUALN2iTPDagH4YV0MLsvWs
+MYwGvQMqKR5CdeG0y0FR5Ml5P1B8Ml10A787Gm2aNUL6MSC7Hoxt1/fyA2QqQ9CVrFOwThJtSbh
N+GqXXfBx0xIumDpmOXMjkGLMvY78szh86WqdrwRzyfUtprI9RnbN1nxRaQSfkcBxziyeC1el7nJ
+liILjyjr+BP6QAm84P14mIODjMhLaJ1IRdfECGSbr/fXc/qbk6kL4XhKPkQlQgC2puWmIf3Zg1e
8QGAiJo2NqKbSNHsO/jlyip0ou2QE+MSSiZ3TwzCFZBSfA32oQrhBj4AEK0u3VFfTCC5/YCtQT7w
jTcn4q4zYUkig9yZJsefTfS1LXiCd2kx+grHJocXdAiAzXIq52zcKLxZZW2GmJr9Z51uPHQ4f+ZI
rr4VgixEqQh7TbbxzKwIIm9RE13Ue320SdrcRfU2DlUw2n95F+J74peN5RvUcZAEmIHratNB7C6h
GyWznLJR0dWFK2ySLWTQmIEKG6nl+vWHg0pUoFVjRH888ER4PaD7wwvmQmodPONFYbOKfiJmqg7A
4zJXoSOGsW6fg5pqNSu6AYxpvRE9XSP6yF+rFXfKk7RSDU4Gz0dRTMvleK20kNAjRdXBXSkanX0G
yrY2QdQyOC3EJI3JI3ExOiwa8bkEDq3FuyNV+JIDoQJfEFXX/UgzcktntRlZiouuLzUTpSdjbFoW
sT1m5dshtnZsMlzJBgBDJFWVw92w4sWljUwFUNWmkeWKmYGgn3tF4BI+Gvxkb9P+CHE8tC1NeH2j
GG+MSAvzBJ60Pf5G0yycKJL+OeZGFWzdCohj9zoqzlvJ0UaiZwiHl89CN8yS5Yk+8zYatAKH/2E2
h9OllJ+57ldBuDp2ZLvoJmoLv87nsq6LMOqU7B7Z65j7P5j2qLPWhP16Lo40LtihfBfPFXLcLpmn
xQL9S9fqkaLCzJedMtC41ossVHDHhOMO9N/nYfgo70ycrKoIejVEMt9U7+Mtr0w82VOwM+7vLhv9
Zr7SMf92dYVGHSWXVgIL2TdNxGVuT4qjF4dlAzj/SehXbRNNedyVoTbNheCayzuJPLyQVimzGEjb
2ONuXqbFSM6hjUqp1cEEayemmAdFdzRz7vANz+tzYTNBiqH4aIe+vH9GSoozzfVvtSwo1SzQIlJd
faftHSSIfgSXby+UvbKh46DVZUtSiJzCkS8hnVDdK2QrG5Z9M7KFwXvWcuDC5gPen42/he0Bd93B
M7/bpirSpVy7yapGZ2LJOpqJT+fIwreQnxiJRfpvFBumCAO1fggwxIo+iPSitPDiobCSO0kUp8qN
iaFGO1h5Rc2agXBtnSJqX4EDLImUqw9CRsdTB5ogNsIylJBcW8/gmC/8YPAwnJVSZ39ERDPQDqYN
3h6hzMEjZYQ2m2U0653+pYDZjasPv4Hk3JmWT7D0qFMPd+k0vXMsqO2JnTncNwgYdD+SCwv3vKLZ
xfcHZS5myi9VBKzGgy0ati3K+1hXOfEySWVhTTvlN+NDRMKvk3h2A+CA7kG5tnD8dE5lSVSl7jGL
VI3mP6h90+DPX6VRqsQmB2UVoJ0T2Mb+Fd6v7dQNLMbEasq1PTCJ6urMAiJe0TFVLq2CCaVkikog
ob9+LxQiW2WdGrMxNr99fJF+ze09ZH/ZHWC7/f7+tStvzZhSolfVbOyp60x0FxeUOjFWN8PErpG7
UlK7mTEdHMitaIoRUmlfW0G1HeeHbdwiyQZV4f6DjG3qGptelV6Xz2QZIEnbisGa4CVwXgKDyxTe
bZopJEeJoqeKG6p+/k/pIGV8MQo+iMLTglnQAiACjjBrtX15/KhhMYuewR312OO9pVDk4nsGquEl
zoiugiZnxHIvLcLkmYSlTEv+6FwyRTrwuhxedd8waFFEvlrSEVAWA1rP5IGEjoOGVUIQu0IqsCl9
9TVVyryQMEXYxz0Hj2HKXKcQr21CLYteMsYN499ISDm9fuOgIn+SI5uo2SkBNqK1glu1bZQlVSCt
tZidpPt6fQ+2Ql6nQTkqEF+prMg0f8rATabmMkuqorwnKV0PTFOLXyJQVvfCqC89OVICVgi8ZNbC
dIgGwEVuhgiUR9lH6jCe0/YQt+cDBrWBI9a6GIRl5py1WtbMQ/MDc9xoFTkA7LfVhJcJuzVRsYjP
x1CO0ETl1KaBzUA1vqEByr6xFF0X5yz3enDkKvZ9gdT1ap7uU9+YqP5BLy8CkXkBeScPP/1UQ046
Ox22f8vNnQuNwRcq73DBpnz1q0RiGDst6hE9DUrAS1HfST+a4ctshdkcB7sOt7FQWQq9hF27mNc4
H9Zmn/NJoypyMuUWKP5kqe9gFK8X8rFKdL0oSHEtmg6k+sa99qfSRhruFpw2pZdsaKuXMTxGoD+r
rtIDqOyvIP4rC5Og8hiBImPnk6k29tItU6vo1Zw8uB4P396Yk72ZHj+IoQpTv02HiBwZ50hhxbg8
WhfsXTtCUuV3C2YI+omyNmCL+WHyVMrlNuHZ0qSsqbb6IUM5WuMgDMupYBFCI5U9vPAQQA+MVc5k
fK40nvEIiwb3s3TZStx9SsF9G2lvUhfMBVHNFDp1j9tjU9pK9JeZ9NhQ7EElMK5CKJjRLn8dGvII
9by6FN9UInkidatMJljShPU5ILxGZ8D9KqzE45lTbYAfW3GiM5xoq/3hZ0GDOOWa2uRCaYIdMefu
rBWw5yLZtDWWLCzUuAaXkwYeFu6DsqumJ4Y0o24+LpO/lUmAojCc4yap47rTdn1qYGr6Gp3gAX+R
zfuTv7RVTboH3CchBOOBLrdkfa+Z04igPvyPYfaDnz2e8NXBgogv4fQDZvK2yNfQzN3oo1jU25Aw
kbOeItC1lsoAVQucWgIUVWlkSh24X8o8KW869BaZiAWSE/eCa5sWDbSiDlzr+M4i4wXVb894d9ls
hoDOBLi13677BNd+gRHimxMuoxIVhf8/q14X9AiDLL6byeX5l2PNxjpml4ASsb5v0kmIDzfr50Km
UQhUxzvWOLxv3AAi9UcxzOjV2bzAcypu6pRtZYZa+L8+wWGRWe9gFjS2QQIk+GkGu+msZOWDPFrJ
CFUax/SvEEuboPiFvY6hdfK8BFw3nnYlDqSLH0OIHHdKdzs0iYbf/u5d8dRWpoSz4gB3g3urRDGW
7LvgWJIkLaCeaJaVzElPQEE1GqRCXY6CADYt3iozLqvtUW5b8pE+hXw96uwtQgum1jCGJ7/A2j5i
nq98N02BEsAPdF4ql14X+49A4qYiq+kqlPuYnk4hLkhQolJ7dcpoDsjUS1McQ9d5YNGvgZnpZfnG
hrqcc1Wa0S5vHuiU1KI+w153Z7CNtsbexdGVGw5y++xVClqwooEDkY/J5i4gke+u4iCtV8LZkN4a
gltU10IIQU1/2UpawmsUBLGlL+AwvUFx2HAWYU91csrb+9Z0KCgwDlRCve3xA7S1eCiTBdjT+Gm4
aJ2ojPResUxnGwYDOEi67dlfQehLxv7OYhSV6Ty4i2Wg5PZwrcYpVkbzwNNFHqHB4F7FZWNNvfwN
xa/3vL++QhQjzsufgvIUhKx98pYR30vJwJl4BO61laRIO0OP0EmNqo79V39Rhua0b/Sn5QzQ4SQI
1w/IVJlgP427eezUpR7DtIKAsjNfTCmR1gIneHEvt0QjZGoHJTNKITv2Csq2iGwi2EeQQ7XE6KRu
6ASzxQ4zWLXNljicS2QEZEryOI4QwEuYuvMbeLfTvTD3/Z0rp+cor/SAQxMV5pqUycPhye4b+bDb
PviFrkx80uMflo9H8D0HHj3UQZv/wWMOC7z6yae1i+YNbW58xt6Kv6Bq9AqbicH3fRfJtAO6RM8H
VoVlw0N9im0JGlTumMLlELDzmSUBqxguLVMK3KIx4AmPeYIJzNrnASs2XpuLiEDlZHc8+2ALDNJO
IfSrYsE/tHc2DzhTX2tDRlIWPuesdXmGWKqA3bheSABnhqzCXKa/ULFGCRya9greTZ5aAq+cENyF
xnjlNI1sOnLvNddezVqt8/kuWxhxzCE4VBPvWKaMfG2iPNMoSN1voUwKPO9gNoUipj00ehUJpjyi
lIQq2Cra44SLsrMleFLWm89/8QRXTjyZqWAyNfDyHf5a0R2tFOZH8WBaHwW/MbZhAMcZNugLuk9t
Ah2cckFl69oJaeDT76uuXTGL9xmJY8v99P/2aGHDYBiFEFjOarsswvYzkUxsNdHMz0kWa8xlhpuX
jsKJialBtMlsmf1g61XFYdtWd5vEGtkU7wJr88UsIA8WgUmHVAJ0SnVvcatjWiiFphYIUk7Jr8uk
JvvfOLL1S35rCw3IiGiqxVBUHoUyDtXL2aIwdxXJ0vsl/cjheJ4x+R0esZrbzByRsJ01VMGXhY/2
nqz9XrcmybN9nlxjPGcgCTXHR1oZ7QUFmhcDjT5bCCmUqF4SXRF2lOy4LKuyDiABQbT/bnd5teRd
1YqoN9ImZPLuMINz27i8elbOfWKbAg7yJrBMGd95s24oxxpaKaQPXo03oFCWKrQdsClItLFdDny1
cpkgV1D1rme6jVvHYSBV6s8LqBHu+P0oQCKWl85CiYTkkgGC93OCSpZPb/g/FaB5n2j180iqJNQ5
tKufNbvigB3ySoGjwKgOjRrU1+9h2vU5ASr+no4K82QrHEB8E9pYtrcFY0ubKG0i8mFfK7YpRqad
NLCSvb3+LNsL0JmvIpg3eCoXNyYUZcsQ9AaoOWzkCU3aB31bKIax7HR+Yv9DLjID967Ch0pHxcXN
QLA2z9E0t1HUBTIsDvmOy38WZdr3hzhfQ9EoxIFcLWF9m8A1ui7UlZlo6xJrYw+rfae9MhSgMZML
iJgtexfuqY2ktX6qCTYzyWL7HQeaqY+K54tCRw699UmYWMakppddt/Urs/jeikQsKka1jDmnnkNU
Ig5Bhv9zXpdZHFgCnxTDqXU4fpNSofaStnlseVAaEc2z15IhkW0Wm4QHdk7ArxQNG3LW+GZV5xjO
tfS6Cgb7+x0pskQh35PaPOB/MsrMHYmRndhMPQ9RPADHaz9IUc/jA9jcWnH/db/JLoEdtHCodNBv
tIktuKiI+B9as3D9CDzBAVZEDQGWJLL2k8D7c3T94kdx40MOH8i289NSwpDxuT3AqBIRZwM3jf9h
oajgx/2+RVN2QYQJig7LSaaVa7jm4xU4dUwbwkLqdexsKoFwkBFBNOZjvtzn7HZKFN5+FQ10y4mw
Wxc9qWsHDPGy94AHmOVNoHYcNba9P1oMz/H1mUJP4+S1g9a6Sn9r2OzUCL0iwGG1/7W2YWSqGk6q
FoU8/NpAQ6DQWXE/J9sHHoKA8jrF1MX8LlXBXbfaHL1mhUHNmnoAIYFKbhoMqv3Mdb6+XIR5/y9O
bB6otEmTnHuNerZ+bt5IJTlzsEoIGAcqRKy23HOtcwJdCnmgFE4GpGtZLgoj1/DRYdYjJUoJHwnt
uY5bgJE7txqrwKf0OxNRB8Tlc0DpJf3Lyk/UyRwNIj2KWi1VcJlILhUmOUrz3q9/V9OCi9MgLw86
/HseTNaVuVCD/SC4PmJw2syqUpz+85PeZMasuGm93Otzysov+Kf1iD96hv4DlbIsGi9fnROuowX1
LTXuVlS8NKysL8AAngkA4bmTANC/TocVYKhDlMY20jdTy+QVj8V3sRAm19jIlmym3dsttHMCmy79
YdZZvt+te9DHTYowQMauVMe5uuruAB1XSVUoItpcaoVYZkSz0p4JZHN4dSgWTkV4mMv1CZqNuIrc
dNZGjpNDLQR8UHGM7q118sEg7O96fIEh8NJBhilTb+AWqX4bithznrMhxfCTmQ+yZvI57Wyl+Fkt
cReRXhYaYgUHUUz6T3y0VNDQfQ7ACdyCz0z9ll8X2GKnStvzHw7h1nEvkBs/y+lA1VbuzyNLEOMd
J0vlqZ6XhPumLcBE4d4LVtN5+Jddx9133VwefzzWG9D3FI5tNnS83SeINd5NwckCglpweqInKkUn
HWpyWPtyFXsH0sVeubfgWbtZJkF4HlEqp/URhKjXaziklU1p6cuvotqb7OY1fudn0bpfuUoVi8p6
/a6gwiEXX3npeCOdJugxyS/9mzOhNjFbd1GEoGdj2ke06lsYIwwBrsMEPx4BQmeucEcQDYLyQIRk
T3qymiNs4WWghiCJY68QmudG+SfV+IIHnT4FC/hHRKR3gYZgayK1Ov/4t75KY7609AVAEx49HSYL
MZjuUTX1BmJDl/RAMKgq9LFkNd37uRMsI+cPK/AmkGsj6xny3kzN4difj63usQgJR3jS3U+mNPZ7
qGFoppT7ix9D8P8kPcPcp5TlgQZZov9GJW8vh8klQ7K5q2yDEvsDuDE66DWrjbrwo3s44hGtfwyU
QxBZnQPtcs5xtcv6R1DZVlW8WKCDaNv7+9K85Ai+sohYUqImwiyEKFCNKYhb/xcQL2rVc76d4bcu
iezF92i/jYtSNo9Kisz3Bqueut1tDl5gwT5LE2nZAnGYSqhohWVuQvgCLwsMaPnYHmHN/comfwmo
mqCrD/46z2V3k8M/fvXALjlncnlnnbkvrZF7Dgadp6tvBruCZ6s1HZ8eTqz13XoJVaqBiHCSM/in
laHcrg9OffIubLAznNBz2TAnFJK1RlinzLvTXTwIbnWq58UvcSX06BG1Y/OUaY3ufZalUMpsb7D5
YSFxWc3ClOwSx7fc7oQ5DA/kHmN3GF+py6fCN71bie7gI1LEaSvuwPtFqEkUXy1kyFBSWl1jYjm2
sSbZ8TA3be4Yc9+ZhSQEV697taOP3i9EYttFKaO6zMwP5QvbBXUtkRKIAf3mDeQzBJaWk4wdeL9V
eR47wP5e8Lt9x/rjY/17poKOAN9fje3krHKxajOb6oIxSX53UloI5VTiXyT4VI+sYJoaNXk56QLC
E2nGclwzpfYpKOY7ta/FufVzfEOSl1e2v8bJdCRFDqXwahBAx1msUHDN3sLLaKlgg1KfmdDuyknG
GSIdISYGailGwcklL2lOqXODYgl578BELStBkEpRLSP+1ui7BQQcYGWUmw4qaKTn5pKszLkNW5k3
i2ZtqLywdyml78SdLs2QYbYTZ4LaYEfUpEldut+49QS8HodxIP5bwIu53pq0rn4AIjLNcRxTb2lX
8+jjGsXG6NF9gOLbynCVjHc9mdoHPkL9haa2cyzQl4+lhIkwHem2+rg1y5MlaSBcaFYgXz6kZM8D
h0PrgVNrNZV5dzTpJpEBtJr0GvPVzn4PIq3gZOwQ2NcZ3KOVGmUs6sYpLYUmYdGPFTHll6oXvgmo
+/KB2uyQbaV3rPlxgdpuGmsxEkBE45A2TjvumiPturZcAyWRLzMQtUyvHMrf5+77kcmIZ899kRAJ
t1k82vDsUdSOzzYSrbtLGHkONnxFHRNFAZj1ZdeQPBfKKL1nyONeLosnneVPM3Nn1hN4ZEX/XuTB
DsA9oZMYkieh+xZIUbSP/3zkCv1OTvDelGPjJfXfWrrko59DnrCSIGDzTtMu8XTXmUpnsqAQvdeL
sHKjBBGX47fMeJF+zLHC0C6xy98WtqXt3XzpASvZNHE/hYfmRM+rDum1aV1CpzFPqKsGbPTwX3Kn
Qpcp0bXDS8zM//RPxLjAa/zd8G/ndXvsxhGQeGj3cWu8n1fjUhdqmCMke2RH/49ceJwTXKi7hPH9
zoQ4395svqg552AJPC8yEEpaczox6sL1w0WRJ+73Unwu+gOt5mZCdzaQac+0AWVOQc7+/797bOU2
WXAg/M/PcWBQe/Bt6LdRRO7gEEehAZ4I2jarnIL0tovCI8YtNFryhJZ/h6U2mSovg2ozxHHhtJ8q
dK8ihBRlC+b6bXoBuxQ32/SUWiaZcco/4+8o1COaP+1GRUsi6H8meNxFY+XqMIP+2xaIowZRb+gy
mhZOO6VHdiRjiClydZcDgBSQkMJIn/l2cZ53rmvS3Sjlfcd7BZRTfz8KBPHV3+owuM8+wbZHya+H
3RrsOEmftOaTBMinS+2wyKKykHZtngW3iPQQzJeuUCjC0XO+RTBBDpIbhYf1hCghqx1MX1VIYgEJ
8hRYCZ9xiwL5JuY0Y1607vkuIfKJAd7MfRq+VQyM/n/PiWIAswMHFcHsDbEnjNMv0hXR3ISZ6QAd
oKhMRM35xStDQoIDgg/0mbku6BnKyY8SYkwfNtOjdiTsm2j+jF3FVRZxuTmZpqpqQ3sRMzsfxfa7
ORvIIVj2VJr3JQjdOIQQ7XrZbyfB8VemnaTmlSwFJVUz0VRcpi+KapqUJmuGOcU0W2PhW74hXqct
XEIz0y1D3liIeEW2wr5TPQ+0D+pqkaajpqfGGNgAg0A48VXlTidxyRoZ/36JfGdTboTbi9a2vk+Z
JeMX2VgYTamBCvjWlnSyj3aXl6qysMonamzGy4l0vTsgGUflMUZcJFhSgxKlVjOfuEcSHwS9bxbh
S3ZbsxOTHdvD5dXYzkSlFd4QYZex8C/RG2QC6UH5VLvT8rmT1jLg9mKWzUitr4A0Ec4nQVhbPfTg
wt8x1W4xTrOAaMCXMPBYXgfkVGx6/p+iq1Okvb8uDnXRrrIuvjrubEIujwMp0XK4091O0c1ibfAg
rQ4UEzqdZBUVc5KqJBX6Rt756f5TByfU2dcIyhUPFegX5JOGH9xnvfKaYIVc72yFXksJhdRJSOdw
vLR9609clb8H7t/UNueDNCwhN6NNxKBOZyGjxhi5HnKQlkX13kQoOL8DhR6D2Fbz2Ft9zJqdZhKA
onXFiBkPhcLcyM6aB2qwlV3OdMPltEtP65/evArDuMmSmYSub9x5g7wD8RKR/Xk8hxl8MtBBsLpN
N2xQzQpGEOAMnkI/rbdOQuCMPYCu/p6zEXgTAbotC71HoXdRSJK0CdBbXW/eVi9XOqr78i66V9ga
SE299wRIMCzfCFIBtKStfmI9N3tYm0bvNF/yBdTWyHGWhhJKLOFfLBNcdpPuDk5H4Z5L4YrCIp6g
20xOnnoEoGqiZhWY9XGRXEgNxpmBpOQMpYr4Gzs/j2xxv56N7EZFYSwewz41CoDNxVPC7ZUdS171
Q2gCUQ2ABb3n/AKORqkMVc+6pbuKyc8lhfSz9/2U6UtnkEqRrqbwJOJZfvb9YG/sLU1jjkbpNcEN
gFUmxeGoU76cZnzrv3Ay53vyMTxtEMv0byeAIuAIc++ECu2Tq26piSGkgG97D7BTXg7LIdNvj2Ff
3CV/VymL56uY59vN6AieHobyfkTY0zofcNGMJ2e5TeH9df3iWvhElrPrvoYHqtqNPmrP1TfQpxmt
t5LnLNEsEei6UY5hR/dXNc2+J5/dBgb4rpR5lwoUNV7Rktm5QR3eCiZY31QFWqC92mGtP1dlbEM1
ZPaxt5RkyesTzx7tQe6hZENp07+s83HDmuG3CVoBJudJS8IlYJ9xRzpu8sZZzGnYDaX6V0QHyMaL
tIuFLFak5SSHl7tNFmoiApMXvT0W4h4LC6BgdaPGpWf3/vJDXfJ5zJ8YvcOIuyn+1cWBBT0j4tds
VcQ+eLyOHo2HsnJMeYsPn2t31+G+0VgaUAkW8oCE/DxJgY55KjCYuUlUivI0zfMqwvl8Bcqgf4L7
HlEOgBIJI1RzAu38wARCewYlkdbKuVRPDaMDqhpzINn4ImOHjN6RY8zxutK5pxJnV780Jv4WvVOd
PXLxmkIjj0O78BSUDnmzzsTlYbe0MbzY8BZJHCw9NLFBJKFyc2H1oI1WTD7Wg37Bwf85ese+9CyG
YOrRcz0doJKsAkwFZfesmxGNXPYYKobN71BL22QCfvGwIsVpJHX40q1qFyKwyCIFLnyXBSkiGURd
MSVsj7bfIk5B6vLvJFFutEqBUPvks9gPnJ9UrBjoatY1GRaceDyWJYch+dtPTe9STpoLWD+E7n82
XHcjA4h3jNdRRoTLU8ikOPW8igWtDcOQOcRZZ42E7jGnEDpv+aQWZEBdzf1o6mjDIeIjFC63YCT0
ItQrv6e8M3FiwqrpHZw95MwzEZnDihl1cYVnlU0gp5Za69LIXBMcgMbQUsqUpC0QpoHFhUU2k7ds
mJLGI23Wb/kviGzI3oHjKM80hh5s+1S9O51HTClnLdgErL4qTspUugvijiu2/NIAhM1dr2QOvg06
aHwAlMSCipl1upTfzSESiGcswaZs3R6avmsTPoFJWebzQF/hcC0otnSuQ5PQaeiX85fzjbisUAwj
9ziuE70ndpJWiROm/68ChZraTW2DZTqMLCfnOGSFZ+3gdVUci92APblpQrzLg3qcNekaF3wQGhN4
4ttzemzsB+bpuvrJSRwduKrRucOE1zh4jNKw9lT0NZQ9qWGeWvtbEDqwgM03/TKNdm1rpWW14EiA
2/o0/c9EGb/vr6msZ0FoEy2o6tYVlRy/nUEKxUg3md96/CQhuq5bvey4lXcniUNn3ygo3QI/b440
BTnfEwcXqc1IU1LaB0HgqPGwt3XeC6OBH868yWP5iQz9w43NxyRuvn4yleXjUQQxIp0SbS6luWgY
nm8syS5BxNYxENMGIY21VDjqOCqE2WwdJ28YkPHwVDgLYp/Tt5z+9W6apoRxkSCg9y1z05NzwiWr
jwm9911nt2Y7fBcz0iQO6+B+zZbwFQUCoIMMb31P7F3JLs/IfwyOC+sCOVqnTa1lFhXUVSwdotbT
AZ2LYWa55JnmCc1DY2IFQZ4lQZfWT35uS9tOsDYYXJ8dp6cFqME2M+CiBUeEcGDpRP8lHn7xmJgb
vEkMvFX4QQ+G1ZAa9Ta7ydfOUDSBqsFgdBm4VSWOxFSqSRiz5x04R3oDM0lHgrFkM15ESx33Mb1R
VRFQWSwptXPH7bLkkw/zk9yfELC/j73gOyUHCamSUyIR6EXIGwIFkf9wVZx1STEEgmAlVos9LAKi
PzQZQ4bw6SPe9WgErhv9xweSoQ19E7hDhZB1zltL7423yAq9s1ialntvsO1zf/WCacMHegmS0Kdu
NVaHIK+Pv6lU9hhp8c2F3iB9Y2r70hADiUE4kVRE24DeQykavcoKXWrZfxQPnnva2482dDwpPALc
smaUZ/JHN/F0odYL0MjZ5SEAusf1gIr1t/Jm4hdG3lKJWLnJeqap/HlW3XBZZcSm+61Waxvkr3Co
iHWBGw0MXysKQ/4RX3XKATfbFpA5EjXdCd4wnmpZMCWphRLGvNpif26oKjlYybapkvpi3b0gau27
hup1XNdaXYlKl+FvrCe6DIu3wqGgifEA625GdXLCgbGXuNuL1BZfzaydkofY4avmlP46OfcuMrF7
Bl8vOizC0QXVtagR7pqDfP/iIxpdhjMpTj+miBAj4pTRiQdHxpo2KEE9ZGylILU0PG08633/FjlW
/dQ/eLM6cgQxq7hVQbUfmk4ltzm5EsCHklQzzo2wfpyk/R219VLSZ97/Hmzoya1jMedt3g1dnt6+
EFjryRmyB3IVSFhfVWYmdqTX4Px0ROZLQDd2HeXPKWkyvecMtPF6TJsUZOEB5fCwttK4OtcJnGqz
OwSVq3WNJoK7EfZooEJhnNHsMSpkfyBiOUMfrBO0Y9ifHff6vOVSvfsBMmuqhxX0bHRJ15VL25lo
2I44HUbnRFEblfS+1bASFR/O3oV1rnaYblbP4i4IgIxy2e/W6wPpp3mPCi5XfkJgzj4sR7cCpq2M
AwP4o4t67JzVINC4VSB/hd/FtJYGHmPu5VXeg6X0hYO3UCPd+kZSUfwKpPAh5cDR3cF7nq4ROHWg
WSePLwN+vQF0spcjkSh2uCIkVw7qrORdOm8yoecy2kIkZVB+9rGS5SyGc3AUIHJRMLiM+r9RCzAH
PzEWWbUJvmQRUMrkfGFM1R9HezeYymrd5FODaH7xR+wTVEhxRoUGtfqxiiuTUoLzipvRxkeJb+/H
hkDwOWlVn+s4qchmf5Mqt2HfqvYUs6OR/+tXBIapv4W9Z7AefYQe15Fjt3GVezsUgtEJu7RDmEyx
IPtEFwQfcUIDeU/EF8EKtr30cX5gEGrMtKwjQv2dxhKytEcprGwALCUuX3Yb4FK9TLxCpc9wSUzi
cNT72UppYMljZWtULTBYuUQV+9Ptlp7su+xRH2l/ZQo5aTIJSXll+5p3AGxGDfVGmLuIOeFVbFKb
A6OSMMHD1M964DBCVGghdiuNsTVZKAxPvZw329JGsFhfSt/ylD2YsDacgNbXK6IyyYUQUute+j2m
SpU/Dliv/oKb6XPDITVopRVHHOZo7Qi/7W6kOvQZtYqE3r6a1NErL41T0DnyiPLBStzrG3xI75Ge
2VZAStfraUA5pxo9EMR6LokMXwDyCzoo2AySPYcZskw3S91/CKge/hrOt2SQGSEYprzQGfl3XekO
6JlskPC999HuyiXxE6gQcSjEVW+6mSe8V4Pf6lIm5vh1fLHMBfV3agnI25e3u3OOlDEl5YlQpUe/
/7J1SPe1sj0Fi709s6XP6IMZXfI2W0OBozpMVev9s7bVpn2Yk5ZmeTTIryc74RJ/yYj8bcUDNIjd
wkDkJLh8i2v9V2FGoQs4feSl7dyaBkPJvKlbbM/NRiDbOmhQkAhE0DtjWHWB8krcYNHotrye9LvN
B8+NgLbyslx0LnJcBhC75Itv6Xz8WyfqPdWXjtbhqa74b45ZuX7atSbtwDXPmQ1dPNXFPqDOKY6V
1HnSnc3zOTL01FoPbdx3pUgnBzu9KR4wGE4vKf80LWO9NAZu02Sp1fr3TZRkQSRCnh1GtWXSlS9b
cN2FYj9LGoOW+YOBu9XGDqbunp+zIFy2ZTUoaYBDxB+6gqj83x+TM4QS9hgNeZjdhkP4/woIRBh2
z1fzLt98m7YoS9CldFT0oASUAsVPWGznSdpw4kAvnKc2Q6W6DmRJ4VCoLfp/WmV5sQftDW5VuQH2
vcuE0x5+2Liu2zPgniW/Rzs7NeaRContyeZjM4hl/dA5G1opbjO4a5uXzVbslIbQFl/dH6yO6QkW
4ikXPH4nkn+L5EEuFx2q3ty8wTKvN4YR4Hf+GtW03U6SqWEpUBLXjxPGaG1ENctj5pXnrAXnG1xP
Ol5gkVk9GeJVJFSum+fkC8+BJEfv5ICnVBCpRAcrs8QPjcKuCXDR1ss1J10PUM+teqE4PVn7szZV
+/o1VRhvQkxnjo1ReDp/n2hnziTU5t5SQhwZkT3HCENRZMXpy9582axthpgZh3s701kRBo2WQciL
h+WC+WciviG/RD0HbNRCGQlGAmTFBsF3JhypKGH08rJm11jImNMrBw0llcg2pzLfA/wnww1GUFlh
F8HOKzBNuasSa42nkPrdVyD28jMPr64bfAVTlhhy3hKdlhKc+iKVcovgQL+qFnPtdw8WhIX/sV1e
tE9akSrjGlim7f8qG11JNHgZokkQUBFpcEgHzt/LGXZ/rkAiYGaqFojk+G5B0ytqaXtdScZ0XMan
uw9cSogm0Hdqv1MVKIL2RpVIOSOERw8tP3bZYN/f0PjPBSiLH8fCzw85URgILdOe5mdl5JH9yW8/
OrlqgKL/KqdzYShDn8RYsxPt5zVVm+1s+d6mg3GRWi7COKlNDrNqXRB4iq6lkfh78D1MAx0jwydz
ZmT4+QCXRnxiQg1Bh/3Hzm0bp7Jlan26i8v6wU/vEFpzW/D9BiC04492iC0WgHNuG9xwwqeV1qO4
pCmruQr0B/J23Cxh+TKKpJVj04GY40uwlt1JybzNMrQUhEa3GWMoS7d0Hu3Qufez9jNxRG0vpXPc
j8Gr7yJpx11xaCaIQy3EiUDFYfs310rfeMakWGgIyN9ifesObmz1rjoyRXZahYOvRUutsfhyL7jC
s7wVJ6aulDu+aQzkxnWi3wyUWT/R1Vg/RFl+0zc2Yx8mXIhqhkmVNDTy1uJHBDFvoCCWFEK1KqVB
SkSR7Z4oa1qO8SQZ11iODDV3vfWV2TgN5QUk7wbzAT9FfiPmfUQI9bdtMd4tCG21Zo7zlN6Wfbw4
jqJfmkGpfzyU1b6816bCpEXarcuzLad5hBFmtOXRHuOEBqA3+SZx2QaO2XgXw/uKPayOtaWtV/05
mvigqfIY9y6lgLyI5OaF96HBTlf3w/S+oPdK1jN9jtLmBhPy23HzoE6qhex4TwlE5Lv3iOjKEFuV
MP9GPgafjBFGkYeZt1vlMn1AHKPs+e6VfnYhLy0hufwEKVWLrQYF+77oCYy9NpKb8efRzUWv6aqY
m7RTbKI+t8YMeC0YDEuD3m+2uxUEPbVPLA1E/jnwktU3h/v4dtImitIjQW85n0xsQQDBI8L60bqe
nhoXEIYV7wEsGVBr3+W2fRPrDsczrBMWveP6lEJya7kiKu4N6DKszAjyxbQLac85VYO78vbYQK9E
Hg47c9o6nFpVqTnAynMeNTSMfsko6KeXobGPOqIxJLpLfk5XpjAa6dsbmGQvMuNyWxNFqIn0V39q
65oVXWzgNsOP3o4Is7+3sDnB9qWQwRj4JC53ncqdwKD/vcyPmqqiaW0aBh2b4kj7C68mQa8xiiWg
KEL5hl7fEM18tyyNeORsHERGE8mE63DCg2w2N6arJF4ENZPfuJFeSL5i5dCHrHMcvlp5ieMTWbsQ
KF+O5h05wUFoqxd5mMLBCNhnQ1P+2ieooLHnD0vQrGL3KUz3IVTSshr3KgCOntULrgABdlAGCYGA
cFsyZQuWobmpeSzW2YvROewh5/7QojrNAS0Q6O8mgLvDvHl3y36sXYa2ZrhsZKlBNgqCXLC2GOcg
Eu9CBjX+N8mMDow3FvEmXRvInAEVmxE3SuY8MJZI48+jIoYxWP33MCbzl7QCu57MZ4aOvOKhvCJl
KtVpm2rLvbf+SsR8ExSYP8k8xCP6Ed2eVhaw5XlQzF5aQ7KXJANWTddujG3vhXOULA7a1jCP24Dn
5cJ6v1erLyhQeR4NAgjKwKMwkWVMa8AkgEw6wt7x0mIYdvBipS6L0QcIycaV+tnwYobpZsKgY1NX
XTrap8x9gxC4D36suoUlEZNV1TNnxzxNWuckDj6mqtNkae5A0Z0kQplDjB9NIJX4iargBubOdPqd
05jhX07U87tn+g2hyhQrIeMeFA/N9q1+0YQE3BL87WPjTX9u92eQYVVbZrfeSxTByQnzOSckiF0e
A6RlrK6AiL8UYjOOmXVjzpoTDSS5xfrF9PlmcVHWyckMVQOY0i7+5szTc+0XYSX/+3HR+LTbLTOl
VOlUzEUPzThxoLlWzp+479BmKTxTjCNmK8ClU6UgYUmerh8iIlw//jQpnr7sUo95UPURKuuE6uWr
Dd0k4VvbBxub0eELOBBv08BmRyV3jVSwJGGQ/ue/5esEiA1eGtGbY7whNwLIOJbOp1YV+2glO9Zf
Aj3aXMVOIPkTPALlSYUBstLhaHIr0N0so5E79Hf7vUlkV6P6VUmXshMy+wwnu7AkTu3ikIMsZrRX
IiGYj769VQkKVQTTHqnSuR8qhB7xtvf7oo3FmlwjM+Kcw6pVu0JzCUb1wb56MSXNerKxZg648+vX
9tDSu7WnJ3DgXBRUimVD5TJ8pWwsOyovpQ+AOfsKzXiT0MaqxViUks+QT+v0NlCLF1Csa0ZIRy9g
6JmEjdWt/ynNOD8X2ol/zcV94HE/eeEk8dU/Px2WAcv1uGe1x6/W5c9kqkCMpui+jkwDmYx/yzxs
pgUjMmqYPt2s0BxEo1TKk0Cjd+TafboL2IhpRRwnbFFQe9J0TsQ4fGxwTAm10Ch6ediGMV1K7bpT
JMk8Js1DUPGwtrm67Ur7VLNfdobChxJQh4y6brTaj+Ig/V24NkY3Kh/KiCQ1mBfDhWu7spQ5CJGf
M/cqi0AqkmBk7PAPGecT0rzFriWK95Ot35XOVWroJTP0D7wisn2EMLlUYsHv10ff4tJN7tFK5w/0
4PEbhH+LxYYlqHz20WZPbpLB3SQwAfmjLfxAXALMU37Y38xZBXTo1yxOALhwSbj4mhg2y7MM+Vaz
IbuOoE7CH1g8TWFviSTS3C29OnP4ll/rywiSZX3cEJCYkSXKsgu9clU1U7SsiQBmnFBig+w2GTy1
XqMiYpoGmo/IA1niMmzQV3iHTxdSX+cH2+R3h7nIa/52zsRMBqbe7xR1elYUETe4vkX0iuhEtv53
D1YnZLoEiFHjuP20OX632agtK2K8CxoGbPT90ppYU57fYIprMByfkzzS8arc3ZOAapQ/qLTSBKXU
4QRQtjvYMpsZZw0Fcg/FCp9Qdq4YJctSvsADQOnPX/4gSR0VN9k3qlGR5x8b9hmuRmIQgOKnQ0tu
ZR2OOfVcO2XZEJMtfzyqmuSm32qcyeSoPb7dpQYp9flCMix7RTKDy97X6lmOpKaASUfwUpwIWl1D
/I4QL0z/tdqvXpAYQKKOG+00x/tcolQt3ay4Qqi0SKy+kYqINmbWHEn3v9/GLJj+lUyUkWWyRY9L
x4jq+rTF7b0OGv1pxLpqeAjUx5b9ui4BTHVn6bkk8e2hTgNL3pBleOx2g3zPCPgEe5M1X8sozLuW
WTFnJhoEOBb2y9l+QAInd/DAK/ahTxmLlqbRKpwlmmvpMOghNv54iy/BhP4YlyVhmLHXuc4ImdbG
uNMqztDD/GO7fzxIasyn1CV50VOYt8kG1wkBRy85b3vtLjhbvesZPQiaTkTZgI1TIJQsfLyrx+a0
a9UJe1b4moyqtZiAnbUK6Kyzu034fvvWppD8YLP5SRyWtZWVPRG1X7z8TPZDJKatHlGPVUi+ESvR
36MW9LLxs8/xIbk4+D0NgyYggeCuaH+kKevdcxfnL8kNbcbDEVtpv2CESiwfy9jnvYvvWlO4/GzI
hharHBNEM+/kiS5MOndzARnPssaRPtXOHZn65gb3Z8wlc7HC4QA718RT/3fkfxCForI5UWVQUb07
nZ0Spzf5aOFEwjcfh1sJKDoJ1Z7xviNROvAtoxN8K/NT8nE1dSUTddDOcfoHzIDX+dZZ/d6q0a3I
Hx8ZR7K6wsMg/rHRKSpTPH1oHZpfqpl/diBHyxbkJRGVzDFwQa5OKm6YDpQ+f+DbM5OxmXcuJM18
Fl/hBTG/YFpAeO9PI2escbiMtl7sJw5gp3cr5b4MDXvPml5qlmLeFe1W3NC1K3oG5qbMjuKWX5yf
xQ9kSNKo5qFcstOL11Qjttaeyo4GII+7NdC5R1MOlfANsFwiFBp5o16JAebtzS7qxRYOZ+jIxY7m
FVkXiWCDGdBB+Uuy7SXJOAX+u2zcXxONWI5ykPBm2mjesGyruQTmuStFUNoLzN+/dLIYYqscj56C
QcLwLpBQhDJAq83VbyQCML1gei8xn4z3sv/ucIn09JuLIS0jAE7Kf5llF5ckH57+ilYI/WlKBqIZ
AZZOPLgb2qCPkx1UBbZ/X8YqUNN9I6WEB/pbk3I0CHNquBZgxhsvMmp6fJzB6om3chyPfqGf8CK2
a27Sh1qzyX29tnfAdFzyTCZ7YiLnXOLoJ2Pw0e1igKmbFvbmxfxGnxqwqUkYbtr4Zg3vgVnK3PDz
9Blg9M9YL0fMpZ730z0qRN2Nx+CagIiUq4sMRl4sE3XwRIaZfAJYVDnQ5/MS+qiboujaSCE0yjOl
KPJQjUjBDn3EAUfVmKj94KYRUaXZKVuGdvMuKIyM1UO2B2wDNfMymgl3gadfWK7PXURf5jZPaaEf
aU9gnz2By3iaIzvTB5grHJcVes5n9kea2Oo1iAOAQ6UET7Cdt+8sE37DG6BmAygWkpcdoqyfW5UW
IDpg366/qYbvC/TAUBL+CQpG+6gRdbH6I2tG2+5jnZudDEeOMD0gNPNM7yG5UXcevcmlROyc7zjh
sCUuUF+b41R/etRPqSzyBE1rl9rLjJYWoepWT7RugfNsiQWGeII/UTi/lMO1q7s3pu/PkFp72GfQ
ne6qgehwXYaokL0Ko9tGaOTzTF4AZXvbFtpRr07B+6hbWcjjoWzSgajASqRGMnzISUy0/jTJhNa9
kJ73WmQZdfWkMM2dVGig0RrUV3Y/csebtcim907yNK7VYXJkuO+4sRRmaGl7pFImGpPd8zNGkFMX
m2coqn1sYs3hD/TRZFAGgq0qoOSGi9NGE62hMtZ2BAAppq2ZBzBP19YXptwCAEPROQgz7uGQaYtb
0bZg3hbHuD6ntRwjQlsJNqNnpKReYQAWt6hBwKMjQCdPSd0XpSrMcGvz6s+1soFrq7EavR3CkBbR
a33dJrNxO7DfDj4UySVLnAH8nviSmls3ZZrfDKirQ+YWElIxDobj+N10RnHBJuUzynFKhogT+QSJ
I6q87hn/qpZtRffn5mK8ElzsUjrMA176uimMbJ2GiYYHJp94mTyMVKg30zIkrXC1KXf5A84X2c49
QkjW/DyU7yCSrXEvoKKynLO/NZ1kzg2Z/8MkIeKGuc5aEJMwlBQEtlIang2hjK4Y2b8IHpEym1nj
y1wqGauiAqLh87pyRIv0f+d4O13/+qCOF3yoRMQi0cNhpnjHopyWWHXTZCyk1WjCWmYmut0lADLn
n4/uHTZB/VNRtoCpppTWP+aA3sUrSWensVN+7pnGBhZfN6+e2Ppk3c2u+ndnY1PL2gcnTE75PC72
S2Y7fuF+/ztQG2KGjlnAp4BLzLhmNx5fUGu386FETys66yatAoE2sRZt5GldQGX272C5TSdveTnS
rFQ0oniGNi5StEFJ1XxNXU/HNLNU1MaHd6YQC7DFyZY5B8UgBbXsghrZQGpKgrO9dTu4t9vN9gxD
t4Xp9Yt0L7TjedgNt6M8V4drAGnpCOQgbvNTJiMkgy2dNQisfK/IROEYQJfm5zy0WIYclsmh9jGf
5EDcULdQy0nzd1wd5ZF2urjDN8Pjy+B2qkJhtlkRJUvM3dH22im75p5pfBNWZj2uJwk8or6OcYxE
k7XgTzeKOvk2vFwBdWYFwvy7Pp8CFqeMcF/woGfnFreLwWfp+xbPWxxGz8fatQ7in6s8XdtZBw32
Py/IOUTML2dDt48fYJewuhi6vXpUH6uZ3nmJUc2JZnBFa5TTKNvn7f6B4ptB4Z3yACDefPKC3aCE
foJGl5Px65HCPtzMLprY5A3iExjfroTq9IKVIJFzg5d4ZRYg7v0X5GJRuI9IKpd2R7vCzPVHp5Hn
gOyXv2bCh/5pGfJXbSZiSpFi22Tcm2fP0CXHzO3vvRdvCQp9A+rMiNI8GY0sPaeEqqiayfsYKW8D
4nLpSwEUQfYb5aaRDkybIhPAHn2y2N394GdJ7S26YJ9yon+jHSMby83veTEM5lh+X1pg0y/IHUc6
tfav5woEhbs/r7IQg/+mgsg/N3RxUEMBsIBP+xSJEUYXumAkbWBo3qute6uUXqgIGq2kzamTgYLg
6kBEqFh35bBH8aNQRhrDMbel59bMEiS4uOSyKuQEq64KZIPUwdXtCM8bi8EynggK7QGcWzH8Qbrt
YiWnuBWKtwDxVMVll6YAZ8WsPIiqEtFVyEdyxIDdRHsKl0HteafJWguBYqHYh/txEKov4qGqzixN
rk2Hfqjp75vHNgO6nUt8qtYmakaNgS8t5V38zjXol9jmqiFnp6PDRq/r9JDhCPDpcJoeDoCDLvoM
uI6jcqUijdAzWypVW1BFafvANyFpD+/+1B7u2FZ8EYjFSt72uP63HhMA4R/zR0bfE9eE7K1vjhy/
0OrFQD29bS29qRHsPZoaL0FALhoqLENpZNnfJmrv3cXhcNr/lrub+LsBwroPmDJ7FGfNo9hJWTQ5
HU4K4kliK6QHiuOM7JltauUB/kjpZkzehK6SYIUuCEAINdNd59JaYy1exVG89b1XXUyxLXwzCGqo
iq3+1BPUhI4rx80FbphjUqDwhQo2VWF/QQPxezEA4hAYOy5+fUZGWndT0Di27j3B8uk0fDVBzbaK
P4DdeIzGjoPioqKKzIO4VDlGfEkJLwT69fqgXA//BfPeutVPxrWAUyF8tngERdDztCqbpENaMtG1
NMMs2US4y7fSLLComh9O6w/tzHJca2fHn9d/82I0ouHw8rGoxCYImELuPC6FvDAs4hHxE4pgXDkj
dd173NNjlKhqaIBMdxaJskApHlO7vlQV+Kjps4L56TlhjcTHAtAoA8puuxQJXWnBeraiZXTo6NLZ
hxO1PLLtK5BAhUhgIB7Mhz/ndnCgj9w8kGEa34EZapO9t/Smfx9KLyP6lmKlayHLFsIALFLwG+F7
JH6rizyNRyqOhjYIFwDq5d+TEpGqXuzEVELi7/kO5+Yj6OfVbqQ7EUKa5JVg1aNv0BheyFkY539N
Org16iPYKI0F3FgV2b5b7RuGNLnjzisKYDhmn9RQIvk7j0v2vy4FNR45hB5z8f8C/XVhE5ehaezj
2gmTdqhIE1CgUkm/r3AHMX0VHC6Z/8FDaZTSflMG7WX/4fnS0TmRB8kFREl/Ua6HZqwPypQpr0Aa
1MdJ/i8K2XUGG+a4hGAOXjiOTWkVcGM7LODyn5Yl9IrZ9Ltxn+xH0gjoBIYM4ELhSQ76awO9T9Ur
eq2vfgk44GfsYwb1p/G4Pl/0w5VGL3VpvL3fRZ7dn2kCJGXYYHl6XIuRbq6dpXz/R62FMvwi4VSc
taVx0Spyz9F/0PQp759R19i/gFoh/Ao07ehbUG1mqO2Zcm6VPFaopW9RIzQ4NtcAY0BKJyo0bBtc
gEYkFYPwEUFehgs9ZaVkuG9IPA/ycTvaSYafq4Zk6c3qAjhRathZQG8ksMhOQ257RZa2bVgbkacz
lsJTa4xP7h52ec2FIaqAV9hk95x9fQidtODry4wVzdl5fzcXJ894NwlrWjjSXAv2qZ9mkH3LeqZp
+qUuEnHPBvvrN5aSFEUv6Y+eOyzHvKESxaZbEnCLstDTohSN0CqF/kkLm9I/EbIaKTwCK/4bPz1f
R0yg3gARRqnm2gr98UIVRKWtVs41jv4Xx7ZCxR+Ad73iB0nhKlrwciuTa8V5mUieu4dEnU4SD8M3
YsowQTeygksQucD0AyyyWhwmGdyMXSBsqMampvgi3Fadu1m4q5TXtAAKRx9ikY3LAM82GrkaSFUp
IIO+A+QBogYHS5RhnAEMCve+7iwkP/zWPHEatyHctWj/W0PMPvjHYAD9DkQQxm8NM0HvB6jcpF03
nTQ86YlZLge2E68ryNFCrhc1cH6wVllSMvkrdSO5EymL9Py+W1VoX8DHWCFIhCCHnw3+9qn6m635
Ts9AatlYtJ8Ud6vJ288bNmi0oaxcsisvSdK1B+H1J2SAJ1KQoEQy2xJC7NVFT1MTyYXxysTP3x5c
6iBA7O//dMqQmjti79LlD5PGLBMwKmCpzr4ukVpAI/0vx4llYz3SSJ+vwofYtEoFV1hqAoOmm9dl
hAuKv/6qG2t5NjmmIiG3gb+pkUlZcKtIp9hcUoJbANwUhlrNuK0uZVlf5TWU6AF3JAW41pXB//e5
m/LX1VtHJiBBwhIAoiV0+Muk7mpsZY5mE0RVfcLPVcNZrFajc8SvQTfcR8us1vmKrNQI9aXe9+mv
0LbZrVPofgMsoPxu9hqbjPXRpD0wVSzHzfK6PjW9BdxbmSV2q52BytAYM3FygSFKq9a5d6fJme7l
ohhSELZLN3GyWbM3Wmn5nXLkcgQ9Z/J0L5//ELY6NP0Q9nFCm0YU58W+a+7+OtInoAKB8DwJ0XID
ab6ufg2q7rFhDmoXZumAO+xN49+3yUqHPjvnx3NCUYoThPPM73B6F6QCvUw6smPM0pinQ37x24G9
hMPlSR9WjPshsbmEi6wxIxMGZ2t+9O8LmrK0e8iYpf2kzmE4gkJEcU2KpdeLT6hswLiGpaoPeTU4
PzAW/IFybl9ogI/tjPy9N7c4RqdvdKXIDfuQIqh7leciWFCkTFNe30pAiw1evqLbybn3JtGcNVIP
g1FuLA/n8SFhF9Mq30stNcrJ9K3XcGdwnW0cz49VoIDNeN8cg3fL1g/EHCVCmvvIyfYRj8vobKLI
ouXov3KHoF0LkUHpleXiA+BQcUeZAw1NCbeGklZRVHq2TPPYOfBw7loi8W3oCqY2rM+OEaq4hk4v
mKlVnJeDIakkYD58abOr3Nlghr/xK8UKlar6DACzlvkiuOQMhlMBLIZ1hC5gCMrufD5Xf4e70VEj
5ndcj6U+jIvEupBY7/eCLcGRPgxGnz7uip4NfhxX2DWDycy3qf0zDdSNRXv+Q5LuaCcHSldbGeIS
uN5wyJ4iXIKGwKYvl+jxAqL9upy8yRUp0ENE1cp6PtyWRFNpZ2/qMUap0Pj47dShwNjPJmgTioVa
C7Z0JVD+3N8oQMpDTmAL5bDhHNmTgkPXFaRpFOifEXbjA0Mvbf+UR+pK8m9Gsf2B5dNlgTotKWGu
Cc/YVRMLik12c6KoP26MJPWYux4/ZQ+fHT5JFmkZPdQ2FNkSE0jAv+NMicOKZ7MqFDHp9rHxUYg8
g079td4dDGPUgxoep4D9rG71v/KOiRyLOaSnYGRGDXhItsmhWNxv2sTDIkkeXu52tqpj4JEd+R4o
ARibq+SiEr3qAg9uwGAWvEnrOJfer9kt/zAZGYGFhkcX6nDIHh7t29cQ1yZuwoUKzcxeQkKX0/Fh
s9NY+KiW7xWPV819Hs7kIaRhgg1GfNDC5AAgAiKFYK469LzmBj4xIL1M9eDGQZi5nNShMbj4BmDH
df7PlSTYja76yjNDCdbPtehoiCJ1VtOb1m5BYjKU7UC+i7UiJcXuKvwvKFpAXS1m4Z+6i0nneUlV
WiEXVEemEe41ioD4ky/48+lu+aDnc99hxJx8Sz21aqFj7Ej5KbjAo/FxoYzaMVdaDSLWWbd+qOBU
ocR9Od/WmOhsX7LZJDYms+cf+hRvv4JzgMgjqxHe5eBTIvl9t4kR9w2LpNMHAu7iOK0IJNK1r+8T
YcpRxRQr0APzdbgmqQia6hjhJS1C/Sp64Q+wnHdtLGY+akAEIpPMftp/LXUR6w8GOrjVCxUkIxat
4gSteW8Ra+K7+uttpUrcmjl/mh5GXCBLNhJvmR9dARYHJax6lyIH8bWSnbZ8iiuiyKjHUcGdNUz2
AOQscJ8KT4cmJbnXGk5OvY7sp2G0jGh1Gbi/N5cjbmYMhzeBz6ReKjivIprD+HSMcDBldiYHK/mf
uEhlxb24OjjjMLaDefmfqVrtq0UJRl/ojNzp3+/MLVnL41Pi8SzGHmal7Jx0WK3yKsTDGhKP1Hxw
e9yLVxRCRkwl8E7fgu7Pxe2c9zSvHs1utyUW1kM1oHKXEagH2sC5WCx4S2G0O+dHH2fMo2idpdhC
TafLNvJOg/RqUkU8o45slGtdrNle39jTQl6s3nmkvQwIdKtIo8x1a11OOW7KrPWWe1jo/q2Kahqd
mljdmvS5Pe0ms+CCzNpDdLfqWdebMOaYQj5F1l0CkLxMHVq/phc01vlhlTGPVE3Mv657hsYbfdxM
WHuB7Dovp7yZCGsF37vEL1AknC28PfUiuMGpgPY6kQ7Kc4xTn7sNKmKV6WHhnViGjDERjDvVu8fc
/WoOE0Lx2knwxVThNN3ZX+9fvDbog+W9B2/lgstAyl+LraYLdLI33va0N860R2KC2IjCb+WYs1wc
Sz3f7agBIWfGKKRxrRpFdn1LW6juryxZdAJEFnmRmnqY7EHM4InaZOBvsxW+yUwyaI+O7tuVJZsm
chBWmr6s8ZDNkE+AflJ965V6fMN152J7F+vdESIg98sCLyBbxPhb1auAEswt7nMmQdaaT0M/a4kP
V6BGaSybEp9IFqgmEkfqaGSkusMgIlxPhaOwKIMvf9D1ikIF2WvvWRwj5zf3pKOS0gc3IjQHZXCS
X9UpJq6FIIlbb0hwzP+r9MCBRmDwLb5W1C2Ma8PAZ/amWFXbMTUwstQsvQKT3C21iEk+nBLOKWbM
p/KBSuCgGxT6FOrC9THtkXH8fRYXs3HTCiASGH539hRBd3QGHjfWP1vQJq6t2/lazSM3qGCLdE4m
CzBfTeKM2LZmsQdUdWoWsdDt8135lsH7+kkAerkrXupYth/QYgjr6hfGQInHNl6RqcErU/o/bbVk
oR1bPHM+srFz+IH2R8GkkI2naMpt8T6d6jBbgcIdUArxEWN+f7po+cpdOuUbTy5k0+rAyxg17PfB
lBXFTxl62kdvnbTPxZ7EFNXSElxa3qJcUsEcxQYWjM6yxximJoMoqKcqKgms+0JzAuDAd1Ly58rU
R/HE8OEawXjCETpC3L0NGKxg3mQ2BM6LUoBeK63WgkjjlXUCCUOf2X7bFiIcB7fJS8X5TBsZaEK8
WZDURD8de7HAAhNA/csm/d+Y1rDZqnsCMn2WahRiroFDvGuI/Kyw6xAr0FZT9GHdMx1kjHxAPYUj
rm3nagaRwqD9uDGWxHFo3wwbDeu8ajMndmwvG6RE+AaAT9DSU/FnX2eGnFv7eCrTgrShkOKzj+3G
zLS1Fa279ane5GeJdIALz+jbnfpMjrZRTdoZRAAQPyXqE3GIwd53fCbF0nvZciEu0EdyRin2F+/X
1OHGiZzJhMQOK6Nsw4304e5BzzZrI60H7vrXHNJRu4rjtFp4SVTXdi4KfT1VSKPeO/Lg6+S+T0uy
0hn6tUai6rFqg70AKCp6CCcuRSvpNx1tYvQFIgBbr38owO4nPujkpZVb/6rwQUJirRel0I5Ucurr
jn5uQH8ZaYkz2HpO/AAIzQiaoxsbDGT/5CHinx/rUZxSgCi74VeygRYkDZpSm6SpvPfxbrvnGuJF
2iZmfeiVrXt++U4HwyG8+6xQl5Db5+s0fUnh+ttxL7Xvm3KdOgivDha5X3KXCQOs6dr8LCDoCQhR
pgusi2DR6KjuloeqoAiVj6G498dKiGkMSpwBxi3i5ZiP6hiJgc/jmKJ3o4ciImrGI92GgyylUrMh
sZvkWn3OXjhaR3apa29q12DMk668H/qhLuEzvvImAajA6KQg00lzoNQn8P/Bn5TgLKRT0PwLayxE
LQOPraJX2zUG1MNG2q131rSmHe4M3NAmWDwS3gEbPcriSa2rZPLBcTeACtSQ75NjA9WL9kxxO/Mm
t5Smbdnw3JYmi9LCUYdZiSTHvEH3TeqA1sFa83RQd7wP+1ySURDRvUKN2kmMHH+sVQbemGMSmiSt
xaF3tZznmjxOB9RkUXGtOz65tPS1Y+ZvNyQzC1C2ezt2l+h4sh0OV0CgkNedw0f1u1Np5To5EUoz
eOXvV8x4LlAsVBb1KmVd7jPZgwMtw/5LgD/MC+J7vZ45c1Lj9Q2VOUWCS97P5OzwtHhFSU5tFZH9
XtM5GzNz0KyZSyME91iTG7wqKGYAWjrakqo1FvB6V7rSX9SAQ6VOfpAc0NWlPxVQIAwL9Vzwm/Co
/0afQf6PsIZDnhRsnmo+7RLROkQ7PuaeQ2iSTypxvy2x4vYIditR6ccN0+upYnbYfxADaDTqIpC1
rkWoy8D5HQkQZ7iKRjnlSazlIZuompH8gKdXIpwLAFbGTKFt6XjLjB3MHoFnctglSMuzLf6vYBLV
4orMJC2Ky0NnCLrS/BJZHbacM5gNglEpgIhEloZRSHUTLWvODYZCFcKFlyhtVaUU8I+e+qn1CJYL
AoVWaMVyjnwBvx2y6LasFsu+sA0f4FlhY9Bo7ZWYmDQY1repTDIB4YpUObRweuFrpvUFLjaZB2/N
9u+Vuzc4BRYsfXlFD4zg9DJeKbwQliLZlk59W1DP9w29wxRV3UxYzf60eRqYQdZBxn7/R8ArQqY2
klQDvucnMSkgFBHagKOsdPsBNIrVPJTslKEvItOsUgw4l7rakPlaTbLZwLrpvHvSGoJ8X8Y5Ji31
HSOTFld5lHIX0Hc8vXbaJnkwgp9ukGpFxZ39zZRFSkVX5FdMicgliBcvkGZ1IX8uxgGxS12YtICE
UuvKQiAD6A5LvQ3Yjok9QJrX39Kt+edEQFnT22BSqGXFPAhCx40NiOAIaGoSzrgRnyxAQVf+55Ut
aP2uUTUrmwnaAIAxJqTr2+0B9QSXgc/Avd4iSDhpDrwao/KQMAtTkX9t6yqklq6LRnmmPx5oBSsX
Jq4sRWAcj0wXolMTSpnSFBq2ZJm4lAC+49IFhZxpuOxc+/68DEanejEEO5fTbgVWw3tcPaFqmHMY
bcpELC65vU43txUDuvu1mPRtTIUfaXui30Uj9aLm0lAH5RnXPfQnAtHag4Aqkov8Cg5S0MYyhB2m
Sod9DmKd3qdpD36tJeUuc2RJ6wWxQfZpdEj8C2n9KtxiZ+6uGxfxaq2EZl36E0AnTJgU49ooNoA0
LfMhqNT53j2Fm4j2cAaVsPubIQhgKA7inPMRR2xrBVt9QLIhuiORdiLHkFuQfH09qRAh590PXsLC
UbDQ7RVdXnlUKyPssuZhtbgIw5/myEp4ykdi7q/UZvPhb8gHPNHp6TyGD1zRXRT2zRnXkAwqFvhk
4JpKVUE0rWpP9eduonTsI5zX/Bng3ugSU45SAC1J4iZ8L6Y0Mvw/mRUvqC7/pQqRgO9vrD084ADp
+Cd1mWw7pyltZLdMhLLdrao6NpLqeTRv7srCL0SNypIFt1K9EEhyOZYKvPlM2M7wjfwJ+I4Vdss3
taduO71U96BarouUfC8IrTXkQU+VwEZ2ZkRMSBQS/JFfydRBJ6nyd5izgASZY/DA+qRwHNVynuYL
bfgG3vfTXkjx9fmCdYTCXh7yttZl0Zo95fYOnOBWggJV1wntgBt4YClLq1N0j3A6o7Ds9kC73DDw
/AuzEWBAUoHtraSESlgXd6k/di5oeG9NfdZpxfjHwh9uwK6hHxGNeB5WYdXDq4VypJDEC+Xw65Lm
MHTCJZi2Wa7tkV29ql5mofuHy8tBIcopo6PGy5mSYlxV7LPf8XyabOH1nrv8HT2tbGqrAriXIu90
3Hd7xLeOrJ4vCcwx9LZPHqzXQtMh5DJairKuMfBOeGUoy0iU/2XU21E0NnYFQC17V5SPIcPe3EgI
uP6zY4SU+uQylz0mxCVVsYfymSX1eIB3igs2GO2UNYT1NlMKCHqoM7JzyX4d+tHQdbRIfCKHGJX3
bLBLixzQZ1eNqnqTiie1POS9TtSxU/Ku7gvMuX5ECXcyUSwWzdIJZY/2S5AGpzoTLrQiZd4yxwzW
lbDwskm5S7TuCeG3/ZxDVu0uHsjUzUuL9LBB3UsUlCWU7rZDf5nO4H2edceC3UDP78GpQroD7+zC
r2kKWE3F4NQ3bzo32TO00baQBAnONJnUgxSAgvHeaUZJ8pcqH/Lg5tV+uILI/gPqSxnMU9OTEuHf
j5awh+WoIrFaTfmHQtW6MeRxm7BesysxawYjbWjz92GIcmIYjzM4wX9gXRUqUBPFcrxGQlxWYcX2
sI9tu7T7laEPS0kwBY0vLGEr8a3MYS/tAUEodtCiXk802l3+FG42vPKH58JbQB/gEwqt7z+CxEzI
OujOt+4hAr1MT5P4t7yr6VdKYA7pwkLmTMxeJdxCLkGG/aG0qKxExFNfYgLBWCdo0VNX9yyZqiqA
8LGM6LbAbp+cBjeRkPnJETaiC3cvl+slGcCDiGZf/QQhRB3+VneSXWYA5XDtfo3l+9F2uq9ClERa
mHkOxB/o4D1W+KMABxXNjz7GbNtavAFeeE5r61IkgFYHu2iYwf7N7XaddDY/aeVfOr//DzMcpbCm
THN4xJAzj7zi8lyJTlTnZrCUPSFR160hRcCpwclVCDIq2rQVw/f+KclMJvEimWdi3YC2+rEO2ElA
fuN3iY/LKW2r0q/T0iXGRF/iRNFPY6KdNsGEwQPuErcMnfLnOGK7r6uSMlCC/cRGSQ2G+hpfhtnR
hmMmNubzAgDeIjvZkJw49XJrGNj/c7ldcn9lTewJndRNG+vSKe/5SssQS3juL49VOjdSWSwqMo1Z
8QOmG4jjryHWUech3ZSZOHe8tpwWgb2KOFuuwzUcGXwa3XMbGILjAgG+obOS3IbFVIpeSRQdY4lN
g99+3CXHx00VoEfXK3V4eiiDPW5p63p73VImXFYnGflVYFnobPg9QR2y4lnlo2wFjQvCStfyZ+sY
5Fqa7G59rXMeLr0uKqzjVpUJVNEmG7RWJ9+2r34G3Ns7R4IWa4FRolTysiSgq1neY2z4nFbzMNZn
MNuhHKxoQZWTjAd9M/7AL4dRH6gs+9rTAHMXcdXoNGCORzH2Q+WaQEZuDSYDp9VXOTi3lI4MIsin
Z+HSaDi2FXP/MFWN5vMio3H5tD82SG4SIkAo6oI9F3+Ymz68ZsEniXdbW/1vgsBTDUHUZ37j0vXS
tndYzLohU1FDzxK/XR501xvQpm6pGLff1z1Bvs6VG0RZHw6SIrQGYviqNZWRYAIJ1Pq775iohoz5
46mvbWGxQWgVySwYEI6P3ukSnMLv/LoWhd0cI5o42bUKLVnMQMK+2MdJmlHsNScBrzlqLt3sTldV
IQP+p5fud9IsHMiAImpMQ5U4VCOarcM6pHal9LLkWi6nYya5FX100t0DqgdKrse/8UOjodTbR+XG
j8dfqIpYT8WfFrErXtwwKkob2xtBlVYqVGmu54P2BecIYKhrd+Ltdrr3GZFPVNcWRg3apMAkoswA
Jqudpp38+7qM7TGQJ+FTu9lmgntR5/8VjlOwQMDFlHkV22F19vKKpJemdI9QZU55kPxMnJ5F30n4
fhC6eXo8lzRGsCMRk73zSDRBU6CG6Uu8E4fi8Faew+lW1yMmIaNhiGpEV2TCleOAWZsJaWC8wfSE
8Be2R+AFzwC/N9vXzbcHyu1748T1odFPJyr48K6T7AyGElNfSMhJ4OeEakKS4BIDZiRliGR/xFIM
w1JpjIYK61k8hpJXeZmIbspgQG/O+o9TI2TEC7NM3md7XO3ilnE9ieuGg9qRkFUhcKvNbCoYwaRr
GLlGjonWmB69zEq2N2Kffk6agQg83Nr2eRK8zF7DVgBpEY85CzBKfeVFCG97LNRh8ueMMMH64jfY
OCZGq7QAxctVBLkpW3Du9/3HNgfcDtw7WeXqc3mT7ZvVgUM1VxmLPYOdj1UKzRnPoMf/SqWi8fay
wobGExDGCW8u4LjOY+hY1EV61SKZuoD/zLCSppY+6x5gHN3VnBiA/AHllusJdpEjMmxQMzfp+6yB
2uOULez61t2SQlTKqs4rxKXmN1/86NOARTcLzIfHB42ubGwyzA1kW81V/Mqh1npkJ2YzEn8afd7E
k/w7RiKXH8NRfm1F5QmL3x5r+TS40xOZeyW+7J7u2LU89Lk0OBoZ1uopVG8/N4BAlKMgToAneNgD
lxH6QPQIfAmS7W/rpVREgqapVvL6fLKNZR1mFzk0GNpziYoX+ANs0kKRf3/za9brbU0VdOkacC2v
wAY3AV8TjqXb/U8ydyRCHDIsozbHGcoz3a5Gd7CEuyumZ1FuH9iMoIb313P+HtPGI+cklArfM5Rk
Vzpzc/fax4+h3vwy9P5XOO08s7oQoQlZZmLnCcTEAH28N1MLLN/p4nOBzIHQJBdkv77w3m9Rh8ED
w2Y3abROg+ev6lCuULoUYAch4grTd5y5jds4OPuZF2vJHt/rnnwETymVE+qnTp/nKeYfpcjpcrYh
mTeCM6oHdieTTD6PII7z6ea/24uWOg2Zl+dVRP9KnK20GrasVNdT9W9VXq45fqwCOE4TL82RTDCd
1/vEzCHOVqCCt/DiLM6ZkSW1Z3DryPvu+H5icufu5Mlgxjo8kUZYcQD3CX4dhFca4j/M1DprjZn6
oLOG0a9ia74c7mXsqijj7ldceXu0/GcwvxK/brM3NrG+AovHMf/5g/NniJFh9WjE3D6b4HK5V3jn
a91Klpeorl4Vz/WYxZiuo+p1gsIwGdiGS1YJl2ewLvD/ynA/Q5XM5DnjejuGAtW9uQs0yxByvgZf
FKHDL13qcpal9rWFMuqMX3O8IaYCBBl4qX5vUY1MeyWr/MGcMBL/aCxIe22ZKXZcYINjnXQ5JckP
4OLikQhabjkKgudxnyk9HWSF6R4Tv/pa7/LLy30R8+We+YXyKMgbQeCTOnDv/3MYY8uS4hl/V4sr
nfdli+7lPejfX2FRmBBuqWbV9dWl6jVI/SCGTsNY98iRa+IPxOJ3BZ1wq2xUEpjC9SuV64hXKj5h
QYBVQjP2cakwSlVBbfPMe1SQFxVJVHLZaz3/mpZ545Rt4SWczKs62tREakb177ZbsT18n1kAXJ5M
8KK2R1aCuZnwoXcTunHjyrJhbcO98mvHyus6aP7zx/JHViZqgVbF0GtHGfm5A41Vj9zuPpVyN42d
ua1Eb1OXUP/4fE58jnMR0iB3BFgxPPIjfDWTu+M/psIYhgh3AMF4VZFoEWRkcqqMej5pT0vxOxQS
srPd6h6b9nJxm4yY3a+zi1juzdXzmHdqEvoYmyf5a4HLGOeT1KCRxcDXrsUusVu+FUuZupacLPN2
X08QWcIg1VFkPz06PbUcLPYi0zVp3JtZIhdbMBWc/yYoif8C5gJOvSBKVyUMPNLPSYodQwR2BNil
vYoFZTXpsJVQ5o5XLJOtzgBgwTqx3vxf68dl99tnfRXkFgF+sdVf8HDiotrdq11CPZdfyILx1K3N
/YTXr2jopmta7jp3wLkRRgQwemQUPpts7lk+N+0JbdCNhu+mHIIIVe0i7CFd8jxacu6dg3hj+TCp
15+knR1a/ohwCag+YdHjAbJq7pQWhlUU1SRwHADBvPd3Ky9nmfCUbpWswG1amZVX7Oe0A71znen1
RrhqJBEblZ5fHC5HVv5rLplhcLExCfbP4nnsyCbNQKywy5rxbPigXKEYwwTkTrajHVVj4J3K3pdp
IcWy2UtF060mgn3nUP+pW15/CIjX8WfMOrChywuGJrY3kNU0ACBLelEXc7Ton0joNXyEvR0JJVTO
5KaRMxen7fw70+66cWnILh9ydp+6Hq2JhbVI1ZuznlFl4JdpH3z2kG31jsQYZI3wkAmU6Usuy7IV
B+BjIIxztAd/ldybScIDkhX593g3O9mCFz4iQ1dlHIo9A5op4WHzAvDgQ/IqFbbb/ZoUFzlqGQvh
wPgNGajVUwRuvvbub4HrRrW1/Rp4ZD7WBx+r//VeNRKktM3p6eAcl0pcyQ3nhuDlpWO8CcG9zIxy
m0MwD75uM3m3SDH7nId/ycoAe86byg4NrsrewJFhQk9WAn6CmyPSJDMFV1NxGu6FFSBqUs/N1+5z
0JZ50RaXxCzWa7xrJZJAjLuKyQcJdiuPJbA9OmeTXV+3GPz6tghDQBTnzel/dob8+ZFSQy+lRQcI
o5yZTwT87U4O3TVn6vS3lCnI1fhoWkj9NEghj9mP0S3+oWhh0TKk8dBaFKfhSjgxiOFCo452gIVN
3cyL23QkGCH37tPA6pbr2iPMtMxJWwM1ehVEeD960zqj5QblFtKEqAL6WZWryhBBUSbJ2MX6gftH
kvf0AkyuRRDjMbmOxqnDmwbbw976kuLU7HYF+c3RFyZz8lMU2u86QYZzkGr9DgxiiJbQ0CkzzfWb
duocrrTxB02ymwPlkjGdsEI1reqUWTYsM9lNA6akq2UJULxiaV4QsLR0z3Y+Zi1Q6njewOwAuWf6
lnmOy7KHmCXWkqKZr2KmuGK7OXQK/rTOgKSXB83kZ0v9X6J0fpv670GyT7ptMcHKQIy0UCGPABQr
IDKrt3pu6I/F8EGJg8KEl9AfWgNz+4jvHF0DVgM36S5nMhQBkBDijWk7Yf5sIMIuHksykAt2YuQR
GgpJ6K2joWwDxEojG8Akz8Ch4vNGiXKkKRfN8helO7gd2hudBNjAdW1oSbNxis0nblUqX8RTzS0L
CFyfe3NyEcXr5iBdgun05JPvb8tgQawe2ypM6kytsAe1T/92kpiaTj+SPL/R5163U74f18cnU4df
ceSD9KmfYrVepQvfR2e2YFlUfvUp9YShGKI7Ua+g9ta6XXeXvz/DmQ2b4eBmPYO+9MBwguL5B7R0
PVdweAPyQaRFmJXteoU1PtDnYVL7ZSTdYqOn4+VIw729q52/aJZVNrTiv9xsVXHMdWNipNVqeoQt
QabUKAFLY92jqDnpfWhQ+A+4tPpTn9+q/Vck9iXQw2G7TFm4dXkMUsZJNLUiCLaAsAdyKZ+9ejwy
Dm4yFHxFQqMJn60oBFSi33fYElI8+UiqzUknacf0Ak76D2Hq3WgYQoVe4YPQB2BUsD6jNY2riCuD
mvCHhYzRgQl1UYkFlmTIBIZtqG5qTmG2+9j6xHjkLjVQuGyihqAH7BPTnh0SZdwXEFlSrM/6PlJt
8PsJ1dVOzOzIusVcK6bLUZt9+UTLS9B9I8jVhIihGs5RRgVwVlVFg9cZSbNJSE/6HJIXQgE9v2Zs
dXJWLpbXy/3rt+l1sLyDaZqdDiPn7UiQ3VIxJsiZ6cEnpzGAQX2cUnQgSLO5XIWAEa8pSdJmGJkn
u4EbrJnrz7y+lSsSu17sXC3k2d55u+H32Z1F7RXxdiR0p2TvRbvdBap5499/cDVu8c/xK/t93SQE
kjqL+OVBJk/pKt1TzOaupUkWohboEpZs3ntX7UI9ulu8kN2JJJSH/eTQuha54Z/gvdfTE+TIHT36
7DSuTnkXO8IEf0RWZwXDXiuVbuKAyMcP20imHbxFm73hqv77udCmyNJBHa4TS70DOBwBUvf5rwJJ
KoWCeWaxvFn3ThHfOTHUSgTDbIH+XwGuQgS/m6s/KvgoMI73K9bvF6yAVoLHLPBXHapNt/6IgHnY
0psczXMcApf7pKW4dHJIjDm/omdUkb/QS8KMPtuGoMELfVGBHUQblEK3rHeSbLQW6iHV6DIeGcnl
bGviTyibxT5GHLbg+pZqNj70IpSpTfnI/HeEDlMKpkQfP5cDf+EqhYoWcfXfzTNFuqf6MP4WFHCt
MQxQbILn7tBcN8J1DSqsuFL/QwoWIRAHSJuuUubLPE+Y8jWqR3Q91gLGR8fYkkx0NEE6LepgtMtr
yIJynoavQtwli+3+D/14cfP6rkA0P1p6HoGshBrkyXqgKltrY6IQosCjaUqGwoQCLJuqsNxsN6gb
Td7arptBTh9ZNDbgeAT3TtqcSUeiUIj+o2pfUAkr5x3gqJ+roXCRvaXG2tIqqnzsbTrzO9dHYEW9
YDKxeDH97X8KboMqaK5vkwp3tTvRHNhReo9E4gfrmuj9NK0OzEp+rIrbD5tQZ2htVizVvwOS+1A3
EQfXA4EgmTSGoSzK/4RUgRhX7biW4C5byj/tGtgZRWVmVVn+obtOxPXinGGHKHmU62NFnJmAjyih
YB+XD08/5X1DQuZIyfj+QNVyZOKZLpF2d47OxaGXJn55uya6FNSN6fG6Yn12X7BRiMMK+jrpQPi6
4YMlBGoQKYZT4OEwQHJuBXX2VQc8sWB/IauWYh/PBwMzDObtWKsMO+DO3MPIwhu5/pMyvXjr4cFy
kpFZmr42YQVZF+FRr90qXuD03chz3gn2lxN21adHsdOZDCcw96yMdJNkqCh1CYShoxu1P/0S2tvA
XIxpcWxAz7P5V6n7Y03QOnHdzxtwXBRHboGxws/oRwP77eUb+BVvrhUrG5wNiLD0BQI2HxhEj+lV
daWOlkpAbQCviboszdpHP6gus+ZbksRR/lyASfi95KiCxJQsDuHbeIasGbsc6HYzmvlg3OYJq4RZ
gyfkwjVuyIGM3J2JWKbCBGNTS59EgfT9EsgXkcPb99XloRsT0GhEkFDX4OTZSR64VaQVfOULU3Jo
9RjgCO7n1LDBKEQhQMxEqp0CG7Gyg/Ukv3OIOipwm391VornLN+rdh3Ada01aMi0BS0IN4L3zfPF
mGEzZr332WlZJpSya1e9vo8wrmZg5L7kcBuxzkrsN8R92FEk7oYzQRm0uYiLhRZK6RgS0UFPVvT0
7JCZlMiGBXLK5BMd3ENWmBY5JBmOHYgr0PrAza60CQ33CfZnKKZwihAs6eoJNBuOPJ7gYzSJUVTR
/xrkLphzdVCpoS7BbGHl4IXcpdYTHJZU4YSukISOzYDWL9BbHMdPfm3Y0X/9rQ/NBSxscCnTOLGD
ugvIWAD/e7BefMZ9q0BXQhAI1m2ENrwbqRNc8wZPqM6Ujwad0FxSsn2sh9dfjliGcLlzBrXauS2Z
NqoZq4D2YRILS2ChkJ83SXwyq/r1km0de3HxjQRO6ONR7n214ykIfpSSuJPQnlcnHQJuMVFkc++n
5Ofcc/iDVXdS3M5NG8+9x0IChVh2jf7Dpk5tTLF+nOpQi9T48ualCpJ0JA7xQsbPYGuQmy0SXGHC
y/C3xPCJvgySt+jX64zjFunryctlbUuYcLnYikZXJ8KAR5DcCgH3ThSK6gYV09swPTvIwwVj/LJm
lgVkGkO0mTXUbpwqEqziw57OhVt9bibbBp9FP4RlfYlN7DjJAg+7eTx/faExM/O0vHFhpPLzwbZb
7H9Szgs3n5VwNtgR54lI12IRBUFnK7vSAfl/mcM1qrIrhtL1aQQvtj+hw3u2V6IVs5vEvW+pDBuB
Px0Du62VzzbzWTB8wtf1P/VjWWo92VKvzK5tdXv0BS0nz4iF4XR47qAXvM4RPre53vSMZKus39ev
X5Ncu/ilaKVixYNtRVS8WIwiBXH4HQS40Qu/dlfByvyoK2jDYrm2HnLTMr7NdgZbye9xkEBZcWqS
4WmLpqzKtpC9EnJLBJo3Ge+z2ZJPeUgFUXNnLK5Vao4huQM75xTxttSbW1WttFrdEoST4Pt1Jouh
hoW8A50vEwHTxSMPBwQlyVCCOIT6Y33QhCx05cANlkB85VD2mU4mgZnM29mAZ0B20EflVawV2DqB
yAMkfuiFrWUPj5gauvisWwgqnxJSgQ40DQCrtoHeAK0Ke5SHYr2qPYIVPkFSjM+I0ABEovBzRniC
jQjyYaDWKPcnla8yD+/ib8pRa9mnatjlpdBbaPkCAgnH1L0VjDE+fu8wBf7DuZigOcIujkaRDf3h
gRgaCkVIbXJYMDU6M32a2KPXuWYH+Utc84UXAhzgtXUQs2B04vJ4wpdxhiONh/uwJpQWILWMzDaE
blOFud7av/0ug+aWbKb6J2vlDcgpVmb/bS9VYv4wi62V0zKqekhkzwuk8adEMz6KBNC16nKKOwx6
D+hcyfrsrplWfzamS44OSkwa8ynNnuLKlHAm+jIUx+Yzza06aGm1Dv2UCa57os5uiZUoQRu5cMtv
53c92zluBvDS+H+oz7Lhi3aWP6PHafQncjnjcLkc+qZbeXkUXel/4CFEaP8HMHOjX6fYnv07dd6c
i+4WAjHmf88IpQJ9GBZ+BkQSiXjdtFfiIj8Qjj9FnvCZL435rze1k3mBUghSJ9/cT6gCg3ZZXmRR
OR9L+fD4feXrKWUTPCcDsJBmLOSaHpL/zgjdLTnBkLhC4eHK/nJiO3hQHiaQzgMx99F3dSCD7wkm
y1MKNmABzdw+CN/B+oNGIZghXCfunGARnxbFJAeZ/N0iieF9JVQ/uIXokrbD0tiLLCn5XhVyCgS1
vtyCU/NUy5HD99vkDWtSTsbaXBcX37KU5EXwVY56bPAlkB5mXOaqIkZw6/S5jwrGAEocrhC/5p4D
VkeSBrPBAy9lz9sHvP0lvo/f1mdkSvdmnTY0JsuqQrEfXf0wYqsd5T3XfOUevLXyAT2YipDlQC0Z
NY6kR/FKVnbCIbRuevt6e2W8ndn17ttBNzPawORu41TiRVOUXRMNYuVbifj/pv4/GuU6MT7qo1hx
5d+7FNmMjViZiIGhWEVoaRdaYMbmla9VoQs1omFtnT1yppbGZeA59maBospzmktwzp0m8+0DFenq
InoZXCcktR+YdlUOCE8oi/s5A7fqD4CuV2tI8H9+/DTil+Mnw74IIaM1S9etHbEm+jo13ANdm4rY
QyaGu3IvQrfTGMr17s8N692h+dcoTW1h1GzGaGbwF6WGvzAXLH6QRdPHJPzJmLZCCM6jOw/iEhXB
WYXBr+uQoXN68cs4a8z40FIA70E5NbnxtUIQ91DMDkDcc6Kop9qDI52ajXmbMoH7Mgx0b6NtprGE
cQP1CHM/oJA9U9GnibmO2fFN9yRHtQ7VNzyIYkXtUS2eKrH+8E1TXJ9VdDf1UNzBaDgzY2yVqmX2
JKslrCCN/cP3ox+WDDSMVhGWhvL4AKYk1UfdgnUQP4xP5oYg12bkfxltDpfKfzaATZcUuYNwXjCi
IZUMuqpqICIMVnr0ssd5MSDTZqzgTYS9MlQSDfjr9cB0dbfZXIDiMlcoENPk/GuLuJFbBxbzSwae
6z9fPaoDxTqE2QIk3GD2uk3z724ogt0p7FShHB5eaQtd/5SK2MDZP38hiAqW6ipaInJ3T+h5SiMd
ejDc9TgumMpzekrv+/97oAyIQhgfUBtdfrUf+TMjy8CBk4q1Rv6bJrcQAhBWbi/kJ8FEhtf6XeDD
8r92c4/WM1XLyyuhhRs2A15h8gdRZRSvfYkp6ZhqgcO+e78q7vZRHkC/VFaHap56xl4FgMv124Qk
rOOUT5uPYf+0wQ7pW3f5Pr3Vshe5fmYePguTIz+bknPtdLEZQBg8W8i8zokQarrC049Wxr7zwoVI
hFlMhLh5slKtOCcAsYgZ7TGV5rWXC0tyCQA6cfO3yz6Z6sxn947xMPNTVPvex614+gZWkTDu6lNq
afOuqjTo5qA1gE8+uOlnSQtn5iIsRcDiq1WttGbJvPW8qCiGe0Oe88az1AeU2j7NjZrsvGirzPGh
xVvCUxfmk+hgxvNZfoeHdsfSqxesIoKTzs2guuu+XZvGbViwicCvlfxE0KErREOBZmMZy5DOT2PQ
6QLb4JTJQTLS9Efi+3ph8JJP/gmilyPrwE1rTQAw0kqP4cGsD3155qDp6qMzdl2l2+oBLUNfLfnI
nNKXvb8aIbc/dh5hdOWozN8BR0Syvlg1cUz35wA5a9/s6pournzNmFOHRZqjljEkQex11m8FcthM
uDHpCJ8hArl2gfA9ROdyBmouqnIQzjycoxLV0RGIUXHYrJcMN+Ws3R73BikegdouOCiK3zjEEUpC
sE7WtItO+TZfAaHJSUtuZi9jhM/l9FXJ2GRBajvBhKDgoF38qnClb0pCnddWUcD6DX2Gch0rHhmX
eEWvyU5Z5rtpkw0Svyy822JKwel3Smk02SSq4ZHtZSVYvxu00GQ5S1mLXdcvaSRQEgbt+ZhqPF7S
/RJrjgVF+56YP86oUjEkN97pHRpBXhVhkAlWvtpR6TwwCOLZ+ybh1oAx2xgpq4Hijd43InOIROWW
QUhp3ll944A7/iEPbT9IJkTx5lz+IX9toewZAGYUOq/NSr6YigC5c5DPsypjDbxHYpWHpKiz74wx
7QymsbhaTWgp220V4go22BUE2xOoSMbhoFyTUVo2Bdbui0LsOUS91zEXRFzbzLk8U+FNukZT+QsO
m3FAy3F+eOpZXcbAMU6z/xrp2nF9hRoSjxwioAeO7nhheemFzvzP+1fQ2sbVfHJMTfrIy6F5avE4
uUFl3iBv/AXRWIXWKZIPKzIDbuaCCgGP1V1CZ2tDqdQRUBOi+MOoRxgRvKC63o2G9c8ZsgKOWl+o
XSw2KBCYXjziENiDpeBIHjR/h1S1eL53OGNxJXoEThp8wht9E6CWp9dhA+hy/WQnUqAeQ/ymBHXF
utM+qxSKTIntRtHgREHfOpI83b7Yfu3jt3rWsa+hJ5xSxybda99K4I4YJFCpBR7xILFQmOTxJTEv
HiyGOy7WLpxCYJ+4lpybykctsNrIB8277ZfOwRk3r95QmWi6enKfWIiPaCpDkt+SjYlsiAgdauju
wYtP71z9lw6kolzTbG+MPSCTNAJZ2+nNv0JH7edfvAn3k8+imoujKb0fWtCJeaB4dLvcULfRJvUl
g6Y5xAg+z0chgpJeebb2rz6QJ58RjplTvIzP+cXpAHos4vUMjkgGa3KAmr+by/iwrQZ0HHkbAiSK
4YS/64z1qBiTd4BYiAP279inOwTnW9RlwNBANbzTL0gmishJEHvvzi/xR4cFeGaJ9gv9ng6pl/mj
SO9kpXtP2XpWlN3oyfiSb9brxvNei4jXv0Fphr1CEJkWU1ug4pItVhGB8f6KtchuLiez8NlldIox
fUw5nymG+Mq2Z1l+E3+1jrbPZTaBwgCqjlK0lC/02Dy360Y6CLs6eYtBm16Bq1GhnbQbWwDNrNYC
LcZ2TBa63De8zx26Cd+tXgLvyg+ZhGIL6Exb9GSBgrodeW93dWwBURQRhp9R4KybwOVdrmW4q/Oo
b+LjC8D9v2UChFkz2LMLDvA5c1ocRHr+VpmfbkXIcFwUBiuEmrOQmuX1jqnG611Tx+7LzocL0u7B
BUhEivTtbf4b6Y7hxPn+83fNGAssrgPc9a2tofagmEj22Jne5+hrhqf94ZDfEXftmkHxWZEN5szM
sE3daDmcxKyyYi1d6t2DZPoy5U2zGmMurZOSdj83UsopYIZ3cjWiO6eZ/WpUySkEVPctz+FsAERy
CJKXBK3imdamE7vKm+Lugil4MjodjgqnkbkKea+eF0GINV6G8xmDQs/1QT7hc+qvSGkSu6cg2MNK
GDrvnZf6ulLchr4oYP77wu6QUmgo8VzPpIrudvskqUEfeBZ4ah8yWEmmbZsfWOZnjb3B9Ql8cb1J
K+doBReh9SA8TZv5StHzQktfoMbBS4ifGRaBor0r7do6xW5Oau36cRxAWXOV+w8xS7TSX0moouWs
6wfQzFQJgfeiCq0EU77OW4Z+oODKAEYyjUBDkcyjtY9XkHUz21lEN2cAOpvQ+/qCjDVl4lTwG7RH
1jYSLqkjoMQAF1Nk08rVqMTEJPYkWn3m0ErqFG/nHPuPZI33YX3vqrwjk8ezOOBrOe8lell+43P5
lEr1CZ7ZwlU/7xMpL0INZDTFm/O4v91A49imHXcPUziqCpj8azJ/+E0tWXRxbgRWb7iLg5Waa767
St/vnlWmhXpUk7e7u20TCtk+OB32lmXRfa02GBfPYFBuRMhUTQ8aBPYdeFxAH/qdgeP6hrPSN2PU
EZn1JOl1T83CoBfJbtHDlQ1f0b0Ulr2aB6H2EXBlxBpuczT1yGZY/7vn4SBIErWrrKaAZZhO9UWp
JM4alhggir0E7MPy5BWXvy1eDfA12K+4o1L/mHcPz4V3opnRAsIoLTyfComdw9MO4l8ChWv57qv1
3/yirOs+Fe1se7sTg759k5JW3y4Sthvp8pk4WhvSbt31SLyHghhhBln0fmevu7qnLnB+6W+k0Z9A
FpBQ6s/M0tJUEfq5x9JWt2bFWT4rxkSqsmyRJlBN5Iy1EU6JCPTmZHYx3t7XPj4MylBGhlgmhzBG
OdKTQxV6yziCjDksuGvL4i6m+6Jx+cKHzplemDWsl4Sy3WYEyfpNAFoowSEuEtN17zGFFD715Emq
x/HckViSEys8zqajHPbI7Y0vNWzvJyIbE3Ah22aCAcIL9W+CB6u0ldHbiygIEhC1L3sjHyhMfAP4
Krmym7pGldEFVVNMDbFU/zWjad8f55U7LbtwVoYMWqhSIWqKHG2SUWQhEetlr9AhcJN5k6GZkRp4
OP+kS7i5YVipbMoV5xmAJwnT++6uoNVejzD1/CZSAf0JG7Ly/9WJEggYn2TdYVrycZCbzmmQ4jVn
Rp5CkNAmZ9WcpSKPpuec08AC450XSpK15YdBiDW9QGzYbY8mY1/yBSg4UtaK8wOErXBpzRiUXRQv
Bzrb2vSLKTDoJmLazg+5Dy5bK2jJ+2Z2MjAU42DKLkCGqpBxqVPWCAh2XoB1+aMDe9WVNOAVbEDi
GnfwqrVlS4zWXm8vyYc2aYTbpO96d8xtU1IuHtZ3MyQWWEvBDTwBlrODTgZLAEzlcLMZ6MEdvDBN
SuYlA9H5jaJi27cQS1XN+/4NR4lNsjYaUrsCZPIJ+aVNt/t3ALuEJJ2e2vvuefxLzsEVZUUP56ZV
a8w5b66Uc7rZsowIbdhEx+jxoKSxjzJGrXiO5FQN3eAGvD/VfRCdcSGXSeNlpYrzdj2s/+C1kxBw
OaAikhdxg7k6xHmTZ4vfYM/9LTyWSVRK4uufSb/H+LmRzHhxqqHw3Df1DacvEwxhwig2J2C4g1FE
Z+qBuLw+sYDAVzECcRyRBRwbsp3W+nxYF+xvvsS0co2D8icCDwGy8GS1T05rHmmUZz4Fc/aJpAxC
nt6J3CNDiEV0wbjFCJWtiLK+Q5UVPAAGeeu+gYaoOf0T1eYEmcnfGiRAEfWg9vnwriRuLZFRiFy/
LUGIJS1O36clK+0f+mUUhFw8ki83jelDJrsANAhpwa2yE7gLMfCi/pKdfvGgSwzQvKksmbq5e7Q5
+mo3SIsE0Ad+jBqFx1XWcnqi0PQ2GJ472hvLoadJ4C8sop50LCDY6H0DOEEaaLXQ/ksik0YRkQrd
y3M+EbJLPvpsJR4cRc89gk1+gHGzcRTWLIkV4byTGmHZEnP07lJLn6gvnHsq6IDmVt3VCcx5mwOo
YnATRCxKW/l+b++E+7COUqPi6M4z9ALwcIEd1TK8DniR2V67/qQ8AKa7776c/65yMPo/OaO7WZBY
uIxf6lHXvDrtHMt3J96yu/DmXiW3GlHFZEyigzyx9uo4cRVUPdcP5Na7CMTdpO8kmzr6itd0PHb1
xE+BFVrTjTxfEiGMnR4w1dwHueA9+uumlDAlfxysM26TlKGTNdjx5wquuoWxIFOZwlWQBOYnKy9n
PAjPFliaSjULzRypisl0hmVhhto/r0dsTbUupeyxXZ3RtF4WJR65H/U+r8GoDwk/5sPczM8CHZqb
4C0UeAWOjgUf4cgHSucoJiqz9TVbCfS7tuPnsJZryQjeuYTggsIDgat6LqBUkbv6ToONZGTRmG/4
WGN+sao/Tc1wyj4SFydsnsUicLvuyVohZmdtQuPMypGdeKJdrwUdGRLgYKDcsa5ed2YNGE7YrKnb
NJxXbYgt3rcL80PQgQmKC6SPLk9UgFCVuB7moXFiQsYHgkwszwByA+SQqAAmCUS5RH3PQ0CxHQi+
azvrfj2bNs67fi8SsXiR4uINfz2KT7aiaiITWU1Xd6B5CP/HCM70rFKDb0VypgVgVzS6jVsMAvjE
tEHmXnvi6n9rMNzIXo1BF1PhikPVV/pb3cASjTGeFy72InX3bwjKQ4MIoNgHtBYjfy9yHmJUFcZa
adWAHHGEZEmQKS8BlbqYyNd3g3nbExVrwJ3IPTr3NrVDOT8Ws78cXbWtlWd2W8fw41Tp65LXOQER
yf7q4YsRsvYFEtgJkVHSVYiPSZnKmUCbIL5Da0vvnpeh0VW/DuvsGzuWcfcdSADjUPjoa4Zm8xrx
nCaXvpspSglQ28X+S3jGPNYPI8ErBf5BDGx0L7TF3lyjEp+n85W9ibAjGVySlCzwCyBZLHxFFZBa
G4YwFCXy3qasAefrSD7r5sB6XtzZQzutBV9vEH1EIvcy5Iz468r+hKpQps98mxsHlahl0iN51Qd3
sNb7JN9qrq7CX6qJBmQ9cg91tos9zXbj3DLs2FN4377alWruH8wXsDYjPNeLMwMK6I/pgv0dutU3
QRNfNdU9PpYPln94rukze8IhuziJvMeTtgIzt8LBanxtChqEBP3XJQtaKKie3lu5NTTORxC3pU8Z
qgPSBRNPRx+pDZRwoACOB9+vKNijfxjRBPrbiWa/0N2Sn7C5uHYl5Gd9NS1lMWPZSMU4kGcmptzr
svKUjbqFPFF7hFwUe6h29kxx3Jn8K6+HczJMmkRtHl1rdI8TNVP1aPu0zBx95iJ6h3lxieEOknIn
Ze1lINsexXx5cpD9XGa+YLDwfHHZTx6X2eYqoCYNO78xy0NAgZ2TMb/coC6HDL40aE+gaBZsNv/6
kw/ZpfEdVrxAt+L5ENL0e4wsj6nA9tP99cKkKh3gYlx2g+YQ1natqT46ZsU1G6S3ivdZ9AvHGeQA
rPwqXETBn8UBT6dhJKewu71KINas4bSAl3xFyhnc43Xja0DvsDKBm+oo+LaUuZzWL98CecX4njve
u6kY3jqxd9dV/92F7MzyOtjFR5VOA0+ag3Ro5rlhQ1O9hOCkjV4ZThI+WkZhKq09eJSQdr2X1xqs
CgfG0p8rN3VqJY5g5IIXd4b0lpm0IrsrdTxfXcBbHMzjVAk9pdWAhokg1rsGXitZkDx3CDAExWDa
jKW3S10hAB64I09zymEdQeYfWZXItnGCWjiivdKTaTUkpMNF6Ljql9ftlyreM170EUlC8Vb3bsN4
DiM0Yac+PORqXy0qs+QLz3vIM53LG1vV4SGxSQVPI9uHwrCPkQXl4IpYEhbC8tC0rwfwwezaYW2Q
bvtpP0zvZNaGSR+0/AvZZA+W7k5mH9fyD7BFITv00N7hr/3IA+k/OrK3KDCtXAMQa12ewID4lig5
NunVVWCM41u9D/O/ekdfXo1AfsnPY/rDtcaH9zPw9QvyJ++oe+xfGen+rdzzf+tnnX6MqnO2at2+
viwxn2d/hsBBYiWQW5EuRunSyq5avSv+GVaZqESMwVO0GDNCsCkBqcoc52gDcV7hwsAJKh/pEL8F
ee2MZJYsx9LGEi9s2aXflevovPA94dNfKZFxcED25on+PxtPoez0/l9nYgQztV+FJ+rRbWKp0U5S
vZ59zg9QqBu7MLKiVDk+CBBikfK62nRaHNNlUnKYO7wt4lkrX2J6ACWFqV5y4TlTiNCY9r7ZMeam
RiYUUVrSLzlW86FxMTK/H+Ot3OJzeQnUx9SsuxICjgNNQuoHPjdjDGUUZSh5cObUrkqMR5m09SIx
HgeyxUe3g+VJtJe0g3lBfQVeoiAl4zialHp40+UoWcFVvMSFRuY3qgLj97BM2Da+MGHdOoz19TWV
OAVbHUj31cEyJUCeeOqNHavbfOPuyjEWVH/oV1a5hsfRevVPaps4m7v6nui1Sz496YOMG2plY46F
Y3+ONJQt9AN2e1knokT70owasxn3T18QeT3/n6QKXSsz1B735npAQdxaSKMqxnVeOhyHME8S1BDR
pXVYPBjH2ajji97WKgKmw2q5DUmBqTMGWcebzkedi6V53x+iNG9F/8oucuF1Acn21TXwZFmfmVG2
WEdEuVSsjrZXHdfo8wR3FfoPLKG/5t3baYgAwstmp/Ym70wqgywDWy+fyZqp2h5+QucukWQd1Azy
CcB7GodZKBplCVDc+7Lfe+tasmh61jqNNQ+EgEtrLi91F8E+F8VC6ikutczGM3D1GaoDiH52gzRc
l/ci2aVAQJ7VZQ4OZLunb4m9+Rf3/WHKA+/+uLAj/xRGe27gC9puH6C3A0p/a12f3vMMDKc2ZqiN
Kk4SGE47vBPg8+a3yKnDgaF1NAu8VNZN95XRbsV9JCZ5OGCl3qn0pQRxrxJ/z37vRxHZZQMld+fK
0yxSElxiMMCznMy/h9k2j7kCOOvjo0NUCl7C8HHb1qIj+lzqiZT7LwM+tKwdF8v9zYYKTGfTVLff
nXP8dighax//1eduwDGgk9uaKQu6v8v8NZ2X7W2mRNZNMABoEZW1QFT2Ymo33fpYiCxfDV+PjMzY
aHAVkwe+iaS2ywCJUwa6SzSOR5MKX/rnIisww+7zAhYFUn9KSirpTzxkSBw3HpAEcUjY38uGG+hE
rXahUoN9YCNElLzznQyNJF4MyzyF5mSqfd4GOuHyg3Iva4IdPwBwugtPQFfjutO+CVkgEFtedD4W
3gmYCCxcl8PRYVGrsdWGrIRqTdoJXQX4JV/SN/6qKSzId0gHzi8GPkP0tCsGNJ5N8Gk9X8AIkjvW
ROUg9apmv3t3Zs5X3xWdoUSKUbQSILB6E1F8Bd1s/lXdUCBPud8EX1Fg911sIXfyejvNFuG4xJNS
kP/R3wup9L7YTpSXSftb5Btz86vg+Q5pa1K6lBIk2UPFfAolTn4neVn+JiSMUEc58hrcnh3N6Fbg
LkKNyeDAu9Nz5cpsNyxCTFvHx2J+tqvfLJqpe+xbVb3y4F9dJ00MwICCyziEWV2fAxiMF7S+TU82
psa9VkCRRQ3WBBvoVLjc4Di+YCjxAflXV5HvwwZa5eCUqsbC7YyLhQAjZRQIKk6Rmp8/vABYnM+k
+IZNx8dvffchfbqQdlV1UNJvqRaPg5NYB47aGlLGXoJoha35dMYPmxHcuKXt0BRab4yUmkRsXpg1
ulWfSOhKwKxqbd/QrYIW4Uk7syp80aqoXXG6qIj7QjDqdBHOWShADmTdin8ZW3ZIrbUIN0aC8tZm
0r4jdiWRa/nifm1ZIQGUh1RLc0MR8aM2y9n10fIhmg7vbV7bcJSjxwnoTnYJjKwUkJJx9wSSaJrY
OqCCO2sMQ2iSEKsAXPO5YlDmlyuuv5SIjJytASF1J/PY+Z/49SotLylDe+kWrI9f2CHGfQkrMi2N
6Jy0uzX+r2hCQ1j/A8GV1gqpxjiH1QOAjzSBcxEyoCqlJlwLiYhDJe2f9an5TUxVAjjhxetxiSDA
AQjVDG27DBXTtYuPKcs7fNr4VGYfCHQxyzf56zcarbkGb7wLBuEF/fDkDYvmbAor7GXcKo2eRZQZ
Sh7WQRik9d++v3mk06UK9fVjLJaL/h8ZqlMw7JOSVChhC4B65WFkgZ7ajICdFWDCxfv3/IliIyYm
EpNDXrIlwXlBtR3b+NRVLgHP3qrDmNw4m4V/qABK0Ysa4jy8pTS3q3dDFWJkf8DbBn1YS8Qzm7JO
jCXx5dU/YuKJUyaczyrjkmkFVemMo+VdmpaTwS1tHLL3ma3cZ7G+k/D+c75BjesQpHptutFEjWNV
jGQnlJK1YNk51EObNgM6h23/vw46gHw4wueRx9LSgZSgjq9Wvy3pjDi+2X294fg5ITB85zax0xOo
K757WmSoTv0QHVeMulaTncYSnjrpxuVbElNp/q8//adocHJMKM4Dl9cCrdB3lhzQEwjkPfrZ9y2X
ZO4DZ7WuL+zdBxuAwaRaASP7VCFrAqw4vItnwaL+RGv0nPSgAsz3wn2Uw7RE7lUsFGXIWrqS4ktY
HCOAJK5USyD1DjP7Ci6YOUm1fyL7rJv+AXaORDnDgzn8xwmixguE6ZA+KNdhNoVWHAmDO+63qNF9
NJinV69rBs9ITiHNSpdV+Ffdibg+3YqadlK/dWVjCxnTXVVupfvv0HBxISGGoNCVXN3Lwhqn32EG
qEOLVSo80gIYRdIpI2boff4AgOdtWhhAyr0+Vt1XlaIliZq3mFdVmEHXhlG/aYvZbpv2JUIp6imJ
4F2uzxE9ol7oBvzpSjnx9ONXGedlV9EQInvc2gCx67N8KnxhV/tyhPQHAPNcVzJH1wcOtF+Rgusd
LhU3MZppzoHW9XUzFlzHTpSklSeQWS4Om131jllZk9XHSZaYHFqhuOAexLB0WENbVo/+XbR02E3P
C/luQE+YqkgbFzDDBsTdWKWGBH3+PZ3gu8h306Cvf+i88Ukw9tOAZb5x6H5aLFoySme3B6ExBoew
uTksnje2XFHFrgZYYxMZwXawu4sy0rMV1yD1nHVffD/Y3pOL5Pu0mBf2CPOG4vmu7Xbr6wgYXIob
+sgVctqHm53vEaopS5ZnsamPmZZCtgTRubGg6CPM0qkezuhzlTCIMbtMmQf8maTK8LUHwjvEJ+4B
O5Wqi5HWE4SVhTPSLoDAU5IKxajzXi9783fVakdmu8ruYlsasFhFJ2ct5DngFafwKFNxlNg4BMQP
G4AQTf3PSyDJcuBiNMxQV5SMVU0ynNKABlygHZDHbtHRD3ZlULCCifdcvsvREov4GUFgLT4oYB/K
OYD3S02WtffLqsbLKf3pBkJeeguN59DCPGVM8l8mabPlaxnWw4P+9GPrrBouMng4QfGu5ZBaeFuW
FOuzQTxoqdXL8yGQbG/TmgWXuH7f3EhZXKpyZt/1YWUNi0t3Q0+F1KTSkNYYMapmltjXLikdUVqd
6Js4QiSri7p8Mf7hJ1prHxhOcAhxlAz2UwRAl2aJwABX0ERmMih2wG+QES1HJYSoY+3EaB+PWbrk
XYKxhGv9HQeKZHy62wa/ZrQlHXoBP26sI3VCrstHIA0iF5RsbWVlzr+ikdh8AQ38OQx+bnQv0c3a
kKh1PMl85M0yGOU3JrogmdGMyuEP1HOzpW+xjSK1IrwLJuIJeVWrft3F6qsuE4rDWjKOJmcGbF2T
xQLGtlzw3jfYN4SFZn9wht9pvbqDacbmJRuPq6cvN6dOqJu/jSZZ+EjeNbALEJz+leYDs8Qwtzu2
TlmnaxbQCyfbwy+fEilWvCfOoZvhnBrtHn2QhR8a9K6xiIcn0os4lU2lz8ETs4Md74DTauRDzVVs
6k72SPQ5XQdMWtcozw6oIiyrdN1VPi+LM3qJdEnMSwyMA/3B0dSEpQVao6GeNqul7cGV3/B5vRRH
KzJyA985+b9C+BSCv1ZXQIZ0VuoEfticNiFDuC9IB+hR+Z+LJPPwp+5nk5J2O9DTqRyyKdzAF3un
OgPfyzoEEQL15qGWqv079bMB0XFBYeHf/Qk0M4qGxb2F547ImZa6qB7czHskqkGZou92HpmIRG0X
chcsqtWWzqQzgtvdlG/apsl56SuX/clyN/hOZvgYcc/c/qOYRlA5Y3Iu14wlXMCCLK1Dfd/uMwje
xbsJl2GHaPq5Zu4Cf5IP+RYYusAG/JbZ29oMXhAuc5c2RcYgyebO3EV992jqSEjB21o4FwT6slRj
ahlG8D8/qOrF1st+TTKvHcahoys3+R0ocNtfK5iHWB/8Ifzz7VQvYuNvzPvdhy/zwD7RlqdpLBwF
PuD5Tjdrm4PY59213PE5fMHWEzZSSFj7StPMu/aMhPgW+CJKCYu9oOvlWEm8c2X0l0/sP8yTzlTV
lL6UfDlVbz4momf3XLCwspvi78ROvtodAtaT36TUGsNhf+3AR0nOEBywu3cZttiyNX6zutpNB+D0
G4arNy4oRjCFW/XWPrhIgqcrfwk/O135X13O0QsgqpINru0Dwo/EGGk8od4NgOzTD9RiTOxopSuX
VJCL1rqr3OfOFl/xpiNj00q4Agu47J+W7F43fWPYGuPZam45SkGsC4OZkPFasVbAB/KesbuFNASS
5vOvgKDXuhndX75/h68awiyLeBb1RJ2PGBWdpQUrShP8ckxnIVtuIYZyldRiIhJVZpMyfvlnpfkv
7+tZ5Qw0bCqLagnrEXTWclDFx7TGsCk+I6UJyNFxwjbS2LrpGF1aVyaZbFi+Ls0T51T8wB+NGMmt
M+l0kdzrazWn/R8DP9Nd4ZQUJt1R+bxjXi+o9rekf+3Wqgw7k68cYKkiO+VXN4queJShw/OG8UtB
MUY7WwKNxdNOwoS+Ol24L3cE2Zma9a3IwCQwBpOf2gu54g1z14Sms78F607ywQe50Do3EY1JP3mY
KBPnn/5QhV4RxReHoLcD5WU2m1y5FYwuXoqcQyxefJ8WgY7bSt0NYGxGswSFgMlAtHiYQbvTKIZG
yInVZA1TNwZfXRCd8VsvBzk6PLnLIRLr+pWHgYsjIcsmITSZCTHqayugJXmgXSOfEsQct5SeLre7
IrFy9NfM6jJDCvhemmjnlg5Fx24UeidDjEEdpskDPhtKy+VqEjM236AcvJFodS1F3qDDIEoqet6a
4JMDH7m3E3w4S27HSj5/ss21KDn2fjZfQFC9ggMLb/fVgqePwGRxa4S+SWi/C/3tVuIuhsS2mofP
r4N3fvMJLqdNv45g4/iOWEEvSm25nEBySYDzKNPtaxiNM3nnOn6fChtV9JO/ZbWlQL+VBBJS+1/W
sH85U4LTDpAQy77wZtCukbQRMTpMZPvl5xj9lmaQd6CrY3YYxvNZk0/N2BIwyoLmW1Q+9dFRMjAu
xO4JyIHx9E4fN3yYxM87+mhzHdG8uxS4h8jj8JI593d34fIybxckkhObONmt6iThlmtJV6GTtliY
s3yO7q+yTu29kU1nf38q/AyqXITzOKBzQaqTx2E2OxIUUlidNRAlo602RDgHbGfkXkneL65krznB
1eCZowAouhr8l+kd6PdmAxB/5XtQLewuaRejLJcKeYCQ3PEOK/AWY4gXnvUah2YzHPP3MH3Dbay6
bpYKP8MHd64cO2Wkzn/xGYsFWDvQmRO2u4ZKp4YPb+x8ZPr2dSPfPlo8WXbcVlSgExeJj9f+7zr4
/etSysgTo1qjx7h4AZsRhv0iRNdoFdsGFRsUQ6sCon8RJWi0/cv6jpQDh9IKgIC7bj5kMlYdGZKl
vRscCZz7Gg4Bnj2I9R9j3Gpu6Kn9PpxyAWIBcKqbUE0UsZ01+nFNFPDSekSNfmtv3uzgCqCw0HEt
u3BlR7W8ifS7ALakcu/EtoQw3URWZ0bnN8RBVQpRMc6jJXwdyLNJMPJbAju9tmFMQjBR3OKgelvy
vAQdcKTUpaN8yCFe0VS082lhhq7RmT6ZhHx9b9AiN7imQB1TFfBtv1CFND9fTIU/Vjqhys351aD0
Cqoy+jFAiswXFhuNGTyfWXJzj154L3XFw2YyZkdXz8fjms+84DR/ObZ4/f0lvI20mfz4TXPHbSxs
0USOFizw1L5WonaKYzD+m+jcgDFV9KdDjdbtYDxospcpGkHOrfsrNxqm8jmwr/D+c9GfpVdIOVjX
gunNPfpQIslTISrbg+bTXQvpAeGcL5UyuCFIqTqNQXoCGDXQhatB2ECvDs59nCSRGAxX9Grnot2j
JRufYYE+gJQfejgGicoTMKcriMjzYsXCfEwXSdh0NP0IcC0DK9rHIZ9dzmU3hhWCi56swZF8j+BY
+DoL77QZvwiT2DnkuVJ0KiqYxGHyjZztFLTFgno0d2yhC0ND4s+qhfIWeWwohD+VDS+Uhdb/B8e2
VVCJ+9jyhCHYaB4a+wzifgVH+amUo2AnMa7GqXrThO2vLQNQQbYAtgl3AwWxkfbS+G6kdljT7j9f
j3sh5cFUZHjti7ztJgFU9WkSFFDiSWiNEngtEyc9Xf+rS0rxXDFQHdI+BzEmkJoqBeEWV9OROaCK
ZmqZqqRNy7yWFHoSyqeqwYlF9/UsE/jgkOOrE0Jx2NRXr9LWRBGJilrd72K1Nl8qayZ5LV27YuIK
Ms0q0LdY+eaGZ9cN1dZNSWEuPD8hGokjz3TV3FtOErV+pVF20BucX8V4Dc735kn7aavaIB9mOT/J
uGyxj4vBbzVFKhx3sSiug4n6DiX8WqfLaWuE1FsmdRn4qUYTNu7FMDis+hBE7ZD5ZlNuQ+gQ/ITv
R0MvjjOlQXPUlYPAw6FPdvV3Fl0TdzlEZQYrQoNMd3e1WOH7JRMXJSzjYMD30SJP2j/9rWAUIakR
M/RuEKxuWAfo67xYFXfH3b97TI+nLheSPi3Sf6NU2fyKczSvZ5ktwE2M7bFrjEvkAz+2z0qx6PQC
vLMYlNCJM4uxfhtFzRiwxNhUBXSlkVYexD1Oe0vrv5Dp1q/wXIp2Mc3GjlUers0oXgRNG56IJ6aZ
cW216cOuWkob8F1QmgxO2rYuPhbVtvnuSaXh82TYG6mQ1bHkMoIJLal3itpJqk/gaQU+8TQevd0q
3I4bnVo/50Dwtd9AeF41kyS/g7R2GCba/GLtZr6DgsB1FcrVi9q/lHCmZuuv+oQqSk605qW4a14V
xZoVND1opXMOeEBaUohw+USmEyhvJ04RBgLjBi9PahuUZrxpz1z2se/cnsv1VbMmP43o90yyW6V2
ZfBP/sf5xN+5nFThZrfaG+MP45A4P7xtKkMT4wXZ9FPkqWitOiaVMOWx9zYbbrISGQ3SYUsMIZ2V
VScEnJIloWvEfxA0tt+6ZA1qsTtieGb1S7S2gDelr/pnjB60upbUbC/2TdGTu8ZRaz4hIwe4ckJK
8NHfrsvJHr/4Wi82469v3hOabfxGxVtIeR6SN8smPoDKg6qamTIouR8TWw9/uj/TgBEFeVK/YfGk
1+G/8f2OzUJH4vzEC3ull+JK1gP+fQf2mjB9ja8wozjW5nYpJ1s/21bnnVEKkSEzmF+dh1Nx5rmB
r6pKwQsCDpIUAv5SMZGYxwkjOxkA5OXA0IHl6kBLkxp3BjCgbiW98wHv6Q0EYg2pIXFyQ7KyIlZX
9PNY7yH24v4+gNH6YKvAHDJdf4EVrtOuq3tGS0cWRMybsvBba2QvDbB9Wv9K/6fG8eD+bZBxL9AH
dXu4Rd88vE0dabbLzX7pMIRcueFQPAaCrATtG/WOPXbLrLA/V8zrLGGXMY9EAkF4yavAFizKpaak
IMqby/uSEUX6jwpUHcjaWQvtJnDWKiPxAQ9H/HHcDRQdwQyjfhUGITFm6CPm7WdwePXo2+Q3htEz
5UukUSJlQtojO6YUnHIKBcFVCByg5zdefe292heTSh8O7lFLxvOHR0IulXGJzIQXMmc9CRtbrxSQ
MlqUaJB/5NynJJmw6r1IFdfxAwCdlt+suxIWZ5xxkXGXbKJvNReB0juBthg2Q5IHG33BxcT3xflg
nXFqGXpbzmXgtPiFDhr3n1pRtthn97c/dXmhaf5gjfgDQmsjH5KPgYWhSMNwY9XO8Q8VPQ2nMCic
37cTi97R+Y7mdmgOq5/tlJJPx8NC2c9G2K+ncfIy4YdczPfG/miuUjOU03MHAfV3BG8l0pInFY4h
RZmaK4R3/OqkCEngTRvyvv+h/Q2DJAWhxyPc5AcJX8nj7yhYCt3xVpRsQv7dbMVJ7oKuy3q64KgP
pzfLaxQPDO9s2V/nyZnfowL2UdOnwjZKUywZilKnEgKgH1EiqhZwqMHjE3tlWuDrNOwPtiEmxwkE
ViZGDYbSQN6S1pR1La1hss71u5EZHkDrJxbI+6xNCkX6RC6L4k5HxX6mqPRQaUmpWbwHT8NjMRk/
3eEAup7zlp6iuwSTRyJ7noYLrfCD91+ok5MC8TPC7mNlTuAaxKhsFiNy7f6/Lop5EjpcSE4UYFyA
/c/a8dhipX8IwxWj5LvM+Bx6bTS/mWQCOgjUmsLWPezkBnGDLVW4sQJdEh7UwRINiB0R/4nTopqc
xRQtglX2d8+zXOZWG/DjsA13SEwxMrIbbb2ebEehHZlcJ/BQvXRGNlSOsP7a0o6rS73pJ86VboQD
tGXAg/o2GWM6ZOS/udi371bVaM+IGlmW2r5ZLs2c11IQ5w5KYWuMgdEXhkBgq1wX6tAyURF5Og9U
n4wsy2SgrE0MTjLQPr8wQYHn5f3s2Rm/82hZbyOJLp1afZE9enm8wEWoPDBQ+77/pGfp7xIHIEjA
xKX7z7/oCH8oQZV5DUarUNzXvBpbT1KMlGUoPTqjKLhErSgr4TE5XLG+CafcYbxofbLN0RESb9Xk
6s24du2ELsNxGEwYBVeSgz5Ps4LDvGs5rz4g9f4ZkKBHxiLGS2dvux/ZVfRgx3WcHTj4Gl16wFOI
gq+e4hHyS0pGu8s5vrmF/hV20uyFn5U9cP2xfJYX1zC3/uRpDij3D60emzwIv/EpIvlACdDFAadg
oZzqT1CvpBwt2ZLj2r/xneUQKGbpSzfj3bmsk3hdBWR+YKDm+jjVI+W9614Sft52KG/MWqQbiFQ+
MR0ljx9l/VHkZNEUBq31BhkwnTBf+KpuOUxRu8Rp9MayZlBGyplRwVua/w2qz4vOCGSHdUL2kHdO
CpTiSMuEhLffVWA4nN3vYRy2rnxhH8IV2GqONtSWeZjVUa/rpWqw8Xd1yJhtXmr5WXDbLsB+R6QQ
Mm7bJPkRuA2ZTnAR5qB2Z9zDOS21PmEEo0Ye/Z5Ijy4/BoC4yAUamAad547OtQMhkdYB+V4csJ13
mbYwl1dLJnEb3xq6FR8H1/P0woUvsg6er/IcYsPD2NHsiNOd4QBQBWqtgMKChBDA47TGFw5geZG1
v3sO76TQyxoX9lkEocIrGSWzhpwUUMBS08dbzpkepy/gKWc0Fq0XGW2B9c0tTlu83YlN5R3UIEsU
aKz2w5JY/2w9Eizwg6hk6VQuottBppJLBwZRhO1VRYpLEs9/aj+7/y4VOyr1ofgEi3Vft5VArnHk
o5OaHEXFp/oHCQeei0v8+RLi5ac1iU/pMlrJKVbzu9q4HI2J6CH+ThgePogE0PoMYDtohm+IEtv/
qHM2MtP8GaAwCB2yZGo5AGBnauQOBKeoH5WQISeslcBQFbv+DYpurmDLSFocdzmejE+f119lYrqn
ayno6XSFFMI/3GZaDFG+b0mZHoOIkx2d7brOv33bu15nPpJbkAVUmAlzQRAUWUOC/zbIIgIh6Yww
57E0mIz3AtjQtU+5xSiI8KAP2ZaNcXfP7xqeYMAoWlhHDSADchCOa/NlSzqF8ekWJoaIHLWfO6Cq
Wlu4nZhlHBX5uxuhc31kKAbavMzOrVLoa71cyO2Dm5AtQd7enQMcU7yW5+ZQ36X5NxGPQf4+uPMt
pNfnyf3mSXfQdXgGVch9Lm8ez9VUmZ4Qrx9yPeFfVaB38Q6VWDlcrs2SPmjBbI1eNM9qSFS8jcik
IyOHJSZvYHgNZsL3jyNk5f9I+eNNL5s/SD9dbu4SoF9ol9Op81V03u/+dUDg2MHeknG6+7MMZnrY
UaTzElVAuJPTH02vrhWglfUs9wkY6ckA7wFzr3LlA6iwGGLV/Y2oPSNNKbhNWWUxc/GBGUzIDdRy
niWr6Bnh+tNhVVrfKTRsNKgEVyC5o3qkXrybDiXTWnzxGobU+IK85Y3Z+vZTtIHNMCeA5g31a+Jk
0kwaZwwQQOe4hGfQXpOr/vkqEzoG01EcQdVPoUoSxbtZet4lASl6Cha7xBWjUvibH79fIfC3ZFxd
oFRoCYCJHT0rx9DUAL2X/ChRjHHzGpSAS0PZblIwQMJUskfX3RcnEaN6lkTS9IuD86nx4c0SAk1q
x1tVtxtpSVfDBWAO8AR6VIa304KPZ9DQ/ileVkE/nEko9/bzx+IUF4KiyCY68WAp5KrFzbhcAboz
45nKjYFMYXFdFtjbJleIMOgxTSpKmD4ou08wpnOFUkOeglqsTlduVKA5hn2ZZTIyMD6zs6XNGNu1
h99jotN5nx5w518N7/lRtY2JY+89U8/t9XZ9kg9/3WWtgjqZaJNv4arVpxXGvlAq+nyOwD8BfSlP
s4XgZFWvsWJ0ALGoEmMiAZOw2anh/QxVMpy70c470fd3F+9y7z6EU4vijJhj1bDUB5G26a7kmckH
ICRxtdMDHcaPr6ZXa4ScTfXl+IDn6bZ+EwjTmV29UuPkqRnSwzaQ77OeuPI2o4u3dVJ4dXFuTfXM
lD7zxA+X3Hn7p/7Jhvc6Sojw0b+PxZ5cZ8t7UalRg8T/KQCJ7K6VzCnOo8Q8oxv+CCNNvTKO7PYR
icONI1eK06x8tFpnjmTguxW3aQD3sdT0VDBTs2BvEpi/7Ih/3ubo8ycuI5wqQraWQO5OTmWh+rqe
h6fXiju1Gcfg4xFmECjMsY/vMP1hZmns6RYiOPzOIix6NLvi3TTrMc3GGPzk641uGbYapgCZA0yX
CDmCzbOzmmBA1x/vamCSBnbCd3buUXi49wttjVBpJ8R5WJPy4txm8pf0H1RDCV4f4zvuBB3rvMJA
RB+dBI5G9ONeilP+jc1v78fsbq/eX/Q4CjS5M6aVO1SGoxUdZkFW+huW9Kaj5nqTtKF56oPDTF0o
b3MybOuo3YIWqHvln63X6rxKo/CinKXoqbNSBMMFqLeaocoNxF1rhU0JRTYAy2HdZqa/fVzYuMIL
Ox2xd6hh/yRlmC6v7sppuWIho4jZKmoju0bF20cEqJLolYZhSCs2cw5X9XGvLtKZYx4P38HVautW
kpfIjS3AK1oSqUS67zuBkfPWUGSk869NARPzcKL9dgLx8r6YPqBinJr2OCOy23usZAhKGpUbDySW
nxspPBowEjuavTUtZSa3RP9GzL5tXecdWMx9L8PpWgMjQitqD77lQrYI7RuOvX+8c5a3LXcR0Dj/
CRvfTmSkGpI06R9rVKzUnq+JvPJ9hBEaAI8JO2VnLQwZkeU7ZzrSiFGQQ62YOYVEv03eBAtCm/WP
SJRE43Hdb+bFjyuuOXwTzZy8pDhvkQeWtHkVVpqEZbUj6Se9FFsIjAf1QcCeXiZmA3GD7Yce9MtL
tDOIAsHnvfJj/AmSV+UjdyeA68662ZKTpZJPDJC2+ROdZh/t5RLyGyjjIXS6/hLqyNcmsa/kFGgn
ROueBxQey+fBXUMO5TOE730Nq5pBvbudv8BpBYmnMkHb2k7rrTIYe/vuepwmhJL+TJwdGwlrlc1F
yLHvDU6q5MqPtOjAMNotMwMfGyLc4r4h2QB4G1jYJMbPN0rOAEszzEa4u/2qLy1j67UQtkg0ikyF
RJKU03wpRvmUMUnIvBVVeUA3Q4DymxIMqepjc2tWs+9B/uloTxiWgvUvKzldPrDvdYdB/5UYg5WK
tqa9JLypDbe/lTWDJM8B2QEAsmVRnvhFbpS0KULbfyOYvvTm2iimU7L84M0GRmcVw/im0TliUkLH
mKtNKSuf1wuqLIkmlnJu9WEl5znqI85xDxzAocJJYGPzRYINUKNWwYi3KdjznqfVMsJaSPXiGJsK
qtmW1gpRZtgrNnzpV9FOBZeWXZQGAjwkHdtO1QREBhnFkiSw1oGmffmPRg39RISu8SartvWyxkMa
3CDRgRdl00DyFU/DOjmlX6Er5F2PFMJ/6BBMkgJP0ygxcs7ioob4gsnBhF8BlbTQw/UnZ9dVfLaQ
y5SC8UK6A2ZtvGOe7halksTL/xrXDkCwROloJ3vTA+l+MKMl9VbaENTQBijTIgSVf+LdGo6xzomQ
pIk3ZqUv/n8dKaKV963nrhyyEsO0QriUVuXo/LmKmfXLwvstBU9UNZ+lOO6YkpSy5wHTsv7CjImd
xTnd4T+LDoulUcUg2fcSET0gW7Val4LKmo+Dpqfo8TLGz0UcyN+hD28Bmh14BBnAS12OiubAjkm8
f3rNxmmdmihaEpQB3/8G9avp/yDEC27okA3f8+piXonuwwMxJMdnuxWEpik/n8o6Y1mPOyfZS2Hb
lO8UmJ/b3FCbrDynAVoLtugl2iOT4o0BrwIQ2YDMx3dxaMSDML1htY028o6IN6dTGa2ND1w9hSow
Xuvv9eDDhEpuwzfd5BbznP6cdZMfwaew/5EMAtNk7CiPcsLAMkTw83pVKMGM5XY1OP6BGlsd71Bb
0YtwF8/u+Nf/eIqdbsWp1akggEXc+RBQlNil4mp9fMYQs4f3iNt7gmUqgmfZxZyFuJGbvTGakkmZ
gS21UcX7paxiWHZDXRoF8VRXDHgYawSZeaSr0m4lPbFqsF5jXYEo/R0V0zwcBW7hZLuEpE8olMHt
MqXretcRHxxmwBrS6O0L03DtaTEW10syyiDWZ5/PCyCAkktqTNFgCLV73PpmjPAn9UNbCqe9j5BJ
bQxjsRZZR6Vv0StxN2aXT2juuZ3bwCKQErd85TW3BHdWZHGTwfnjQcCmDesg1z0yHju28IDkVvL9
JVm2+u/FKZcqKttk0rdL1py+IPf8m0Y34l0aw4IDqGfCb6v+Amq8VbVUO0vyYxD5CoJ9w0IwwmC0
EP4rDC1Y/oGf01FzGYcOmBfVRRw2T2c+iu/nMajbGAyFqajY2YBAlKmN7frPIgMv5ub5aQN/8w2L
NmucxfKLN9CPNol6hntwjHclMNs9X9rYmMSTQgDCHr5J7oFV3etTcSCFl4N8T6iztHfIgl9120Zb
2BayFPTPhgaJ3Udy1ySuEt56xxXFB6lVDwXGjNEmmmqUnxGQysuEIGDjPkuvg/TGYMx6wfULWqrH
QXxgX6zN9FLzdpP+3K5srpBhcrTV8rnvWCCF0M1ktD8rlYdP5tEJLrOdicnca7rbtZ62GxMqODJQ
KI8OPwiTp1g0Fia6+2aPwzh5yl5MzqXmorQOyUZ43abjU9+n8jJ3Vc9gIgSXmA+CwA2t5R+wI2pz
g/XPewWk3xS/F3zatOxjFzo+4YauLYbcEkYJUkeXl2yXg0EQmU27CUmRZTIRmYpS2nBmDlrOFZB9
EODK+dGYFfVyFqn7VO4JpCN9ZA3jnoJCPjtrnBRDXcvn+TLODUc3YlBw9kIoMTtlHVvqfG0L5I5D
Nhr8im0PpjN89OaldDLQ/0JKS77nB3mNscci2WPkoCNg7FMH50lbuETTWw7snVW7BTDYRirdAG+i
WijQCAZDZLEEETkMDS8cEvuqRGkqAXAfXr2NsIb9ZZFS4MkYvwhJGsIoCtyFSOgUuEwYbhmyiUqF
8IZe7g6Zatgi8bw+pp7dPk7Xvh7UCC/+2Ih/ezGSgIl8pA6fM76HbH/A+j40q8weo46lEtZMUzRp
izreuWdZDHOHA7fSlJM8Xpud65QDwOzU63k4B5deQc6fKvLxe1qjXZ3NimzX0OTYa7qs43ny6HK1
LRm3tgWAPoyhMrG5EpMr6i+8k4Iwf5BZ3CH23sS7nibZZa0Q5wJQvI7f2I45W+ivfn83Z1H9Wibc
+lsqfg6iROPrllCZS2txCMawHQR0J2wVH8AGKZxhicP1lgVxxY/XWCvZgszwyvJAXThjUYDlvSuz
pPAy0vur5Dy1bHofziZDG2VbiRRNk/h84nmHUoDxFrT6VTrMv3MmlhuMos8ZzsuqgArPxAE6iNwo
gBia7LKGJoVzrhHvXVZOqH06L7gf5TGX9ROlj2bV3yBFe6ZDDyUUgkrHpCB/HpNYODPOa75IkiE1
A15Lg/G5C5FLQJLu21ZdxMn9hyNe5Dy43JKZj3KzGfGRvxPi72CVa3Nd71ChZKiw70NKKJlbh4+c
BSFBx4KdZynNa4ACv856w5Irvtsexqc0CoA3cr96z8CM5b+RMeElXwkwAdWIOD6JvZlC6c2DBFHd
uWRSGwEfFs+gDKvVDKn+/Sx/vOB8x/3/zjZ2N5R8/7nVvDzl74oGTIaue7S7cMM/R6l+12mtYjIH
7yz+5D63AVh61Kt3vJBGWj8RUQBoQH/+QzFxhWzuqgddr7ihw1KyOF267ks5ZL4V8MQ7wbytQLFw
KARNMJEEa2GuHkaYKNRcsI84PsmihP5X1cHSoKePhapBGkLRz9Rt88PwuuWRiaW0nqaJqymLCnTS
LgK9+Iwn2Uyi/U+RreG/+P7Y5jaxGQLmkYUkYxHWNSLz3rGw38tw+n2U4rFRxY12B8CEfZpAa2Zs
0PtwBw8KGgfNh0ZTgnk9B7A0Qv5KeLA5iNG0oa+r+On+CviOdHgnJe3OG4jvWqt981jwVafrkkyQ
RBgtjTMBoH95fWSrClrPANaONk3o8xb0mzgsatJugfTQ7/IT4jF9cWK9uxvm35zWLdBUCe2EqWBl
f5QS8tEZ/GKr2jNG4xBf6LvvOpju0qIxCxTrP9cNnXA2jIq3pyiX8MZiUARTSNr74HDduKTmhHja
lwNNhYq0dPIp9YsNbUcBDGDvkkd0rZn7uTbA2bNiabrRtHmeob6WBk98U+oKKD/DU/nge+7fQ364
rrtNLQ7OifdckSJpyVOeu/u/e8Ua+PDarPoNc4LhG+Yjjay16zendCy8fbwkzGWuudia5URH1ufI
udGqHcbHJfXx8/tWNxMgbkDIuZ5y+hXGHBtMjnP3vPk3sgB/jZUZzugAvtd7KTZV1GIDJoKcuBWZ
mRQnLMZ68Q1nbZ2n37gl56RjHlvqhh3Zm2/gi6bqB3OmsTmiaMp/Qf6c/YtLKOx3LW5RqFQ2dTpN
j7r3Ny2PB/ljbKwxC1W/DNJ3IuAPYEiYyFcNdVPbdm/tosXHWnTwzT0yCTJLcKJT9OlMwtgmrdiZ
ohDvnMicyIUnnFiWfvlUuEJFpTjFgkW3Ij6TwKN5YmjBZPCfSsLnU+6iiwonpy4euLWT9Nr1kLA8
xHRUuPJVxYW1mr8jTRJqd6XRnjlZRJ9EDp6jYAnvpdQYIzcw+hgb9VOS5zjvJD4Up10ClVCt/3+I
cUIqFDEtDlgT8lOSU5rhgETR62AU3Y1/N/b3dB9YT7BwqeLqI74ovY61q2NO1eyCpIjZN1mobvkR
6jGNoyYb4fCgFOCK1gnDlsCi6JTL50mWxYykZ9a0Z+Q27Wv3Luwv+J86nFWdIgVXwP4PFXdaeB9f
SGgR1/WmSJatU3d7FUS1Ff/Weu+uX8mRGzTi5H029AAhG7BGZk4HzD0q9TyJooGWjVeOGW5zVi06
6298rb7MysDwLxqcSvPhzkAScaiaT3CqHVv5NQVAUL+fxJaNpREz9V9st3IWsAEWEe2y6O5Zl54o
KlarR1HxUUsegcanNKapC3JO8gzVyiKUjeAK8BmyP98TDerm6bagy1YlbQ0sNdYuMxbA5wk0ZTEo
EORUhZBlc0g3Lw6488HZ5WK0g3Hs1K3Zng9UjrC5lSx4aEs4J6opGOs2lCxjj3XG5d71PbImmW8N
vMU4seE6hhoNFLO0ONu+tL7XWH/w48W9s8rbNGkUfrmfaP0kvxkwhwr2C/uaIP0jDNKt0EU3+qQ/
8g3jI3Gom2b0AzT8yod+buB6isFmTW9TNrUxUYBAMbwD22W8EKTV/e4JShoz++1sIr/KjalET/Lt
GWwxmUB7HRgu97DtxFWvDvgLU8jfL4Y5QPQjDZSSUoFGAisDFghsVNHHiAaXALigXv1lWsyq9av1
CEsqJ+TGXOKtUxEjRsfI1Rmah4dcJo9gb7pZKGT1/uRZD2/+i6fSYTfHGH3IBqhkJmiWfrLnjJL/
MeFSUDLdFh5keAPt7bkVVKktX30H1hozRDQolnsTfUXn3BhqA4Lw4uPSCNLX2m1srpjI4rOHmYXb
eOL/cgLr4D86Zua7hkPf0F4Z7bkkhDuEz08/OFf2ZgVnVh/uW3BhHM400/+0nVBcOncKyHbSEsef
5IBw2YCoHXnbaAk46rzzjYaNQy9r3hh1GdRn3iE6q8jKIrIqCMU84UwnpCdh6uG3zLuG9Zk+PyAI
ypN8MSby44pruZcxgxmje8vLko7g0up9/x44WmN22ELi+ZVpYlF3osRpEPHvn0QK8oWkARWVpDxh
35XRSSItG4pedtABQ0Oo47rywCUh3+f9QTEM6+QaErI8AX+I0ugltRNKW2fIh6KzYOXjZCtnm8nL
G0I0a7tYZPpEX99qRhoVLZgis4SgCUFnSvDwn1ATmB4RzIFqIQOhIU46bCHPliBM96I/e2Y+4E4q
VtGjC8pXHjYo702sve3uHiktWbVaiEXL9PgcNzjuZB5VRMwt7LNsb2xsdzga3/+6d5wDFDITiKAJ
eiIY/8oKGZh/gXwTTw/Khdl28nnP5/mhX8s1vRE16wiojr/Q6ApIQD4MUoECKCKLlHzvFJ3/K+1Q
1xBMc6kF4y+/NZdKstf35oH9R+gZzsMgNgJC3hZMIHvZe5srSCKBlq82ogWmBrZ46alsPpOk9WOI
N8E4slT2vn+WIkZwJydf9CpE2A+iYsVXmMiWXRY/KChBgaIz7Lw6HksDz+CUCrAjOHqiOQ4NDs7e
6N40f1QXzgSrmI7NjH8qD7GwZ9yk4J39DMKZNDRk0YQgKPbkM6HslKCrF+a+K0w58UPY9tZkLGMr
gSrrYtZgpPWJUIH2XUdcKPfOKJiPlcn/GzAQFS4dj8jsEpvAf+piqlpAZrxH53SkdZnzf34qRFNu
H7CsCA+VC9ydfkBNYs0icvs9wATM9qhwBvGvpkO+yCm11F/a616/bmls/FpdvG9nzClIT7m9MgYB
/pIXvvHchoJMokT9u2DUASM8Krm+ptFA+KbnLpcCniSdu12w/hu/abfPx55LXVrTc1v0K9Ngshf0
YvW6cQ8Af45yZJj/ftWovUA0I4X606QFFBsxSflA1bMTF/8oHW2iAZ4knNcas5QjIYk8DzYIXDPL
KBVqtz4FopilKtkr3KNo/rel9CSs8zkWHSq6GcdWpql6VjsBBsd21X0istlI9aUsXLejJePDeoRg
T78ZwDPnG7UuLeAjKO6J3V+fFdrzP1jNyW2cEC/Xk3dA/MHZEHUJca3A0Y5kc9WF8/FHgYnwChnj
ppDKTTdgiIziRtxWZC+gFDbZeRTSZ2FbIBZSvCFqtY03k/iaJ+AxQqa8YvSbszRqyHXOytC+HRij
JTJMkfX+6NkznhWQS5QeqmgG2vqqSLK/REk8OxnkPWg23GdGSaxrZs0fkUSG6zHnd8clOQydXb7h
JvYSXacoALasDvvavudw74dcRna21NwcZ9vrHPtItZ5elyxZXIn3r+8SStUlKpmtdKD3cTo7ZEtF
y8Bll9UylM9Lw8koit6Sj6Go5iKbW298GIpLZyhhtp5nnixkWqnJfaTsskQkMi1hDDgTiUivIGzj
AB45BtS0FZsBLuLEawvgAtKOqYfsGRyDdv5CGaCYxWQyUy3JHxz4bTdIghGn2Q1zsblX7FwJFc05
bNkk3mEE+Fy4WnGs/DUYfu20hDggBi6tncEvGZmrDEVizzLL0L8mIZhDs43LT5vWUIkErwfU/tah
pSbFxxMR6/vq5JLvfqar1YHskJv4LTEOJ7JBYwZ5arn/qjQN+fYhgopqpzWvobIOT5ewX7YZeob+
4HJqL1BNseaPWRvyt3vJDdWW80nZT5W5CqBIl/NdK2SEytMK99UW6bBQ+HcmlA+3J8WDeR16keD3
afYqZru6cLrJRNAHfBtDPVuBURWBOE+5cvbrM661hgSSz27ym8DdhW0h57kN6cDPnSh8eYTVU8Or
I14YmLGzjDd378fltkQJSM3ndqh5G/9nEBfU57m6PKf3GeDR8XN5MFQj+QM0LwKYN4WslSHbZTtK
ASmg0/1KmyhUhIjCDNVSuilCYv1TMrIWUsFSleUePNXzEnGY7Ukxnexm3rElcvcQEfy671ak8rhg
37oZsiWsuNYT8wb7XF+QQUUFQDzBJoWMdvWHZADlzdKpxLsUUPFMXuspMI8bWjNR6nJ30EIOcwsh
AartqkgAQjPAKo1tzXiIaXg3eu7MGngG+sc0da4O9V55+SNoh/3aS1oFEotLK1z4+AeRGexrAs9z
za064qT99UJ0HxEeq+Hyd2lzD9QmrruH0OviBCh8shg1oSXK2C62EYz46t687b0teslUoKD9eJRa
qMgLjl212b32WSvuRn5k8dcrw1kPmxP56J71J7OB9gCot556zKZ9ICgKP2mHOF2B77Nek/vNNBHN
fXt/NJpnou8VMKQjmUYRo5WzUzHpobq1lOHv/94bTqI/tcA8W/hFw4C6LBbiEL+hr2iea6KmRNja
aYxWeOGrdySE60LdLibhwGFwBXGoQDTnJq4/iwbrmTSi/dvNLF7pi9/vvuO1jB5/KyeKKNd3D6nC
vqJcb93hjbJl8aiw+E3A7tRYYBloFAceDfFZJ+AZ3956IxTl8dVcGVwiFxReJbhsnUfxhWdqzIZg
7TGsL+Mnbdj+7iHBFiOuo9Oeha1RQYDvMGA9piWn6X//PBudLoj8W1izhCUNGPwMQM966zzzeKjO
2EyqwiWPu/gC1hlydSxJFdzwyDZZzXk9MwHXHiZJEtRkM5MTsKkcD4xeGTA7iwzvViOpvBKH9btq
ygw2YxHeCWCvAxU8mznm5IvnGx1FQtQrypRkDAQQMlPsvCk/Qe9YWWCh93KIuVCI8dAcNiSpwdlK
4FRLu87+HDFP5HlwqXG/YszA/5nuKEef/Pd+EcUat7uzlkVdZLrdOWcdJIGRFd2BlzSXP68sOS2B
PCkffocZGcBjjOV5o1yP1VCmG5QjPLUXKZIHgRAISZrH4e4iQjqABDai2vkmmSbwx85zZtW9jHY0
RrAVZ6JyAiLa30riI3SU04Pzr88y/T+jKxNIBEKK58jbyNSpC+l2CPGjwwSpcuJIkvqOxsuoXdod
TntQRcwhQIMTO66mYsdXPU3+Qx9s99My8hR6LImN+dRpNY4ntLKZlgoHZIUvquq+BLWMsMu5YSFi
v5dmXAcYdfxgWNcZnsTRS0JoZE6wS8JtYex75+ZMLzt6Bd+rxlb6jK15b9Tda+tJSF1r8bdo52Sp
OuSIazxvQ4uTUgJY1F4+GdWxlMJ0Fdx1/NFG4qJWWOJ7eltEFSmLMoSNcD0Wx8GLjOsOYVB9JGL+
u9u+aKpABQbGw8N9xL8Jlmpl8v93JmvHSGINJz3IOyVLhofbKqaAEGkl2BolQ9T/G+JabLDgM/9D
075fJ+urPsgjt0hOTWnKgsowV4WdgKggjhMjZYVonhCbnvzeCZslCeXnBF4FHeISGPjLSCTjBFHv
FpNhcqPSzYl6DFyYtkXLKvB8hTIdO8kpEHt4vw1X2JgZZREMHzj1IePqzsm5mOTJNv+uyp4D2P0o
yutP2YlB88yGLQ7aSMGdG4xN0vgS7RnMX43NfJrgQ1ae7r1hic09mFlX4Hx6/JJQqgpofeLFLXOM
FKvLhWGp9byO27U1xWw4hTou/F11NrBIOd7TRuLoAQKP3M0l33FsLhKJUqZHX7SiYdH3/PMuJmsJ
jPWF9o6zHcr1Gxe9iA6vkB051h1DuATgM/8fZ/zb4HstAhaYpGlI4yPkdzfEnrgFQHoAFXtW2W9C
AHF/TyAodAajFnamQpO1tnBVInZdq6r69Jp88cS8BJDJl8CXc9ntOM5k7PiQM2o2KeypxCFQaAtz
o28nxNFnOUDBoLJ12LxTCXxxURkAvEjMshKngW+0a2zcYXcAgTQKbE3ZR3VRHHV5HhPA5Yd56HQ/
8zS+tjq0XcoWd+bGb0k1s/oKwpW80NeRD0GqjYNWnoZhiPJeXjC7H5qIgYDpajoljmNxE0UFJqlh
5cQBX4BlWbN0Dh6Tf2V5zUYk5tl/78y4TbZtp1LxevQNkp7r/zdyzne/rxf7drLeHjLy00hUPGzi
0fwE4VJAt9lerDT2gHVwq+k9kRhDeHUQ4rl+h3PZD88QbvqPc7t8oufPtMrr5XYejHjUI1AkUPjD
v16ZiL+cuipblH2bKJXMBcOLrvl7CgCZEYok3e3psVN+vchSRBI1SPDttCRBSNhko/7//6pHwWBk
nDjAL0DCL4ErJAdDhd6N/phiEy1Hl3Wx2Q6evJKpPK5WuceiU3/y515ol3WH1erz8PASJjh2xrT5
0kGxe6GEWA+CN6Hn0HOZDXks5uU+m0glywo/rUm0hPCr8DbaSnbIF0aiubvASJ9c4qIVCTqUvXex
Z9qttPQpWIGXhi0vTL8r6+DhA0TddQabgIHT3sZ8Rye9klBxr/w5xaT+LiLqw5MyZYTTEFrJE4/a
6aosUJQ8juLsera8sgazX9IIrprAYzVpHhUmqS1xJLQxWBpjGbYwnw/21BVrNW03T0j2Oq7fTdCW
/Du4QQGfixORVUyXtbuzgtMvqaNw1WXUIHmy4wvN8QCyO7Gn42pdCIDsTklxluQGam2Del2Uw174
G61RJWFlWwkgSfsPco/trXUowkacPKP9M7X/t94Yc3KmirDRjAyYPcc/tVbJVEojKKK7F08ZYqYS
q5RCqNpV5f1v0x1w0HVR7uxRPKuWKljC1OLmoDEHxHeCX365w+wKRqwToNGfHpGdvpWd+tcYNAbj
gw3DfqmDK+LOq2UPxMgETPNrA5Ay70/xokuhsUxMb2ufUzeiwWjdZ139dG+bUtVeIu3cb6yROd7f
dJiwiibj4g9B0doluxB81+zh/Fhk++q1Ap7v98025ZCCyZvXCJWD13mr3GDHNrFb4z/CYtnkKJ1G
ykTDEKymeZQNYgd84UArlBZkSBDvbY8t+KCLCmT04vVhzx835JnV6YMsXIDYDsoi+rMg2NIdJWsB
fVDJg5QNkDX8DXpGT+OrXvTJsqYzAEeVn5EImLTbL1JSDmq8Jbq9zK7YL6LXmZX5pzVpSMUh1hv8
DVSuKyHURcJRNIezHPPlVekIQJLy7RzMdScsDIQWFHuYyVOymjJCc3HLfAnH4iJBAvI2AfgJD/TY
T/HNfiv9Dw6JcuwFhswBssLWI5MuM18KLNhKpO+KIUKY/q/e6ZMGbDL9MFWfiKM2eoE+ubJ34xnH
tHJsGneLvgGMv5IxHFUR6qg8JeX4e9bz/q+GXc1ijIWq0e23MN0+Kka+qN1+Wi76kn21cMR/5CCB
GyirjGYfKSguj7L4xRR+o++2TX6XW4mHa5G03E68srC04WOiSi3yKdcLJ6mFtaSizOIdP48cdHya
fUbzCj7NMOAe/j88auaTiLUWKn/HBFmdUyGe9KYHnTVXvtMAyA8oN//MlSHXNgjK5/GMRI2SxOH3
B4kPK3nWO4kJ/+Jv//3gPaZZQRCInkHCoEq8I5AZfztVp50O3u29HUG8RKffQk5EpB5ME2qsSdQ9
JgrHraB61yl21JOIza9ANglXm6U0JVZydy/S/CRmNnHpE3XcLlC5jNWWCDyEztgOQHYk/5C1XXxN
BurkLLOuznOTwZn7JIsamifG6i+O1U0tE+k87CY7MH6E51vmWUzflprMesWhsWT+dDz4wwTTijS1
66TLQpIpepnOpPk19yXzvjJ2+D/H6KJRNPCv+qo62XuMCj09KeKwJlS9XowrKGb0coVSBegVaOzG
lDdkkPq/3LN5Blkit7roYiLPjHtvIhpUQjcrGccuT1TKsLEL+Mv29wl/G4QSiD4oQsXOlx7N8BvJ
M5SiUteUEwSeqO3l/bZV1fi7RPYi1DYaSM0MnwjuZNgf4/J6+1y5OskwXsqqyHKD9B6b5CWy9Atv
sVd1yytEZ1hLSC74IKrOwx3Z2PgUQFjnO7uzfDUtJbaSXWKtl2JTLC97J5Y/aa8IdH1KPbak7egG
lhH45QgtAdE0kdq6XSz1BTFI5FmpxtKYHU+1s2qe8qNRftXK+Gf5Bd/xcPzNQh4MFV0aaMh86ZBL
UfbNeO2Q+4XS9GMNaOX0yNTrk2jfGRsvN+xUuRqukIPbANDcGBdIvZ4K+xb4hkuuru21r+hQhtHd
mXcIMljzjugMs2T/C6/NXv4fXSp+55nKfHQu34VT86SetDD0BYxV4mY6jynJkl5s0WhGATssQ6xb
3btJFNSGuYRO4DvGK4MKOsZOMysNs+WiNGLxUIHLKdSzC3qVMCKsuIzNHhLYhSbba8ZITHK0LSNk
bFIGqBMj+E3IctCSSTLeTb4KkRbb5db56fsNi5F/m92d596lZHM6kybPehErCtlijMY2L8950qIt
i2WU3N8Nb6CU6BsYVnsfTSgooSKoNvIhoHhqFAeirMnuE0uxwsHYjq0lY7VhBOOGXz/yRU8dZW7+
fqzErcj0K6GsVqX7w5qwb4CMMOIHGPkK6cEJ9DbN9y37XUloTax9196fNAng37e9mVwrhPKUmEUA
SUAM8ikbCb097FnH61FKFGUb0dKTLS58uMQcnyYrf0cmx7rhg4PeyOAnSb10QdDgqT/T/MsVdDEL
is7D+ZnkM1NvKYnqICemKUfTYmN1NHcEeYHrU/R8kMKeWgECNOoxyxl2K+6YBCnhe6dL87aU0doC
UItyTig6i5wxjDdlQsqgNbOPw6XIFLciGM7fXoABmzQnwonphQw70GpT1Mo4ShtIY1I8fj6qqQq2
zRcRrgfVcrAE5/iaodGnSjRlhtsGZ205JQQ4KI3lJnMp0sA26IruqGqSkYoZT5JlUW/5as2Fc3M9
YaTgTuE0UZUYJf0xZavfBwOoHe6p9xlkBO/BPqv+CAG5fRah3rBF3Xh9n5BVZJlL8CJjIFu7svId
5kfD9fDSV57G7fLn/l5RilcXzdHnl/rOoIdBP8ZmMCdVRtNHHDkvGi5JQtSZdSrR182dyB3r2stU
df0eJYQRaM7ss+lSxkmmBgTEbuTrburCG/sFAsdqzBUCQhvI/wyJMd/wWp/8d9wz/zRO2IMDXyO0
UXSkNTexQm7FIkwl2RKc9XIW57n/Zx5NlYKCTkbl4sJl9NvyGfcQrJhKDh+PDjATMaoe7H11EdDu
ku7sbgdPsa07N8L/nZkBgumZGcREP0R5GMJ15+YjLanlgKMh7UuNEZsLMnhxYV8ZMwDOEWsSijKs
ody45gvIB69maXsXwnLyaUGEVGyCGVInDwPdPHzdME/+uuwl9hqjp34N7Nf7tcCKIE0IqWmWNaHE
g2UHIeGSrSY35OxnhT6EK5RRSVhOZx9GSK0yElv0k0GjYHVLLsqRYRRobsY4CeC36+XqweZtl3Vj
tIGHDF4A0qyOU3YvXg5tT5Vjd0TAPoEob0zljl+PCTzZv/jR2J1DA6sIVer0CKukwg+ntvwyC00d
M5UD7XBhpVkvhtRKMxzkpZPlYSfEz12LjNrGBKXVRDUInqeaoMTZlGXLBjAt8cT/x7qwAS+ZPNaZ
gs3xgrcyqJ5EORoKysWvT3RkA/EI+slhHPmD7YfMvgvbMKMTzW6u8qHqvJi6aYg9u8gpMgRFOxFt
xMMVJn3lYnT36WaMgWRGck22dHirdkbR0ad39Fwz+QYgbYb30uaiwPpdC/agx7lcQfkpd3gV3lVS
/Qvv9iTETxewT97BnED2mIEJalKxfSFdiPUhsrNljRlqPKvXH+bQu3QVML6s9g3MLYYedSRkfMwL
QwBCcuroFACsWc6qx2uPsWHHlI3NY4JipBHrj1Y6jHcLVp0giO+NJ9RtzCsrGt+TllqeRU9qhmk5
XrEklMv0ZCxrrSoOqBOqRPqwWRxTZE0FVgf0vf/rpCYV6zbMwxVj2c+5IZ9mfy3QIJ3As0/vxYZL
NmUnrn+hAob1psAHqtF9yXXBKwgju6lnWA6aXLcRC3HQIlr7MYLcGxKlbzcGvMFxIm3O60CFWutJ
5kqWgrWVxGHbI9lCWA2IAPBZzjBAYu/EGyWCuHItJioU4k2epNOkkxYIUoTnvBq8eOQAm7cTyW04
lYNBXp20U0vLsfWRvyrdxkA90m1KPE0J3W1vzS17mFxagF6SOERA7zJK+u/r2m9X/nMayq4w+sNu
Cfqfxq3xxqsi5xbFljl99yQ6KIdN9wmcF5z9GpfO5SObMtOpWejSb/QkuKbaIVgvl4HOVQD3Qg2K
6skvpufda0RwZ33SFyzQW2K1MEey5x1hGdIFGAt3I5RUWS3bcedTAasA++T0UdRn329ZgWSRS1Fa
kr/+9DldB9bS1lRDhDPb1hUnFQMiZJwsknLxY6o+Vf/DHw3xlxG4bw8IOz5uepkH76dVaTI1ykzN
SGNdjQS9momh556Z4+P5sVnliXU7ssnpIkqUs06wOuEW1gG+/ZpD/9D3rtZDyDcHlMT3OwxHuHLC
XbG8kvI9dhT3AlUSqezqN6gTdaVJTM5ufdjHaFcROfIFFU0k814c8o3ks0auimDMRqMeVO2aiqfq
gIt71aNXo8wyZd03CCEYlTbLcqg4PdOBOenKtSnwy+nBbv0EPdc4hrRmapgwp9zPvKI+NCpfSmMY
ZfNIPCU5bT6PH/W3WiT7eDrclu+xU+HQKJnXWyMtmx2x2tmu1PIFACsxSEKQARIqWBmdj1qmJ581
/Ryk1efK4y5LcCMLtYTvLy8a8iAG2XBKUfijJqC3rXA5oeQ+o+6tyNIGdSwmcdjQbdnhwPJoJV1y
pBS6hhEQpJHKB5G0ozZ746vYtyc7QmWJBklhmaqERNbgMhVoLdBCjbTCB2oamdUufxNTZ58Gymfw
6Vo27Be35Zwj3Pjqp0TmB5jRAaf1aNlgB7BKirlYRKy9hYr5RggOQVgjh7IIO+iZOXHWV7H7YLGA
pVNoGWA0cNNRRaNYB5fmCOBVRr7XxRHuudys4F7pUkRSnPLsBslNqCpARpC2Cxok2ukCk8qEK4YH
BsvNN8JzmTp+oWTz3MdS0hTSTDctqPzwlbtEn0HtqBCQjq7GAGqk30vghoMube0gD3tBdtU6CSZa
cnHGwAhidmAUOamix7HG+ZyZxuIZJTfTQUlh6DHEfJe1w1wCRpxnv8hhZMqpX61+P0YvUneKLxpA
03g7Ju77NSSIoZNoDt2iQR9Dl5YS7kFMYp1SgNjZurP1GOA9PDKkqlF02omq4Sdp240gxEmRRXpL
fEwriviiVaOzo8uNInkrvNwEIlyRjykGJBh4krUrSQzKF4G3NPDfgcQ2ejpSOVZ8IbwwpWFSgaBV
zJRM5cL8VWOcvWO1GaOHGuDL6vKhGASuSYkaXnn9Mlwp/9wt4//Ug8qUZKHtTxoshO508FKLpX0D
bb3SCNjbkBGIim/ffMSmXw4oahMhZB6UHeUkz1mQHNZvMiB2w3pR9FawjFQimQZn72JGFICgglm8
kW6M6xJu+W7gyuc5oLfcNvpB4h5Lbagj3JZhxMphrq5Hk1XDnYGIDjnEILpQySrLLbuAX8FwGm1i
0dvv8Q6MU6bRAtAcVuiP2/XOwvvdlU/tQfsjxSGcXjC0EsDnqJ/ySYfe7p3xUPO/CRYOZS/JN9GG
ySmWAtRJ+0qL3On+gqxqgvt4nU3z/LSxPTSnUTBGyH17QL28ib+gIegSdkROey+uuUfQixeGdgyo
U+PgP8iKTDXu9eD7ubxjNR0lu+DECkAu9BqCrjkAskMX9ukOhIHSpnJq2H3qhZg4CXVlXtoaj4zc
oR+7X3rvuCw12aKUbOv9y6xGZU7ltbnEjwSEJOkl8oS4yr7JDOXpkVPaB/z0F8cew/aVoCniHP/n
8fQP6RwZlkpAo6LPcjyierntm4IkW7mB+2gsxbSwzBpgZDpDEdlWZZ4QwKjRfJr+MxGq5XoebZfu
hgFSX54cxWyXQcDFYZ1lVPWPXLAdZu9O0yQ9Q3OaELP1fyO85LTDLiczoLaxtOoLEa0K8rK6ERua
XEEi9/SEw6stqdXfD+XVW4un6WxbjJmStPmdKU2G/Co83wkuS+0vLF8kWtESiXK7uW25dXtHQIFa
Crb/cpFjGqlIZbi0x2kATXu3lahILremmNrKVukrY3z3Xn7VrSfNprNV3wXGwwMSYryCDxgHfFFe
q+oVQ/Zi6lxxn7RvLHZOIBBMqoFqClHQT7aawhLA3DKVHbfhfR/4x9xboScO+z9BM16qu9elX65I
DeswzvqSMlEiyAOvMPDFqjXFGz/VcR70JxvtXv+QRtQbwbV1tfwdoaohNuiWbuPk2DWWZdeRgMo3
cMAJJyrtgdeZb3mu7CPZ626sFWdEK3uBXlFaFGvZD8LReD6dPirqd9ZXuPQCfnziVsZSJk3IR5Jq
Zlv0MOH4C0uwuJT8SQDmlMmpJfcyl1iPHJqVrX8yVLl1B0nhUAn1iRshIEpi5D69D7tt1SQdpz9B
GwK4HkTvqRlr2DjyiO/KC+nAJVcEgT+6djjnlerS9rffw6h+wozc7q5pty2N3wHO4TxQq7mw4nwp
wEerHpeTyIVX6Fq/PG90O+zTSHiXyIgqx+lgSkfmpkWmjSJ+Bddznd0xHufsdxpVfyqRS5GtMDHR
MqAWR+M0JlktHv21J3Lz8rV6kolkDPE36hMnojk89bkaAo1MJMZyaEqbNBmQ/mjOz5vBl6jPy19P
yQwMW1QA0gYk+JTtakdGmcI2O9vSjBn6F/En4GuCa1UgSI1l8UuS5jfO9s32h3jgkzFxFwsbWh7b
uuD+0XY7K4fAINSnMoRGQA3m2tvxbyQtGlFmnnG6GnPE4mAbeCgyixR8undwU7ldmpC0Qq6eb+ys
XXnd5xd5PIxlD6Td0FoZW0N3qtFh1DwCYEbJbKEZtAw9d8bPlNdOwMO+6o6Nqkec3tVqz1GPNazE
vefuMZEj8EXFKmTyoGXaC2lq0jJ2C1z9Uc3zswwFyKMvAtPiy0QJ3K3F7r8mbjefah3QsSN2T3pY
0dLb2jJUKGZN31sb7FuWHIaeNcgTxyWMIrqLQ6oahfeAMCab7zepmgIjoK+GKghDk8WJzhGKHL8p
tsCfwY02WpzTwWRjUeNo2Buv5zeDKX3g2KTb1AbEcehcO4+kfDmrAOCqydmYSwu0/Nq2fDqCxG4E
3DQQGOoYjToLN1wv72teKXBph3CHcZohZluWBLz0G/VgV8hk7ernuEPOBGd+uK7Jvsb46KWLxHO9
ugTmDD790NZyTMMyJrKuKNKL+jeYKNtCgXfvEUCdMQ3gU1h5QAY09a2WVGDYygH13E7/0u6fwPV7
t4IvyJnVVD0Bfj0CivJ4lv9+DFTqX2cJKPYym3IKaWqcID3b0THz5QF58yvFDMW1dOJz6M9vWZWa
0pl+UFhBEVcKb/Yafd6u/dx2DMVAB9ZHbc/rB/M6C8t6BoLSWmsa0mKykGJxlxIPb3maHlFDUUXZ
oagfs1YrAFr1+Ybt/qo6so5xgUdYSqrpeGDKVXdOA5xxXirtFy0fJkmKoc2kkT0SPyFMoYjJwZuA
OCPMm/EAehU34Qni/92SkzpgsfJY4Sxtgm2PVP/DRni+I0LyTmghgeOlrZM0KYNZetCVXQ4dUtNH
Yj8VF2WB7SsmnXBraMnqbwW6ghbykgFI9GWBTOJzQDWl5yrLUDIfMKtfrp42Tqj52vNFI2S4syRe
X566+lMvN3rqrAS5nxH1Aj0mJqBRXU48ohgXoTs+U8mfhLGUSj9b3l03OV7N68xVRJb+X4RFPY2F
hY4EowS3RtofR5i74gGyQDpJfJf8Jloj98pk9wH8VsD8SEUGLxZZ9XOPXgQu9yQNezKy1uQ51DK9
MFuRXY7ijfUtuslMvCBuzAMmocHe91VjnkhneWNk+DtNyzmiZETZpAtw1Jd/4wrDt41AkCne3FNL
sGmPXjjy1fctr2elz33v/UuI75hrtKDm/edAbeIeVPKDdzoNiK+5hVZMlVpMIV1Vw2h5cw1r/UnR
ZtH+kqEBvDQFfHRMWtokAZKOnHeXB4mqf2d7ixB3nuO63Pb9V5sXqIqv6vGckAMXzzif0OuXYu8M
qgXxV+Lhj+OmN6t58LjpqIKpFeIVLRxs+T6dx+HxLXyQXESaehMChANdd1I+iMbrRqPZZk23dtpG
78+pJ/frwpGdow8RMvfp0rRSWoVujq8VXOpNtYac3TfCEbnvdXIUKWkH+kNLFqNyuM6HeJDv4HPD
9lIqZ8FRexR+zk0QOjrrfXiatvtGJNy9swgvd/CfxvYCgt/Tu2otn3XjXOSU2tPIqTh684jOMaD4
fI/cBguIVn9RNILJ8TYYI2UEZU4p+ycMNxOSGfEb1Pnfxs42HstC93O0VF2+yJf6oO645ThUjTOY
1XqiNQKL0Dq/E2nx2E+zzOr+yPXsWKdNEcT7S8dy+p0zuWqqhAmZM4eUEZqWSEl3m25fH14JHi0b
Gvdw3IJUrX89PIWOsWJtdE5YGxP/eeyEnCFCPOyOalQa/6z6rLP5QfUIkNj+gf7tZK17jYbGjb1w
s/aYlV2YeoNKE4DupczJNscfOs5/dE+V+U/320JSG9J55vWkHRwMi6MWgwe2IlDgOnllt/qKXSZ9
UFWmFCFValh/8knUbmSjCI93dE3j3UQciwZv/HfZRa8+LIYqYlApd810VxUl8k+sxfwG5s55t2yS
NINAJUHVkSoDiOLC6cgH6FMZVf6fskdTbuQ36S4L5LE4YY0qCZgqmZjdB3YSl8TvGUURD/sH4s8w
O6moZzqNhGTtFNNOP8Nj1HV396MYaNtQFYo8vnqlwoR8/q6FuvgWZcOvv87hNbM8cuG4ULg4vGC1
QS+wjLZSNNFejffvlQ8QlFHMEBaLhUhHQLqVrsKY73MVow0M+BEmL6N33pp2q8oKZEfJHJDX/JpN
nazsokmk+KGdlddQ8RV9tKoey8j6qtPhHF8WRhqtodGjalhG8LsNIAPRwtgrtvMfT21gpiZa3W/U
GaStF0pF3ICF/GOshdTstANfMwaA1TkPPsPnJw9xuAzNd0glKhOemzMW9Phm6goYG4cq69/qNwP3
w//tagfrcPtWyz3p8rmIZrnB8ui7hEaRaz00smjmeFBfBMnpQ7woRjRsV2vrH1ot7K5jyQbiVpMu
1udLkPvNUftqnfiwIPEOusjC34ezK0tVFT46wlCyP/V9xbP83iXzbvOzIkmpECu1JKx9MXNqz0L6
JM3C536ZTVnobXqEfd4zmobH5boDvB/Gw88rSrF1cHDRdJhuqfjPTqFj0mmWc2lGwasikEcdlhRo
ZqOGRQhW7gOYeGDovzZDHpIrKILEe+z7VyZGg586L+lqByymlzBQfnuSNZtyZxQ/8wecdUu3JuTG
dgQe91obzFNHjl374vsnwj/dKMDBqQ23WHBALkF8Z8JkNhSjloPbg6EGhuenX9skHYj+JJKLh6gK
a2Nya0rv0JmoVExmVKwZ3qQZkA98ibZ5wEGwBDoONW0FDaPQ/LpUH6BQjWGrmaJhlbrYdjcpQGlg
1mVk56XjstVQrFX0OFRdqOLco6b1HPLN93zwb50IeISPG0UoabX96TtJrrJt1KXYquEePp6x1++x
m+FMz/2f99fW9RH06Gm6ziUdFH+ozUosNmRItf4NC65MZs1czRdFqAB12xYONPkWIOj/idyJ86m0
iIls6Kdnx9olvFKDF5EQntfc9BWvFVD3z0y2SWS93lPdouNX8CtTpT6hPBTWu/f8MgqygvqtKPf1
jzyX30MuvktNzaCiJBVihWDENQ6us6qfP2JaHJy2JGa7sQFTyPd1cSloguu0mj+4qxfles60QkB6
lxgQXnpRB16JUmIiq8Fa5ZsWHBJceoGAJmUwErhqaexIPy8hSeIxAOZ7qUCta61vPeezXr5kHt3u
u9gKethO1ZQAxOJR8nrhC39dOkxXxsRN02AQ+FEkrw8nk/tPhuCfMT2wbTnAO67+N/+SRY+BumQz
EhHVOUaQ5yRbMDRVzbZaaDCgCDD6XingUVf7oiooKABIDtiZJcmnfioDpFbPlSVLhmCGQ/hghFsr
EaQDhpiOLoc9KuXBSNBae50nXWkpg0TIBhUKlCP37mvHtpEBXGeNMYx72vXnBAGV1uMOn2HOy4mO
bf57A/vsImKfPxLcoJtVE6CJihpD7fYXHl81p7aQc2U1j+ztGpSMvxB3PT/nEsdH9zUy3EOp/ovl
U/tH1nt6RUBaS10difGBAYMC55GNVychd+iQRZ7vM79p7FucrvFK9xaHelXAzIVh0MzB51DCCPYg
NwLDJDRQoPR6qtACVMs5BZjbFrsksncnQ3E8ctUWZeTeGE+0VQET63lrAvcrv6qkcnkwdpwUDlTr
EpHckR82Lb1twhClvzxpDShITn5f0qj8wdRUW/iEMPaPAZEDtQWaZkFUMxqR20tORmB6OrY1RGM+
f/O/6TZMrTG7LhlBqbazV9rQoMZNci8dJ8B7z3+vhXiet3GaNS3tx/dwdHs47JqU8clrG1W0Iomg
ZGXcX96p/DaFiVrkIrXu/xtSpahmXpKtIo+H2QxtFiBgihaYSBjJZKQmKuEu/J9WzuIRfDuxqSqh
Y+3pPxEr8Hl836A29CKgIG8x8pEdrFxxIx2gDt+lmsM9jxEbrt2rLyy4VMb3xsxvoIdldI8Vx1DF
8xyZOjqK5D9Vyk7pa3fc8IRDdlRZ56ZaJFqTFe1RUuF7+3DmU/jJAsvyuYsEYPgVdZow5x+4BICp
7v6p/HQaewXXTBXd2Ub+gupgGj6PaeY9bY2ZDFdnEwgIlR2pAH1V6udR6O99nVJ2qY0bzNQ/Kklv
/P2UWt4/1dSgyKAlhEs/G975PZ+8C8LXDbJeq3LkSFFQvEEzhqI05Qq8SFxBsW0YSm5y5iPW3vrV
vUReLT/6EBzno7l8gE2t2ULThhcYXfUNROG3NGsxTEqd46pZ/q/SpH46lg1CVOQk8RtJ9p/GEZxL
jbG/Wnp0OKD8yrXiwxnp+VGvq1AZF0iznrTVSHTbMtDY7fmFCewACOR3yGjnPkC+9XKe0zyTt1lG
sFOryLOSux2/g3yXk5MxyHP3swk6AyJv5hlOEAylLXrbzi5SF29l3zP7HHLLMoGmsaSA9xf4w8B+
31X7GIoZqduZnOCT918bPvX0mSeLEa4tfgEegwgITx8I94oVdTSvRduQDu7kVhYyFGfpRLCn7han
wMfCPSLpxxyNZ+qQFRySBykSUu3MqVK++fr3Se6QEvCpYKiBwK0YuxAVSB6v5wrmab85Pas7TocJ
oQ/NJ1UtdsXoznw5uga4ieYmSj+QhlUH4aPQcOHfg7ctU6H68nbGmepYl/q6Cm/fD7QNX10qy8Ci
hcy/+2X/iSmRCTSTVho2K+TGsDk0DGlSqy7f6kVFU2y9qUjWnm7eoU1u+KSnjhUE0lIX8WJgmarZ
CSJZ1wnQIwMvnnEVn2GoSNQAUIMhrU9fjb/C4tOliZxp4KL98nun5hmeTCDlq5UNFll82S688GiY
wFZGUUJ6uiMMhX6IOYyg1TRoN+bmgv1zgfiUWM2TnVd9oZenbYFHugwuMhdV72RGx7QNSjRrb2dc
uTYFYocwL8i07LP0o0XPBGhjkLdispof89rw1cl5MryrJ4lFDD/CpE8fUdkN433x4NT/zgJhA83T
sCpzL1/bt5p4pDweJor4sw2B8tccP4MxY0zjyg1BJTn6qVgvry01cr2qDprw6rJq/KMwL8r64GZC
AXmiPkXFd8Td6WCNiitwrWWcclui7BoAdHaPLf3x6XjW4U+wiSta9jBrihGc5XK6F8gBcbqpSmoR
JR/wwCDmsVWsc3lX0XucAZNlSRxakHjEXPwbcyJUADxoEF0e2clW0fUDjlsQU2YwGC32ORh6Xhva
IPehOiVmwq6J8mnIkEC/qulRSOXUOnrKJYdVqQcifwAoYzMBrnZg2MwFS/Ytlw8SU/iWFQYRS3EO
N0s6HzCakcSwgv/hNHkmp6bjqfQlXJ4kpG5iQkDZ4rFu79IEgftv+LamErI3fWJDGrgqLK+JEwQJ
slYHOShH+DDgrYh6sKWXrcvgvmymWWf5LuOWIYa1Sy0DUV76u9gn9YFC7+qQHBoeCJJpTo02daYv
jxuoNXh2nbGEpM0PBkQLxc7qOtkINi8S/2+f3me+sNz9sCCcdK4FxXcZOteF0oxRSFzBMFkx2ByJ
oam6L42YrWPDW3lN9hb/SxcYcvUbcKqdnO8P7ODGLT59mUJP1wdSR7WlwkaMCeJsMTjZJ3tSjL2u
b1C3vWNXxJiQVQD2XGY83N/YSq/xJv8pe1snfHHpyOLyKg7IrId+ipmfeH7REgC2lq+bKb3ZMv9u
bCy2qWyreBSdFqcz6+b78E9TnF4fN0csn78xEyumPhX1Wexe3flgEMFWLARUiAnIEswlhf4WRjqK
/3tVg9v6P+pXF0XakLHDwC3W4b9q9zgFzt97v23JK7KY5G4AT3DlB+2vuMboNNltc9e1PtU54wDH
1PLlFuBblnSNZbhcXoJYzvrhizidhEn2Ue7NSHVcytGHlgpwP/s5diVRocJAnXbLnxdeBzZi5KFH
036Vbxv5JO9JIEYYKWn6/ea++nGwdbhZM5kotBNcCVDfErsEFc3RQP2YICQW33ZS4fXbSslbrL3K
IyHzftjQJXDpwTym8MuLbG5MB7m7EdjDgRKiaOSwS4pNfjrgwInUulf0me5hzuWCoMydVBOqUKjI
7+cfa9EeCzFk5JdGXPaPN//5BL8VlIBUt3GpUPG1u7Jeo1BWPhydTCte9oN94WFqiMZfg1Agr8c2
gt6WgO7t20fbq7XZg4bnrZ+ZXgcCB0B6vr+FlxUNxLmHU9buMh4QIHjkKJqLz5v3TWVi1H51HUZQ
Azq/uVWsAz0mmnCAleDRrWsRfDXtlrMuIbFH4MyJGLKiHGqs41Vfk23bOI8GJUGtCjzsGSm7OmvQ
HkhbMgWPMpPzlVTN5AIxjXVVy3sTH6OSkcThEngDijV592QEW4MuS31Rg2hhkhOR5AuZAmxode1R
FDld67/rOzZ4Z6SaqHrbnIN4vlq76AXN/mCLJMRUF8fom68+ZOF0XAQuPIy4nUj2BtzYeGv+yZA8
Qt8CNTd1hKQPlaTwYIwTmaRT0hTcTjcOBK3yqkqjjaYJRhCrAbVqyagXruGEF3uaw8RO13D6rFTh
zpu9VUJBD6blaYOZofUnBI35TRRsM+aKiYpsls5Q7K4WN76BjXZnDhe2aMq1eYeg17MKojiKrIIE
WlRqH7XQ8g2y94lcXPyYsZeXrEHHL0h0ToteUjm93NjWtVRWC0Dc0x//vcSwvjti2cRsjQ8Tzm2h
asca8TEUE5zkracFyRcYwa//kDP8MPzquOYtep+yV49MYCkk2BSxcRlYH96d8Rdfi3FANam0QW8u
5hQLCGJMtlhcihrklz7MZp3hy5H5pVUmPbpPlx0/IHE124+5ZXmPnxrVzQyQ6c86Vcnf0JeotNnX
kGf50PVNduJEp+5MlAZZfxsksaITOsTwOx/6Wr1flMbR8do0ahPF6NVORUAvprkm4fFHEx4n1494
4jR88vzV+JhHjG5hghauXuApNORtqLFCObCq4Bi4eFU508DjSJhM81UClwPmOJJxR2rCVSDU+8O8
YwJ642XW4nqsrXIkin6IiM7Jkr5aAkc1acWnGTBrr3Ar/mwnCPPzdLheku5/4giw8BOFp3TXSH1P
yaVmzq9TxzjVEerGqgvcUeUh0mvOFb2ME6stUgvsQ19qOJZSq2t4aewVEvjx6c7AhKvOvxHMZQev
X+N9v04HRi35jSKJzJeavZF+fHr58usZYqE+vmGf9pM/sNEdq2f0NExD/Cq8mj+Ey1JqMJw0d+EB
aMFIXMvuVJ8LsU0HkPnVP8v8stgIYwYZ6TmooP/vJExyHDVfyFMUk1vpl8rVZq1m6koIbPriecVR
Xeqoe6HvDDFt2jGcLxE4xs2HYgb4nilmhPe2Be1HsAO8mZjZVq8tjT1o2gK0b3kdyI4zNXPIIPH5
fkvkRuUiSNDkXTAdxB9orsqkCQ3dkwTMY1gAv7nDBNhvR3RAwOGIvYcd/lTk8NqLBPFHgeMmIFqS
nNS2m0hWXjq7SI3HQSRG5mSZyJR1uN1FPORgGyCsQSlLZnbUIsD5jXWGtvGke9KfnA8fCBEplO/X
H8G8RKfkYWnYFrzlIush0zzbMrTVnOY7uucOEMzL4rvCbhyEE4zVjQqe8sAuHV1WIGWetgbwsbU6
1wFRmq4ThLf7PzqP5Ry/sySg3faPwrM/cYVTCOEKSwl8CqOk5E6v+PIBAWJmlKhVSzJRxk+kFBgL
Kya4LFBrfwjX5siT+koSEo3jXJ0v46xTASo9kYDI+eHK7ppKBzGdWxWYNXo37SMufY1yB9jGzAGG
fcwr6vbWV0As7lw18qkwOI/8RBw3niQ8DxCLsMeeS6EF6McROSTQ2UQaxaI+MTFnHD9YccuWQ+uV
KnOEuAW7kItVdX1UcvnmLWwuIawvYgD0AS/Y0/1c1t9IcGMi/1OPh4tjwzyUpt7b3eB23kJ+EZmM
vEPSf6lXfyEKWHWx13jubS1be52Y1XymBcZh90Wh1j/p6Fih+KI+q+51+1vIHWhcebY6IGCT7Sq+
0RcqJkvXqnPr2g2fUIZhJrh7CQF80+UNSbe4E8EOal3Oc7+v7Y+8SK/O5dgQNT3NbmwMcoLiPmjp
Gaw23ueUbnt0OXO9ItORoWyU9NOMtzYbScQP8iMIlpp7MneIDw0MVcz+HYtf35kCS6jWWtvUszSv
uhmP1PFp+RXFBqLwlArN+65dpdozHIawuVjZLwYoOKKj48Qjwv733TBs4ho/R7VDjVcksXxu6VDW
XMhFocf4mhqVDgPcp2wWFeTF61SmlT9ZGj/YLHVpf8fwC76COokKzhkifcYfUz0y6Zis1VMVWG4K
c3mP0dQDs0C8aKF5IBafgvjBxO2DDt61ByxkTgHZYVfZhWw810nTrruIp4hLMmOnuNI713GYLEii
zJo8h52ueNEeY3Mxezu1tyGkswCsOuJpxq/52cHRdUaQXlcUnZsXrbDet8siTigkBgoqhLKyEPBz
nVXhv/qTBMJ0Hy5p1HyeZx02m7TS5Tp7DXSgQIyD4LXTRSUfU+2e0Y7sccOdKEdUx7QJ4aSO3BF8
KGnPdBMytyPjK2Yj0Bn7maGoKNQ2IFbr1CkONBeyGgNGr3I0oq86ygYY0n0JFpASvnnEK5HfN+gA
p0FfoYXy9dYaLWPVxs8QqS2MgIMlAJ35dh+Wr57XnJ5grLNlKM3TeHfc8qqZPDFJg59Rftp2un/W
nJ+AQLSELVlrUe1F+L3+vTXG9QhHRxXvr6oAJi0/PNPL+IDnP4Iu71yxY1x6cPBKCztGXIJ4vhe1
ZdNHcZ9e0uqT3BhcWLSB9ckDc6/Kz0YdgFJ9rQqLiHFdNHTWRTS3ys2KVx9isA6WAJypXjqEx/Np
i0uGVVW+uTpnK1tlHlzWtuvKGkMPBXpSNQAdBRwZRwVmGHAN6LVg1NM531DtJFd/rwr9u+gfQl4D
eHoWyoL1ga8SoNKc/9H8aTmGVQhIMh3hhJy+VZmKAq/tyweW5Ij0ZcfL2rCAIkdnAuIhad8mxLxg
HhELQLDt9PcG09yGmEPzvvKdBzl88ym2FzdyUnVt2Ip6IJAPvQEEEcIIaZwwg3RUL3kHjZbO+Ckl
bsMU+Gww5vUTfPyuKQFn67SkQtDg724knAhKjE8fMGyQNR3vi40SaHdnvBVqHEV0uvykHUnvcOHL
sHSKNg8/UAabuGoTwQ9snVr2qO4zY0h6o9/pYinHgQazDJtVPFVmkpq/JwBh5BRkdWhSYbNcBgYx
kXGOhAZx+s/hVmJdHVzABM6037H+amM7e1Pxv+zYlF7seqajRP4l7Fbqsb9AvuWQDIbS0JF4ylQt
uhaHvU06owT+8ysf6kJo6NsT0wi3UwfkI6u+NQqyO4lyiWV1rga++NE32E3/cOJR9By3qiqqZfI0
67AOMMcNxmwFI4P5IcLMfBVb5j2tTpJcDEHMkgEjo4jUwfE1cvLD8k8wxaB+yka35nvxGrWMxn2M
Q6jXioWeLJrH6pQV/g/HcSePBTnJifgzmu8tGVQ5zFdo0ZShNkzH8Z/LZf/4tLSu8bKVyjv0NlpK
3iWjmwPALoOwwpsBOEkwrl5P04k1uqePQn2e7EaBYXeaniE1aR0nb4NBAyM0d0pWWJXp8Pwa3AwT
FVNroGxITMraU2ghLtLbIq605jDk6V49wJiUf91o+1lntrPtjgvy2d41Kw3p0aFRfknl3MzVnRvn
7is/HaDXfYJ/NEEPre71Q4ttu+mwaSAsarRaULa3YPFtJiR7CP6jH+NQvP+3fRS+SXHzLt/yP4mP
FgRU/sCe0hY3huwCxftv1Lvo5pOvhJ9FYOAasWfp6DNk2sA8fkoSl3a08/djHC1kVobgjStO7/Se
gFVxYHpSGnOcLO/WpWVUVU24IQjLoPUDLwxwx39N9H8+NV3Pa+Pj/lZwT6FLkiRqg6LBzowZ2EuL
ZqWcfg8VaUIbhIrIpLfBK4d+/1nMp2dq58kaxNy0u3N9CFjxgCHyrH9KtoWfSmiIqg/J7AwlomDE
yiaf0guGKNOa2OfsCZ6YDLZdGmgbSaej+N9/Yype+RqH+SDVAn1wHUVlLjfIwS8fTRqtsesuyzs4
J6hoYo6w1uajJlgODMTaz9mxDCXMhEhq5DWqO28DYqYYeTSut3FGSq7Qts5cDgaqPYbpJY7HwLbP
SUAMdKNfv5UgvDQ7kROQxJ2rHAY+dH5KObRLJkpJGebbuqC+917nkPoCmc0wXXoDF8vIFLYSwTqF
qG61B57YKo6SGktNv3tbQD/sUd0S6YtjjulUm7dlA9BWPoX0foQcYfwHthW6D1URYZfSIqWqwzUI
x+UehNA7QfgDXMA39pJ5d7DNQNBnf0uiW+Az/iUAjOBs70wYreTR1PHh2kgLR/GVugVG1M0xhGCT
proTJBS/uuUzfMOddP5XnY7AF1owbDeMLr3qPF/jb/Q6GdwQNtj5W5+FV9b5QeNFODRkxobFnPYe
8Z7lGQi07N3bq2fTXWS5V1W5i3BTS2zhkuItMw666gL5uzuxGj9wyIvf6kto3CxFhERzl8tIPKXM
7HGvaGqj+ts05dCZXEqxDes29PvCTzWT33cRtn7ZBn0eWt8UqHZbUmFHhfHtfjWuBFOPg75GFYkf
COp8/c8IZiKTaLrjNhLd157lSu58yJGXH0S7QV1gYWKqBaQ3sJVnIBedyUzk/eSi/MARiQd54az+
MD+8w7p2Q9wAJYM7coJ6jynTZidl0RnNjp/wibGLCEWybdr1EoNxLQjBQN4SZIQCSdIqteYOI1WQ
N457LQjzGUGs3wO3G9ge9L7U+f5qVqQuo+QE0D85q5Kqnf+e9tRizuuFLXtCnRsp4nb2MnqhuCdI
p8wbrYovXEiEih9HU7SRR95EYawpdq87Jjp0qIRacHOGyFocDanrhoXv+hjxQNzvhk6HzIUmzU/M
ZLZkZ0npJAaG0xo01eUHGkgGNN3MszC79ZddlsD+y1aKTtIBnJt4nemtD7dHY08S7QR3o6HU6ZLP
CmxQhY/AgOOXdhxHiU98J1lLo2s2b24CN/vMb5E19U/fU7txgYca+jbhiPg+NAOUtlN+vITwL4Wi
ebapzjL4keE/nSWmhfjPaSoec+i4WqjbCjooUfRDN0BioXzTmCGZIY/4XIj0Dv8aRn0LtdB2PvPB
yikul/83JAJm0p9+hQVZifcL05xVWx0LVTfgr8X8yo3lKLyCzpHDA56oWUF2RpOQ3XcrjVbG/OAL
wtSqac5FTNIUzz1dddKxGSgXpHxEYclnxD3dqKSurSpuiboIdb1GqM1PnxvPgJgJHbdGvwhXGhDj
BbvIH96AZI0wt8dgwnPa6zeleDs7UflcVNmdcrXgiVXGVwbiB23LN65IjJB+l3qHYXO6j/WA8KRf
ifovEz48U+ZcrSPuJxI1BEMekoxBBcC10hzu8x08JAfaQSoTcAbUXuM6XYXsBo5TJP3FpofSdYj8
c3BuzpfL8EWmZusbjPho1MeReVGyrF3T1OtQKsU0ZPy6JElMRPyFwmSg1byd5l1JKpZBabjzfBn4
3WRTl455zwkmSwDK78q4GrTEjY1cm9JSuL+Wlo1XUl6WJclGl52Nk1fEiAdeh+vy0XoAAwC/AyZy
IcQIHjgyIVZJyP2St05KGl8G2d/m1baeFn8XUMgGosU3pQn0+BnFkGVxmgsuwtGpLtNtBLAo8JMe
au22RLdp51nA2a/b2J4DctioFcCl16F1Bdm6h8e70whoECY1heWWuO4Wm9dF2ta1HPRBcknE9MGx
b7NhJQC3z0bBJ78Au9Mq4WIh2jlVM07iT/fJwL9X5IMwz9dlI9b1H/rQzxuJIEQIhbLDXhYek6HG
KUBip1TuTqJe398KQPc4Xf1jdgppQ5Jw7VAvasrFyD/GsxrNO87Dahf4RJM0Lt9B3Kj/eZ4sZoD5
KDwvIuUOCUxfGrIcSdZX8lQLu6onEqsaddpeWoXIsmHy8IPk8MXlIHlhxYsxoe5wvaouCiPRxI/z
67s6ehV+KRbg0ww2l8PrvWNA1cnQdtPKRqWrlyC1dbT/te9zxZUESAldswrKHYPcEgh+aOPF77OZ
4Q/Wgrr50Hg/lrHMvDaG3WgZYlJsJyBu7iaxf9wBcuuc/rPF53JqDrCv+YxGIl3cRoAt0gf/KihA
0KY9VUv+LKJykkyLi5N4BWAXYrhcqM/CHGShVRNLJRbfgch7KR8zaLePRexTHoOxdaSWKaoxtmGS
DNkWFoAylICAyzzhax6Q8PDW2JeCcmCzbaT7dPnhzsZQgt5Z6O7SuqcDxYchtKp9eSZdVRmI4/uf
P5qGZRfsXO1y+weovg5RLHpgJlWsJjch73szLPKO6LSiORlT14txsnQiZK6mtvHc9QwXBakmPhWO
ut7I/MDTrou4dDzbyC+lBV4TwLlfH0pu0sdkO+puMnSo0WvupqNzRXN2KlwVbJjaKzhvp2N03jAX
x8C29ma2BrzasnewFFtzlVpMEpl3E6yzNLmyOPLLVQWsAEHGyTL7wqEj5wWHoH+aEzbq9EP6+c1t
eL/9+om+N0GCCAolFTY9CDAoatqzpuxZv7VLPKApejIFleGm/S+uNuPrN40wVLw1NxANn6GGepSQ
kI2Apx09e7RExmd4Br/PIceb3earGE++WrRZaCZNtH5B1E2tP011+n0Ce+zLlnNIw2hPY9liHqxk
K6FtErifwU5nM53SblbA4EThyUjEHk2hjVG9R5/LZneEp+CKFH1k5IaOjsonqWH9RB2JD2Dm5pAQ
rOvY86VPhVGaryS73rmMAe1Ep+pqlIK3z9j/kEVGw0iRR68YY4Ka2bYsa2oGjk6l8wBvJz2Lgz/0
XwHEmmFr6lMTCP2ZjrnjevFPIoT5T+IwhAy3ABxH+WhDdXBmHQ6G0GBS0T+pYAHpv/4H+62djdTo
TLMvPQ8Kpj94GRYO2dXoe9dRSlD3A9r7pTbKms4kvTEWiL4pTWroTAhTeyOgg+r3r/UOHPJhkJqm
DN2i9O+DKu2dJ6xxqqkTdBhTWiM9/gr4O/xavyeHlWHS2Q/1M+kS0ajruRL6wMzNwE7a30kjpQ0t
NlS/GUiRDIUucMsIC7tJgPTeebWQDsg8QNsG6i1tlyAgKOjUDoe5uypx58fIccubs9eg6Xly5iyR
09hbJ2L0kCkZRrKhnx9hC/4SPM9JrJhWMaLzId1Kbdl1kjiJo8hRxlXAnjZxoF6epzTiSeBIccWI
R/1nZZy4KyjnrS5l47hmDBP+xr78s8Qra5hJo2iEryfPA+GEZVGJwdFjF0NfVK194eF7KYlVMe5u
UxoL0O2HWc03wmXjFsYwaAuiErZHZ2dV1Mdps/bCeb9pTDYw0OLewFf9cyiTS2obNnlwOw2veTr4
RjfbvAbP6itlAvlhlgSliBdXRvHEH0ukjG+np6N6iY0T1qrVDkcjZEaFMNmRdZ6putVjCxp/UeAy
BTZby+dbc6GJISsa8XOLaC3LzLupr9xJaPl/4KL+f/4hBHIyM+r9oMP6TmQ/YXd6MyITfxG/xyro
ysAH4qqNMh+XbTFiJRTWbt+9rGaLi59eRJqveqilyRUyLqGFOWDxoDuNrQ3s4SvkWyKJw3OPYmJ0
7BRZ92kRKEVfCIJ2A5Ubbz74/Kib4+hsirIwL5GN20BGSFASIEfmZMxd0Zn2rcBSUN6XNDss1hF+
F5eSU4lQrEv21G0iXCoyJM89wuH/O0mP09w9OZWzKBjL6OxnvuEMus5asMSe2AUPd98FxXsIXa8b
3U7bS7aH64RPpeQbv5HkRqnZQkciHi6oXxiZPYT04fw1hVXDqr/3cK9aXB/h4xDMuW7/3JnIt2y5
AOjmGgb1ovDAi19P9Eo8xufvxqTf75c6EGtP48eTbPJ6VPoiCHE5KhfvCnP8ZlQdIuGmAdKrxzC9
yOSm/c4VyL4BidWriDLjzz2X7TEKbFQtWwE7YNvwuVTxCvQBzm0DRZdkU9M0gtrX7uBWhUrYT1fL
1BNzxnyDnSzkLOWqHKLO8dQaZVF/Pi4yDoaTQpKK/9coYr2+vs2fihPIK8jmBJ4FrMTbEMqnbgba
Csoehz3cBnNOq+nggsblwbT+rXSq43dV0uFu1t5M1tE5KyBqq2EsLky37ICVJ25+qsxVztLfnr9h
2bc8eQ73TP6S7+oKlq6vMaLho9ceYJpsCOTJmZs7kXb8SX8yawvcnRcP/X8Oy8nusHDKBuTDiGM3
7zIEMHZzQWma7rwLgcwrLvcYBicnEYfquLwPMlXY16UfJTYX1kouXk76UvLM37s5xffbjTZ2EPdQ
WYBoG89tuXG23RUd+7EuIr40YLueaAZK01iA1lJ/3DgQa0Y+1UF3CTOX4Q7OkoxG8YpX1mC17P4p
HXlC/RFfuJyftMhYXnLBwvMPH9IELAtFlVeeQ8IRz56evkXhmi76SDZRg57TRvJHdhRuTezoUwh/
5ntvJBcIqXp4nsJMRrhKCYbQwCp0y0KlZbtvUBWZ3Amb/Spv1VHnqcXDAn0NrStFHfgZ+W8g8Obc
kVcLEqYofe9AcAtCGfU2b5YhTSsK4+7x7tEewPp+bmeusCC09WmTiXmLqjYlPX+39+xIy7w0xbOx
VFkEc2V75RFtDRstFPiGX6l0CzVAi/3OGzikxVROBuFZffcVacY+H6bYLMRAoOnFBrFmxwQ/sQrK
hhfTCyq7zwNWPmj1q9Gipsl8Hs4d8fHYBD+E3WZnq2n9B+Gg89+ybzOARlV4Vf2gvvi/9/w3d4n3
sCFNc9wDitKtpyQ5Y0E0wpEXtbm+QBrdJXtcbPOCHCnG2oQP82sz11zWvUnfHDs4uqTSQK0qG1dU
eFPnYofWTTobIV5b6yiZcG9DXTM4Dkd8/5mpdI6yrkyVNIkrW4Qj/Zxi6TBQGJx+1NugRKQwIAja
jiiGOgz5fwAjH/ktgUMZBI+FoDWXgwqkZln1g3Mydcw4JSioN2Vv8EQHiupTlLGWKPNIc51OjkwM
v/nVuhgqss5k+AlbKCrS5ITPr/eIQNFk1bpQyj6lB7r0KcdXwRRbgh3tS+yII7nfSlgmhXN6HVW2
hKw0GpgiDXm/C8puHQ2SSJUcoP9FIuytCn9RwxTLg+z9ElIgVEX1dgy57B3QtdL/rtbmpVDS7nl/
ZlWWauRrrFW0vyczgtuWO1FW1+TV32ypG8l8OZEM78GHUU35xjwBQEET2yA039IkkR+x7eBFR8PC
RjLT0b9e6YOve46E99cjloGQy1mPQUbMmFDqOQ7pZopUpPkftiTdDZIS3tJb/KLILIqlNYu8dKOk
EpdUR1lA2FmHhEaR0rwOmc5hnOpVThA54sspUggL0GwAkyJC/wF/2u8VqHmEOHip4PgKdVpjX6Sg
NgY8/2khHjPDO/CAPIr+lcVw15QF1WBCuEU6AN8rtBFtZLPWOs528NBbvlT3p9NTN73cpPUHGiXM
KJ6t5KHrZnrgnHSkQVOvaH1OqQsohh920PkCN3ARJnvhEViSScNxtT4R7jALoWW3Th9W4LHJGMGl
g74fdcVAjSAHHB4sKu8HlREyd94FUrx2gru+GxnuwY16MNMGKRAy+6zBet84//GTTxjTdCWk1fTA
ZF4zJo7nqNrUzmH6XwqekWdlf+ZdzsAOtt7hnHB7Zw4+Puom8DwdS6XZi/tzHgPC4SYNZGOpN72a
wrWcAvIvWpBZCNMeho4H62XpasDBDW7og5n4mxXV0t7mV+dUmnVCAUw/1EK9SpdGnn21xiZFFoJ9
thy4FZKGsYi/1ptOjXnQTjJcHEzo/Dx1SWvaziP5Gko3j3IE40jCumo4WHX0qNh62fy7XHUIyO52
8+ILq+8GVQK7cAyLxZAQ52HnXd+fM2/aQXem7JRS9o4s3qpEh/DUXfQyiI+bj5f/AeGs+Qa7Y4Yd
jqv10O0+94sjCa5vTSUlWUT7EWPY5tCy3vJvOgD/lwXc+zPRDC4zjnay+PJ7p0CJ1H7QEQ366UsC
sZZGe+Lxqb1HfhcZJxz3qpQ31/M4sLSIAnOW9UVmMy7gwZJ+zoJsX2Pmv3Z02NYB1N055/OeSLM3
5O/0SAMAauOLjexroaKdfgwA5Y1P+3OwCiance4z/ofWBTYnYJ+q8f2YuyaEp+wMeAPCQF7N3E8x
f7Ei0ZjpnygkWE5NHDYK6+CSdLdL1bx5NsCKl/4xXbiska72G0qYlRxyOFWkKLYGPv9NM/DXSBUL
CDlwuxEfOc6vEvBzO3lKai3jYJeOVuA6zN1eSmkJreWPetpExXQlg6hyodtRZUviDJSyc5Qce5vg
ef66TusTLvPlTDCbf76wcdvubHRbC4utKu0SIkkY8niHsarRka2LgVQ2dkZSSPf6BTd6bYk3cbn0
44MoOIYzx264sXh5CTD8REV1sfnu0qly0A1/fBX1xnPb4xPgsi8zQFKeKoCuQgljgI2Hi4zdGccO
TKYpIRc9cNjBDmbx2dkp90qDXeeDz95Lp7FV/kAQwErTjM+6a6zlHABdj/9/pjtZRyWtcJ4V5EuG
+kL32Xlvr7nLc2qi43bhvn0BfFs3DScctGm6oTnQx6XcmJqrYg6Mrlck0c0iOhU/OPb8hy+3vUmP
rJezVBOmBn38fSCT0auE4G7//zjbwtCMhLVS1uFxDZwOQGf5Bo6TKNwT0j38op6TLmmINV8vlB8f
KPSF9FxJUA3SKnqwMOejN6QiF9/qDVWW+VUR+T0Fm+YE0qUMB0C6noL330YVI9YuyS3EfLaDCtT2
+8j80akmh8T4wXRXrPwFThS5g9E0UWB0w0y5KU0TglqH/OW6So9X9nSNQd6ZA7H9turHzINEeZEF
S+F+BTskN2+rsbyN1bb1IjFYC3V6wV0OzckCEThvOeYIsHWIV2Cck9Kb0xO5fq7RVxYlz8xUMtj1
lVFduHHDLa7wXmqjccFVe92GboPF5Ys2rVxilCXZWI+W79S1q1qGsU0EYK2DmC5plOidzCJOf9xF
zLNStdswkkSJh7sN9vcEg/n9nkaPNxRKoChtL/4amgHWfr3Py38ChHEgmuFgnOFjdJ5P9b8n58dh
hjJ6dXC9WvtVL8fVcPjX75q3wqkrtU/XACCuv4MC+jbTC4QYN3n+NNnaNyL88WsqIlJf4+b+7tBZ
Sz6VjtFfIp0OUh8FDJ/nGL5vZNQwJ9ZwzTYRjlKqeysphHj1kr+hi+dlnSBOPRPNc2B315B7AEB7
DioAH9uixeOcn42L5bcYa6BwPGdEMZTUdvVu3r6hy2w/7ggDkvM5TRsR9etSxe9VmBrpTS09i57z
agG04HUoi9VZNMfDU9mfbex+HDhQ+psaI4pF3+Pi+Qkz8tLJvc3MBUDvwySj5TiPMrBFcsjFyN5X
2PQNrCiAvo9/lZZxlHH06bmYXZhquENOws01pCEak+s8XM2yZZFXpdwYM0JVWuVMbja0qd4dVZWn
+CKg3LoxLF5IpXvYMdVIPl0jN4OKgxUf3mcPn/Hl7Bh6Q9aqDcfr+sY+/24yIDTeecoGz6jEiZJ1
qULfSCtZf3hUl5RYCHbk+C5scPytEJyyJc4/yz4czFNjG7OM4CfR7r1UXKnHIUR3RW6xSvwUj/xl
xo7/lGObWJMiOWfa6l57YSX9TFlOG4QKRYTfd5jUIJZSbA4zgyUuzVqRMoiFr5Lje+72q84qr4G6
3uMeLZOveUbYZfMM/X4tcyogz0cF2jhOQ8ty6FVXLE0WouXGZz0R08p3zmHlAph5exx9NrkFBd9b
orvTYqhjV0UIt57vrWjK6mY0miLIm8YGFDr8EY2UFAUOexVA0+k5DMXcmtQa8AjNZ7zhSrfUOoI4
RmD4WZ4nEE34lEe2xiPxmNSgDK0fzYiODl/gFOn86bmtiAgwZ/C4Op6t40c5wxwrVgo0+f3+JbMr
+qvp6foynTjeGUdqNB8WH/hgVEc8NeSz56CFN4H7tvXL4FfBGiMwS9az5QS1u2qHHzx0yAUvDB56
n5JUqBZbhKReRNOBh2DhBi1WifCFgN470hR8v8fji4JKvhv7XX+r2Lz8bJFaJzDS+MVGq7OGduN5
VRJE5VS0AxubE3fr//rvrG7I0/yObCLYlRIUzktDVvpMNUpfx2f7fTs0mP5bpzyHD6KV6PfFXZu+
Ui6g8B4HwGCpR7zWY4lStJuPaOGNZ8D8lga18bb6BwYUfK7gcCv1ixwiDpJZMMCbpd5Nzhl+SLMD
m5qCJ2fo/lIEovgfOCBx6vbjy8k9mRLvGIRDJc3iygK5vc0iA8BXNwU3N0XKuhFnlYHcaCkDJ1sD
l48T56e539Gu1m7np0vGYLZqGuZctFeLFQ89cs02+a9I1NvMYQ/4Z9N6qDER27s9yWNVpnr8yha9
4dKDQkzciYOEAeQqzLW6DTahpN/pZ354l425NBo7llTCALUY0QuF83Ix2n+a7wDGFirSmt7XhaiC
9c5CS0dENCfZpWc5LBSSlWlb56px/BfR49VzX5az/KYxFVsCx2qX3vq3ZBARkEf73i7gog19nPdM
au4x/gWXhbOuMyGOBnA9i/7ZzAAUtwsSQkpTG/M3E26sLxPu4D9XWnFfNGL19YVBox1sOq/IU79g
3J5+a9OhHn3SkufYVMfniQ6/msGZfC3lHkSCn7SVmxFdJKKQYtsZFR/pFszOMI4m3Vu4Eha67HE9
4tXZt/hqebsQmfQ5eHdybc2pqjT1ZZz+xOPOpzWREy05uRgafz1Yoy6WaOSnfomq5UThd8eCSS98
oDTbi7q6fCqs+0pWk0TsPMqgbSDtmxmW7TvE6JYdzruIMi9L+vnglgCVq3Xe4rVzQb9dFSLyEFDh
sCNngLnDKnOGVXFKzu1mH2m4FnRHx/knZ1yxmFZgaC/ayfvhTp4fqcSfXmG+Ud4voLl/KB2+zhP+
CTYiPG9uzbGzou3qVDqtJPWjO6VAem5QpvoQPtSDyRiiiqrrpjTYuQrgXWeUZnp4XExRTi7pi48w
cAfJljVuBg/SUtVM593emZnShyOBIdm++2zfV9v9ef5DXBy40PGpnBvZOSHQVjcJ3XJ6soZn4DUZ
3GCnSCLhPQGrJvsBrJrLQOp/9xVwMjJxspF7yu8fZN6PITz4MZHJJg9EdZ8s2q+77TaBb7YMVhrB
RQ2SETpHug3242rHexf6++0lHiN2pXxFQZb2rB1Uq3m9RaSI0s9pt1rFNkmQse0c6MizYrb6o2Gc
LwtncMZLhiTrL0iorTSFI5Ff+StukoqFGwGLzD1jOjtB8XuWlVvGu6o3PowLo2If0ll4eJXhqdtm
jZLl5wPZWjVUjxXxkCNG+kSOzsX03sIsETUJOx0aKW2K8rdkl9WlisxLYDeomh0pjexHD8WC//EK
zsLcJ39wPk6k2QRttoFuKnimAbl6g2viwW38uw269GoOm6PprBoxuOrJPIsrdwWT3IRfvu8mN9/G
FZLND0fiFYvxMVZXm6v59FYazWn9/sE+1+KC4hrGjeZAAj1qERRz/NfSjPO2wQkaW7wwl8kXS+KI
iRhBtXj3vLE2BrBPulxVsOcZqDKND/wjweB2co+v7T679Kf72b/nMZTt3Jt4YvgGno/zxLNlKogJ
jkdIE/spMKTxHGkQcB2roe40F1TgQ3by9Fw8qdWhQaZ4jh/YwL4AHP8VzVwrqgS9kPOABcrIZuZq
l97+g8jr3xLLPSbcNuofylHdzYB+F2QrhlqOQbMbJkwmt3+vRk/hUAYGPfli3wAWbdO3Y3KRioP2
fLD9UGMUQydI07BXSVmfZLTnKE2kF+49VVj/z0LRUwPlCeBlzxiCPDM6tqhNlIIZvqHK9jSws070
oKBN/CG9+RgQtaOJxkzvdcEt0z6zrOSU3oxfT8qnZb3VMIjJimeblmmgIFZVaG2jOf4Eti1xeeET
pqbtDSb/G6aP71WMVhy7TIaj+c3Bxc+mWbg/m1q7v+ofYuVkSH2Z/YF/5c2YG1QBFczTmtEgXwbJ
OAZne20QtC32vU0kIxbcwxYnlE8ixOcaHaMmsuV75lQoqboGiC1tkYF1ehZ6F6jjYbg0CXYcoLI8
fdfJfwPdwbWJxpw8bpI1BjeKFSOZ1FOhYlnNDq28vvI1BWgEZLcQfZ2sMDMCxkd1p/c2PcMAWyEN
+5fgHWB3TVfN/0+te+fThU6wbwBmhGs20399JPfZ94iSZc+Qh5zUlsc+jtR6M5qj21iJFvrtFCU6
ys5X3o7hYup9Q7ZsHSbO2Zr08X7sLlOGYv7KNqoNQqmve3JgDOtsPIi8d8XvKXg2hm78JzK5jSMy
cW5442Mw/dDby0O0X7Lu2jnFXjxnnmX/y5oIzYuwbV4+Wz9Cvcqef9IWj51ej0gffNLSFAMEIIqs
hZBDSmWXmqOwZCNTHZPXPcmHj2aabyZY1lOgtVhJsGc+p9EENKWnwMl8FKNxwvkZsrFxlGbiRV2C
UZ85Y72J7+Q1/wHZ4DP2wWQflrsMbzvryO3KSESzTyt6h+OATsaEteOoG6WGm73P4Z38mf69Uv0N
13PSgJvZcqBQV1HfAbUFUEkig9fjocjtayVb06yy0Bk5OLooBm9esF57WZBy8myHMcDUImGZQdYZ
2sCROdfwb/pdLHXdf3E0pSMXM5f+79IFj0Vq4yTTjyXJSLpCm5mSKfHYa7Ap5EuVGyWC/R4mgis+
NBteZZAHHtSE/iEVIy4w5mhKTNXg4WIxuPJgJ/a7H9We49gAD04up6uc0b4plf4CKi5Xff9JsqPi
qd4f6I73WUVRPUcjb/pw5Jo1G+s+R8YecPyTkmJ8Bn/ynmTqgNOAI/SV8e4k0D9lvvxjFEqpZImD
wpc8X5ofWXHX+7Z+c9kz4tC5WN88FdR6vlOEFGQ8hEVFJE3h6G58RlpvNNdEAyy5XMBN7SRAFYma
ZcHQL/iAQWGWad6IRZCt1zQ8moJQdngly6/Jabt0mVNQ6A26bPRW4aEvX59/i6KQeddJLLRBkuYb
K3TTakGavUrc/BiPywxHEbqJokiCP1IB+ml4i8pEoUHVily3exU/5M1KhMGhq5SCR1KZe/JgGG+e
abEWGCvKfjnjUeb30Ur3uNnCF52+SsKJZFWQdLkeyWq3T5G+Kzt6HV7JU/yZhiiJnBTDF1ng1FCb
x7HGcHunlXzy3kmomI7fY6AXU83SxeXDMy0EuvH8LA1uGlf6IZxsQHn+NNBbjp/xBkkf0IVdaF6a
k7BpKl8jr+8sdI+LDiHEw9BWGg6Ypnoe5Hu4Jcpr8SPREpz4S73Jv9Io3ZeKITZsIskP6pL6ckgj
QGy9fBO9Oe/CUmE1nEpeWf2Zj+ocw2SXyQ+DWxbkYytIgM48nEx76JFHROfeiOtgQWz5wz40g7va
ifro850AwrCYqljWtSwvGESexTPnhBJU92Yp92lMzMAeNNGyyHpYFmu2bMTEDoAIj04ZTEYXNhYV
KrPzkGQlbux5QWBhYz2mqt5wCTptgctU1ayN40WFvYYa+/ewQJG47FX1nIQbxzrQaloBty1DrhvU
fDQCvumn8Znz5p694OTsBnac6dehDmGWu8RF4V+Xe33vFJTBlpYcihlyk9GaX0Xeuk82e3j6Kryk
0xarEpdI7QGqoVAKhZLZlpeIOwtcxWJBSTuA0JVR+N1Qsl13hi7ojrmI748hoCeEmKuHkkKnir5M
IRHjT8xoPw89EgpQinGXvqb3PocDyGS2GRO7QDCm2DnkO/X/KAlirvXGXW8rHVTNTpTfUYIsSMpC
TI5HDxmDqQkYmxzc7sE3DWUfp5b3exJPjNg2zMI2GQS7DwvT9XnbFCeEvlbc7xxOQ7Oi/f4XQZ8O
bROCZUCS8O34qvcvjnfgCmtc25O/Ejz3Gc7ni/HGRcr+zbz2cVWCV7erLs2dPZWUPIav3RJYi8Of
1docdslx/Dwo1gzVsAVdZDA23atR3PzwHPegzfw1lqrKXdfvk0TWgAFnr8dAmzK3Okma338nnJkU
kZfanKFRTjfVGwL5k5K73Fhd9j+4Jw9ruyPhf0/sWbHi3grK5LHt0/w573lLrk/TaHlwJBPUFb15
gGWqThCxlPQeTErmPy4QaYD2P7WRPHPN1wW74Gy86WolwI32mx2IuPiWom+rS8vpKAO6c5gH7STq
4qp562NmAKLt40EB398JsopSiCuYEkILUkYyM2HSXxUPPSErULIhhwuB01yxIU1SyEVz5qWLUIoe
hFXyII/9q6Js3RcD3VAoTjxHHp83wSJoVM6gKhIOpLyzdI7lf1lvLUkvRqI+WHZKSkxR3daIH0Nr
l5saQR6QIyz0+5rVsLS266UMIbLr89HL+bdnD7JIsxoUL4s6ISrExgRMh+9eP2RSAS216DZAhoza
nPrcVJwn7ciVs06QuY4LCJ4ufJAQUZJ6Feg6iZmDcNpj/VeVLAbC9E8oOEgHl6Rb3JZ4hmc3KKRI
NGkwerZB/sYECKJa+lKWX3/r7I5ECY6V8+uf/2VNl+786RiATlG6O0d1lrBDN7MusELuT6M7WcU1
w7LSaqHBxr/8r0Krzn0UJNNVqTwIF4b0fbX86beaBtQ53BJ+08HOTi3NixaCwr6LJmqeipgFsOT1
NFT6dZ5+lqS0UOqiWxTI1dztwDqeaNlK4tuFTFf3yIHlFeYAudbm4k4ASV3wKFhOAtL54BoJCWdX
fjp2lUB3WAyYQvJtXT8j9pXqrE7TvX+nvy4B1EqSPxs9IPPyrCzygp85azcs9SPBEyEzFI/Tj2dC
cszaIsc6XMUevTgPs+kjqMQya9mRErZhNnRIrSnYi+IhtH8s0Je3qAX8LtuxYv/14/gthZJXufeg
GgMx94KvMLogGqHqNC5rSra19ejj8O3gMGPLd0F0aGXhbPl18qLoIpSEr4yj54DqPp4IZ/ZYeORB
JiOS0zHVPydCcUUGTWbqna7fjAg7zI9QI7iJ1bZhSV7I/N/8l08KA+yrlQyph8fY1+eK654OwGBj
BK4dzMP2PqJZB3T8oMR25ClK6yC9fxvjB0osjG48UbosIPIb4kTwFAL6S8Yng8Y6RFu9E6kEUQdj
+LX/dhvEj37tqvj2yP6XD0b8wzwBy9BJwD3gXJZNbhVncQl12AHo98GJ0ETJG8nu4rUUeGBRxX9E
KBZ4LkNIZVo0GTSZ+m3qPR7Rg2LW9VkaKvL4B1qcrALq9ozPlf8kyLLZwlNiOQ5+32BrMIGXFkkd
nCU7XQsb1AudWco9ZhMCB7fOHloSpPIJi6c9gPw3+OINAd1nPTsGUKf+3fVqJr9773hYWolE1CqS
yADi/EM1zFjzNQncYwf6Hnxfmkua+F2UALLIfU0alzAfSQmSy/gL07Nt2JinhjDS+4LDsb90hBmf
1aSHw6l/HNovaRAERtPoauzm2cy9cKoE6G8vDX+WusWlwSFF9Y5h3mAit8+WOE8kDyfmePN6ubyk
jEH88WkYHZpomaJrXm71cbHc8pfmh5DnCyQ9FtGCnNKZbCANADCxBaOAhoaF4KQOjuRakCNKgr2V
z+iWDLzYhb2J7kvs1mNQmt9RMsgoqqOTssMNo5OKJ8V7U5QgKcmEG/0anHoV/DpGLrUN8TCvKzMU
YcX8uW5/kPcVRao2ohdMQCioCcsuTqHclSabqHU2h3tIAugsrURaTPsQyQyK8BX3ZpOu2Og/bO/b
6Qbde8t5uRE/pQe8QnK7buFhHF0lmdibxxzVbN9MDs5RsSY9Se1bYnRyLTlsmoX9uULjY5Q1lbRS
B7+OKpd2PfFFWEoK1CxprCbqXmhmKnH0wvPzuy05GovfLPlgGS5F8hMKfIZ5ZNM7yWTOf0FJ2tgw
i95IxbxhoKzTpsNmv/mxY7jG8iVFBHEhwZyl6+Kf9UsMPMm2B/z+t0d2PCCmPMp+FpPGr5WKOHx3
f0zFB/OMTUwKlZlMohXB601OBmP4ucPVgqVR2Ldu73r+gllqL1/0S6Pz8JQ/0VOKKo9qRpHG8Zyq
owKLEVZi9z/a0xMvWe0hNrYMnH/me/ZQWdZ97y+GhSd/si4rzEB2yMyLnqevRIbtqq9oEPckaUh9
z84lKC4ALnu4dys4lBRudZiB+fLZBIWN6Kl/ZW5K8kneQDgPBLYLWBed6YHDin6aD2t/B0SRth+3
ccijqO3D2WHiC//+q59IfpEtyrUXhJIUl3kaBZ6lBcjegwAkC9qzJZAi0p+97EGfj7/xHtX/gkSC
XQpQaCY66nHDKtccV7OLtJiLazzhn94Db0a3f0m5/omd/FaX70qquUiijvARDnDc41GGmKWjToie
lWypc/brpb3wbGtKFnvVL+19dzUPutlTRpAgnsz46t5e9+QpXk31CZzRmjB244XvsOu3sxTVjePj
+OXD08iEZjOk+8vznMZThEaaPx53zrqJlw1/tfMfPn3nopRT1XMrVpcZytSe71thUAUs1m4a0QDW
HzVhRJhDOkIPek11DRKSCbQGx3Z6djIWWHqSdfUE4xKtXIW5/EcoX396AVpmBcJ2fRS1Ges3u2Tn
+Iu/NwwwniXbeioFwAtjTULvERJ9Xk6noGHlZ0KYL+dWtm99TlqB9tYsQv1ssdtZRWd3xAzMroQZ
iS3OecG7KinYZigWvT1/dBp+YjH4ceYoGPzAtExe+mrydIGB8/gampG/MKw/TlztPD/zXEokOmSh
ycIybTVdxWBhfc4+mohh6uTI2pnjr6Uv0W7aAkCLAT9yBWsYVKliQSQ99ZfKGThBvY8JGtbdYYOs
QS0JxE3MEQWXjJKMwmPnBsfwfqZrGHi3Mil35R3WeHIpsxdECs1BCUVYV8piixIbf/cwOJptXrV0
FvbDrJJ2CmjnEvgyg62S9HqRQa031GH29Wl8fY6BPRI0aQKTmjdPRmN+dy6rM6zmx1Umw6dsBqS9
Fx09y3gApoh9S6VwPeUS2qzUEaGOfH1U2ozRiLzvtHMF8TPiwYa358hAgmrtp0BCVs1LN0ta+VRi
/FPHZtxbtRx5X/EWhxB2n0vjWciEgPYAoZfEbYvjcg3OLO7PJAjFIXyC2eUmEldF9Lv/DsCBj8bJ
XnQeJRw7tA3RGa8qRdMbUull128UoDxva0JQ6sZ5BPsDlI6xrfBbPIsr7rlZB9CoM93wv+82T/nV
tr8LlaO0Fvth5AWwtcG5amcbUDmb5mvmNdzOMhUbmBjtFRX5KHoer+E/UZyRvq8GRQxGRfXAaOfk
E9M/0z9udLWzHwSSefxo12w7zHcnO4u5AGRW/tBCQLa4HFqrY67G3yyCmwKy6FfTqgd7tWuc/baP
yBC7yZxTiP8qIa62zxq5MwuQ4vkoxqHdl4n4Bl+kpymZqSkW62EdxyZVhytzrZ9WwUqHckf2sN+z
JW/mF06bRYRCgIO0tPZwY8BuKQtg0BH+87r76bXRRTuCP7pXGyMwm2TykTXZpT9mvh4RQ2DMaCHf
59TlaAPG0JZpvZlSU5hsw2nBhh2ItULwpagiH6EL/g08VzY3lE0xARljtPNp2Rr4BkFu7+fVpNNb
/BmiBJM4ryDxhmVSxh9htMCNr1OWN5VAM+CNJs1H/2evNNop02HbVjmUJbzUMlf++kkwkYUqdsfz
BUpbHqiTBp6ablHvDDxSJr3BJxN+kkZ1xRSEegmrE66u6+UkD1eOiiXyrJa6yklpy5XP4RyZdX7B
d4wD2/8cmvMXfnGzU5BQi6hZX+447Y+NhRonNceHGYeg+8lzEdfLCr+XJqkfTVWczX8tT3dYwUln
/qHQaOkS60IH9rZc+ITaEwrNOGUVvZzEw+e1IvRxwrbZksIbtb8AAPrBgh0/139hZIfSvK+A62f+
pdWVFNTM9xmxlTUkbaD/8ODkGHja1mnMCm6QA9lEI44PpyNclNtdA80hJQpIchpMSJrYl+ue8M3i
Ty1hY7deE3ZZC8Anz1fxjQU1PgBfJzE4VeuIkolD8jLRft6vWJttTqLjQvhKI/rGem8ORXuzXMX7
0eJNyZjhiLOQS5GWt35jQLB2c8GRCDWwdl7AgGsx7bTIEoQqVG+bGbiyNnNXOwC32WixM34mDbTc
lg81W/11bjNVnFjVNFE3qxAL6kNcT2x/LuQobvKvPqrVT5pdnn7eyZSmsaC0W1xAu4zzsaUjmN0h
VfUa92CMkhG2fbwMcpzHVYG7T5YWzY5OGEZ3Qo5yoohe053IDbWY4fYeMzWnxqhnzxTwAJamP59K
VHkYK97jaoEIrOda5wA7Mo/PZQNKFLEKlSCNCpMzwyMgAKm4iq+beOFnBV7QXJEgkvnFA5FbCDsR
SyYZhQYdZPJVzTQuke8gCG6/AuNclGR9Y/l2Hzkoh9OS+T8aWBh93x8VI96mDoTjvMl5XbZt/S5X
SbaTi2EVEYEbT+IydwWgoE1Vcky433mhvRk7i9jX6oDCA8AMFiyq+ZsR9e+tXPUd1rOvFQLN4/vQ
KGsG6xU2JEX3s/pIzRg6YHfy6MV8wpN8eqn4gf1YGgLKAf7iqA9UmnQJgI5GlprFi94Zz9S4PJOx
z6bR3l3WYRrzpAaQDV1SVgY7Cxg/vrQfbb6Uwfy496QU+iH63JRBCYykIUbcgzgblIA09RdH6WNi
o5oPpnNlDd0UcQhFiWamBhV2c4QTExTiG1ow8hRYKb/k2QIVKBso6NYGGCG1wY2qyGFmkl6Cc++E
fnDEZycv4R6DBVmOpjfOfCcXep162ykU39ZGO94/ODLGqQHhKzGP7A+ec3jFIWQR37MOjcB7oluU
HRzj9r81SyhykelpAGmEuAYoLraJThE5+UsYGFUrjQMSw012Rjz0iSBcppH2ARlBU4Yp5/ad1XmP
ZxCK3QD2rtzYWkJnyHv0sTvGR8S5RDIwA+f6xS9n3NRSskVe8VsaxFuBCWuoqypLQNeYVLW766Pu
bINDcv79n7YcRXU1B/zQDmHCvcSiJ/cI8uTgU04AQKstTHMmTDXA3NRRDyIewpn9B6La9glh19qh
ff5QoJGI3AI91znvWIOI8xkKj0mVjGR3RrYBlfaiLgrflCGHxKyvo+Y3dNqxErz2wdYTiM1XIj/E
EcGjB10hpys6jCeKZKZK5iA82JhaI96ot6ygqTdh0E7x0jJlLfWCFPhV7VOPQ4BEytSDCx1jSEdJ
wZMN4HZkjQggMHGs+dll+OhI7Y7LKuoeICeCTZ+ierfqMF0RG39egUDOMH3lgAyD4zHHExKlGpfO
4BhOgu/+SYWc7/ugoekwbRvuevS1/Z2C6ECptvi0z6wCvMzon7k+wjUsG6h6xR1QpuUOWVrI7D3P
fgIBGEEdAsXDQaJL+qaxtIbWty/kfjnxi/Y2VSweqc/ZeWYESEyxtkeINYKbfF3p2PuHfxOZl13g
HQK9f3hBO7Vwq8e1THRYA/LE9pbCq91YIbLmFd3o0MDoarmBzTogPa3nAEW9SA7Coi+3+wvjR4X5
BZZNpXrkZ3XODubzH93xDHEKVpSLTrvsmtdnM6TaTQ2ESIArcqTLEX5xhkhR1jTnQ41JdUxmfCve
aTufgURElbA1249xqd8PQheSgxmXNHWfEVyRC0ESTjCTFEFpHrOs3B4jh0dqbk7R4ami1aAjG4KM
Z7ORDS5QCCYJ5k98B8Zvh4C22cJvviUjNmGLkzouIv9XkSdI1/5mGG+H2BhAaNrOLVddn7TGEdH/
2vsIjrWFZENpAJNRiQKqKuu2Jfrkj941X4f48B3eA0kVO0JAzkkZJt6PjePXKqyGZdkfQ+Czu4hv
jeox2CSYy7gGgAdQ8TZvqc5aExdoBqmG/yJrrkey/yReLpIHxcOwb4Ta7Z2NFvjf1bd6+oS3TD4q
aGO1oXMBrJSD8YfHh1uJMr6KmjOK0/LnV77iQqMfmJh7tulXcTlp9VtgrFIrgsLmdkf86b2zDDr7
544slA5QEJ++CABG4bhnQT6AQUlragEUjZS+WGwFlQyAiMg/Bm/iGYjcoD4LcNwJ7SCQfxeQgYOG
YQ0ovnq6FGJFV/2jFJx5ZneKFBxKYJ+Tce/eajItpMbxKz2EjLj11MnJ3/uMaCCUQV4IPc1lj2C0
tdRVQ0pMgagl9qsfBDdNlujI0j60UFt089nvg5kFcz3Q1bX/h1gs/sdDQ1uBKUwlxFcitDVo+fd3
YFSxkWnQXNCx/m7WUTEfH5Zm3EVH7QfONHiheE4KO9/LfuAsgtHXtDu8igtjuEe5fiR3vWvIkJf6
zUkOax7SZGzTR5SZYZvYbXeP5ARVDoySXdrDzpqs6bc7zoAb7vMwJaYt+zsjQYObUqRMfyubXb5a
HELa+nREeVN04wJDlb4z/o27nTTQAG2FXRXwxvhVMbIIjmtMFFljhuT7lcuNkqKB1c9eIJy0/sY6
JsRd3FHNWo02rfygVKd5mzqiLLv2sO8qH7W0VurU7//jVSEAAeo3HqHge2c/DaMqgt09kqME69Ci
4XYSKQDPjcze0RKP67Kp6xrxTjraluJOBvVIG+LPjHz34DsjjtI3fp+fWq2aGfel3jxcToWam2FD
534Qs2X9p2I7YHaUu6DgxBYldx17+eSTCvJeUwzhn3biukVZxoZBSGhXsIGvPsmPVBPi4QScB1MD
lm3UwWS3uabn5O+ZXJU73SFfk2WMuhoZBElJXzqm7oDZjTGB91AGf262xEyCcOzonIIT6YpVsAxr
JpUacBYTP/dNhktkyydpAX6fKESGJSVHnfJtwAbpsq3OJPfhPP3m4ezxAABCEaAC5uThnhmmQCCk
ylm6zbiq5BPlPcJZRJhJjISpxNOtH6guNm0MlNmP+ReErr6wq72weie5o0VuN/6L8nY7VS26wk4/
oT0pDrdPgLKxv3Jmoj2xcXLsNUuj/u9FDdXQA3Jxyh9jnd336LFm2weM7Rymy7LZudsBKfnfUenE
1dQWaFLLZMxFJ/h5W+pay5UWUvRja7MhVNDHqFpNTkKoq4/EtTfFJeg+fUvBqM0XWS6WKO8wtEdF
5SZvQO+O1hQo41irbOAKp3Cib2f9591ut1A99RFjpdOA24D4IGvEGv2Y2gAodsS4+sGzexNM5AxO
E6+oLRUPqqzkcDnvgEc070VYexAeM6/QX51sdIuoMHEGbE8atepmFpQxO/QcAX4Vc7JqafnQxFPC
oSGz4B5sn4uwWCPDN7Me8gOCK81cn92oEbbux+OSJMPXcgB47332Ngm+NOjPIc3hmcX+TGwSUf5/
J6VTPPS8UEm1vs6OE5jvkIBzDwK8ZM18owvTHkLd2wEvRCdao1NlAQ6o8K/IGqjPqOrFAC1D4sJK
+Z/NsmjBEn8x2tVfLKuOemntXpiRBLYsWg9Xa9xSuomaJUYe6hpgixxj/lpp3JtPWZhcnQFZg1v9
fe5ACuu7Y+8KuR0MamegwSc6f65S0g++W6pGlpWk9xv8nRCWW5uy4ssP10xX6TatVRe09Fti9sxk
QDThAm6MsVbkDJtWnMCS1fD5koP03Ix/L+d6GLfgThMY9tNAAtmJe0aXew79lGKQUKSvYCqbhM65
V1nAC9+SoM5KReJpHKR47geGfmbzo0XrxbuYsTpfm1QthBgfgxfN7TZM5963V7aQEXNjAzvsz3CR
ozC20+CLBO+jpG4Rp7xHcM5sfZuR/izKI0KK7IXwWG9xCLM76tDpDvCYo/K5kh+54NUebtrwembi
icFOSIxuuVvt0FjOSfpxIVOisiBgwgqShAus+lzZN6SL0Kb8CFHcrr4Ujg2gz4X6iCG+IXfH0Cri
j3ZhaFeXDZAAUxICsts/ylu34qU5GY5WoVFuegVYoekWBiKOkQHZXPtSxnfHPjmYvPTypQz+zE8I
O+HYJP+vu/RY9R9eiG1JO/wVcrTnJ+EnJp8d09Ox1JwKfyyijm96sxHDTeiw2gQBNtE/KfwVoDDp
eFHLB+r0EekTIKqg5C0o0Fokk8BZn/1/DRKYuUCe6u+Kr63b1EKqV1cYSQ0mnZ5EzVRazncreqpb
Bbwrrah1AvPIWCK4VralHIKmx3c/yvsPOce4PuRWuxe2PYHkLAc4mgBQrMexN/7o1W2GAwNh9sVk
lWirZ4Os52xLH/yGCdc4Sj7GGIa/yZDbWWbS2Eqr1sPDMvun+CuENNjio2uGTfUf2Ysy42rI9SAm
X+RTtJwXz5jcKvafWbJAwAvj0zSGJuNBGnsWd2Yg5h3Hc6yqD107kIGx4hmeZao5ZHqGGQZAnSfS
RE4OysLIauYklZFZfDXtfZvnT7VZJAmlUHDv13jqghca6i1lOcOt8mE4Jy9aZNCcp9eaqcJtmJP6
PKiP8JO8G51j3ZNo0i03bFs/gQOGNVzGb/qoRIVgImbe32KEbO1IoQlsPZsBw4fMsCUvT/PpmmHO
8h9kzIicpQ3W85BAoT38S4FohuxlhtKM7IGMZQD3nPWSsimFYEqg5g6VCx94sLe7+eBNvMY4Wjn0
dyCaGIs+ys8N+3WFa+C4GNkDtQZqrSWbEoYtGR3SaugbCTO3g2mE8QRp/RvbMFBFqcswzpUcTi5u
SIGp4hl0hVNjkWiJh/9hhqVx5SATijjv57MkAEEdGhvW5Pr+pCkNkUcvzNu3w9cjwAn+4buPwxHb
PVY2jy1O0cq8c1LrRxCrcAzUbPDerz4AbupsFVpw0zC/kv42oPuT5d9iky6Q3TuOGKZdeAghW/as
ddd36pZOYk8CvneVaCLEKjahJPGCFAzbHFPVItOJFFYHzvTaas+jGJvxDVTi+GJ6FE3ppiQSXB2E
zQ9jSpQuNlJyktl10MLll3js+iW2jAVngobb7sGKGs6hO8spTWVivU5OFAYMpukSFUejO02CMfL6
ewRLEim1rzOT7DrrxETnd1ncpXlSAkgDe2Pce6vqDyOumhdjvfK7g/Pedve/f2BTPG3VPa90XFi8
aYeOcYGjIK+8hMBZB+qK+l4JvWDpuGJsmd7BOya9UQp2Ue5lzXb/8QvgQmcpCWtuQOTTd7snHEFo
Z0Gpw0cwURMi22L9jgUI0wTe//yNoWk1ztQFLQ3uFk47PofVsceydhPUyCo8NaCWcY4NX47xqCT1
FBUfr1FEo3VqzTZnQcNErEZzRWgth1FCUxqtaNdQuHfstXZJfgs1bO6qXernfNvemnZQAfJb5ZhW
yr8pCZBbvbNkt+WoZvVrNMT5Lkw6Hr8Ua0HiaRDeK1MyL+3dDXuF3NN4/+kRAqQ84GDpAcK6pyRc
csMMrAqpfuvqWJTm255KyAmVTmyAmKRfOD2z5e95S5PJ/6HBTfF8JdVn4Q/t4ECH80MKKF8ccqVl
4/g5lN4/UG1Dv3L5PnCzrXyP7NFsOihuzs5va0001t+8hjz1yYCsEG57aCReB8kozyMndgXwJrsA
dReWQgr8uUBJVOnaauQcLdn2Hy4PHd236T/22R/pfu/SR3pguv6/qCl65chO0IZaKKtxqEKTl8Sj
zos5IhmbedAPN686cQBrvfeLMng1LdUn4GbBs4AG08py3/2tksBVtQUeHRyL8tYXlpP86GRr04+K
+/LD/2twDysoPOtum9RV14Znuc6CP712TBRAQsjmJqBPb/XXh7iyIIL6upf0nT/VCt54rYpjGfvk
1xjTRsB+z0DE4RP/peVA4zEdqBIddR8H3+8CvIK0H96ldMp2BDZ6ujALMFc1xir0OjkzQCawxxjK
31XEwluSSb53FY2SwtXe7CIoIQiYkRbm9+80pdJbMt9NKgMS0t5ts9ypnBI8MJC5P7ckSAjDp0x5
2E60SSamWNniZsRzWHpDWb3gplWmNLyhncOlWSNePciqRCd7bVEmaxS35Moeeqjo/iENDaRkxOBx
ZyabKxD30uVfbEG+LvCTjeeWNTCXQsN2aQMldbPLxS4U+gCtyO+zg2zmDlrH88UcylzIrw56Vl1B
YnlA5zuoATKhhFyAlL8oWlSTW3Pf0pVCX8aZZYt57hK6iRYdHEFRAJ9eNuAQmj0eLEEz5B8IjWys
tqdaKGlTplauY2UB80hxIedGOl/0zC6BmMOiFm6h69e2d0jCm6NzRaoSNYmVs+KSAWqzVTdpNgS0
xqvUHWf5lNI5HHUAXnfi7np3XIQxtCZv8aYm9NuCCYNRNqbrVDioI6g0TtCGc46DJmpRWpAozjB9
wT/qT4KzJbaNlKX6VW4NxuMaLAId5cxOgYxrZVYgzAEQ2ECGWxXuRLpxGc6Iathgnu98KhawCfyd
XYM++skiTp4kC/xTHegdBNR9yIbwV5wSMyCiAN5uuW9gYNLZFAv71R+fKU+IgMX82jRazHXZ+j8l
JGqLCmTUGNus8ChFEOz/H/1XG/lHWmIK6L/TMhsl/L/YFfRaYDou85mJQ1c4vBDd1ulgW4UKQQJ9
gxSOJREUAmdNCiN9Dnui0thldzaD+cQHh6EzcomUaRGYI+8hPh/v9PABCsTNHhWqO8UhlsWRedmc
UCqJeJwX9lqqVT+rFYESjTHxfSIULhBFw/nTtOde+pBOLgtzMfhfuUDreEPEIu46PjkxKqYsIr/E
dOF+stI4lo3GwYi+amBLbnRulEUgb75CX7+bkF9ziWOeQBFpGRgTue18gwp7kQPaEBFVEsqdH5zh
buMxnv12AtvFrS28qDM94npha9RSLV6R7VByeVTDxa8mYp9VBL13pmJoVXui0cDdi/ykyhU9b+N3
5CzjJojmo5HRROI6mumbG0PyvbWy5m+vVlrxDLUe0HZmEWbxOxgHXRjPFlvEKzVRBvhWkn+jgpCk
ZFd07x/CVwL3BcHeCcl9+aoY+T+m+vNzONRNb+FfDF4Ezcx5gXDiQ8wVfm9SEIRTTAfF4k9R7B+D
seO+K4CDkmpUQCd6e4WSdmymLYd08G4Wp3E0X+UiZNjoSgFN5564c0LIWIkUE6gnqO7g5L7RvUgb
fdGe8I167SN14jwekzgXQGXjU0XSCibesvrNXmSbgBobtP4ZRvykpdf1cHabGIMdeHSvQkrWhNNo
iLqOKYH7KufwSFggC5gMeaT9y87QJfFZyAipsrVmJUhyRqHA0EBuJEnIYEOU0u6NZoydIzU33+ZK
wbrI762A0kNktss8f4KvMpHdQo0v0PbeoCXkK8CCKTnr8a9x8G2pKmo+Q3eQpMvjRdXLOC1VN+QY
hd+xTFchNu3bIDUPBLhQfMfjhz4gM/qIUQxM4BluBzdjasNLCXBXl6Le07kOla2aNIIs9mUDVP6Q
pSrzPqKbA9+BN0Rvx3NjUOFaGd9L2pJ1o+QLbaey0CtmI2RWN115h+ElpOsLGvqpoqSHRhJarDJ6
Pvlgy+Xx0DNSIo6esot4xm9cFSUTNR2b1lMtgbxaIqPCAW2g320GPboYoa/WdFOez3FkvpgxVzNx
6MueGiRbOwfGMwllBdGuf6W4o7159jgiNUiek9F8bJakX8tTFk7f0DdwprDx9YQ+1ahR7PRTMOHX
rWMalKjWP/eSkOb0ojvFqgZG5POZiLw56V05h5pn5jip42hwgyBNDr2JiV82q+xzgRCsIwvmLS+e
CVXpI2BYhvzRNdzODYNqtCjpDLVOacysXxxSk7NAG+5pcovVChvUNfA4BFDJfmSyLxV6MXfDJr2G
fQTGRaj83a2PyrZDo0aahQbw4Ak8r0HGm+4P/4TUTEnxYfFzePajXzmTfL2+0FVSfkFf3aXsdZZQ
btmi14IbaIITwBFi1y1g/Jla6oleyQR+VNx4hAotMh+r3nlEUsupR5cc6PmjToyrjQZ1AccgsSGi
vA9JqPM5dM8yVzuRrtSBcR5+gSHc4Z/VQrrZChrzWs+tjGe0aFPmIsrNLLiQc6LU+VO1dp1Dcdyo
Jrxas+p8yB+s51m/g45p9Uavv603O8DwcCbEGQYud0CQHS59vVDO6Cup817EqNX87JetVZxKanOp
EsnMWAg87DPlQgRbAoOk5PQcat2dxj6lta79TnEa6SrFSaJBKoF5JdJsBqtymIl0xjd3ac0J/qtD
hp19UKODkqiywSbHee/+xKlwDlhYJyHtpAPy3CsVU2OJgISb+Yo2cDtS0jP+tNkdTZSMJXPm8RJ9
GHgxB5gQdy8Az2VkHb2frVEfJTD0/PTYQnUUeYDbkrZwPYQ465rUSY0upNboXsbzuV3K7zoQJoDA
x7nTKBzh5AygG0wAhh9NjKiHFhu6EuT7gVUnMGi82rVMCkIE9RXLAtVSvE28N/qKCnIRscFGB1BZ
FgB+sv9Fp8VI8bjQ4byw3YfEgwRRYdSuSNP3O0jIVsm2s6LfH2ULXynjhphynouw50S9AfF2vBSj
1MuWxMXwX4mxz57c2FEjdKDLogwhsKufWJugiXb3zpcjKwPebkcp6awLHP3N12xQhDXxxU/lbrIX
YOAnInp1+L5qBW0OF/Yo1N4Hee022RdgOYzzDnHDPsJ4IsApcU9RRKlbGMC2sZwo8RriDELOjznG
MTtmjV0ZRjeMPGqhFLlOYE7ojuHo3K0h+Q34z87W0pMENL/pWem/SD00JEZUsSRdpG3Shczvwe0Y
p3OLJ7Y4iQegBUtKt88B5DzpbqohRYNYEyA1AiWRzBNwKb8vhG5W7TOskiHhjIpny3xLW0fC7ush
tfrATGdQbvcaLvRLqBYNFNq2BM8eogVCUujkyGQ7Sl+XeN7WaHq1cNzqyzQun43jsBWSVlWxaulm
HB0z5AXqBAKBAj0K8JbMtPaGwgml/srB1ztMwA1O4WJTmOGsckEtKyMuK+XUwcVdtoEFLi7gZNKH
n15FX3xKtjfwasuZElwjeC+MB5FLmzuUPHyo3PQk2oHR+ZrcapRmG2Xaw4YLYuoj57c8wtT4D/45
a66FkC/IthYtFTMVe4gZaqg3xyirzlDwM/m16CGiRto9hG/IEfsuj2P1SD+MJJkVARZ0Er20kVR4
W62O9k4aqCmPvWAGu5faZY0V4xTB8D5Knon4mvLrr2SxBNjwsIbsQxulwL7znbPDXBgJJpKxO/0R
fmJWD9D/4wFt0ZZzhKf1bvaOIMSdQLQ9CX04zmt9gv+KGOveFfK85Tyy6HFlWemSnJueKkKerFad
Lo7ca7F3RLx/LcdfKT7iRFT0jU/wKxK22kADFtoq9oZO2Lsokt1mSogFPg/QMQLSif76E+G7TgvA
nhN+xXQ76K80OVEwKaNql5I8dbQ4c4ge02ORSoZS71e+Ktage5kMLsO3qkTLbOnYL4J1oDMUTmFy
T4SlhcwxKz/Cf9og08MwH6/0hqJHfc6wikodjT64bYn8oJ6YKWcNPqIkXim+hIkr5xjMK9T5pxNp
v20nYiLzVmFgcxmdR39AcqcyqaSc10eMbWrZbR9xGoJY5CEjM2jl0V4DNpbzeFE1U5CjDq/nUbie
5sf2QN4iY9OjepCvm3fzRbDebIg8+SgxES/FRCSPJ4f7hqA2ZpbchpVXB6I+s219t5xsEi9V1Sjl
zUmh1EQMFI7VoS0xex6HoEbkYhLnwcXWUa25LlLIx1UKyRu0f0rMBpkSL9OQ0bqSRuuphv3gEROW
Xi+e+SO/akdEIqZE3b+Zsw6hdK/aGzsY5UiVBl0CoZhQ97HHlgf4hPfTTgnSQzSEUAsjNZrvQlxC
N1Pv85LrsA4HOMsvc9Tmaxi/FtpN3iPuwiPwXFLxFmnkrXu1h+jvRXAXEQcmXuoCxrNAKLfSaf+F
nnp8FQEK5nCMci8qySKLhj/xB1eCruAq/3TDlbyrqc7ypH65bsr98NYgj6gXB8zoHuvDh96XziSe
eXVO/OBx3gnklg1lu46lST1KVQwofxWTj++5i33zVWCSrLMmkGmDBnFpzBHCXQlHULVqNnUyV6lB
Q2AXYisRN82ufbHzEFXnBJTV8ZN3T/PJJDdjqlFFYdSTt5Wcv4Afm0EtS3imleSNqwR3Bo2/wlTG
c7fw4LLJGYC/EcD5jceXtiFKyvXjywCoM1KfnXELs/TIVy7vwAc6l8rRgGIc/+X+SC88q7JF5u+l
cgQiRIQD6vFKJKmisoXt8EBOh1K5xv0TUQ5QROoGgGHTUli8QxhXFD6k3ftjOWx9Tj+mxZ9k/t2l
VIdLIchNwd6G4F7zPkR8qLMjOF/MLJQvR8Hy4nDktFHRDzF4qkw0ozdyqnAg5dJxjHdk3tkRiyNb
EpLw26l1qiGaGaAZ7g8kxpFHpbJwJPl/ZI3UaipajoDQidqcy5u3eQNYr2LDwIJb9vbCLPt+EslC
pneuUGUTuqVW7hjTPHRO4zfoTfkGxcZRPANfWA7l6+B4HLTpGR72O4Sq9zjL861JdFzVnVyDqMeI
BhRJo/jknjCOYf58uCmcUZ7JEqfrSTu27tY/AYdOie+XP+Bh21H+0J4dv/YAvP4Xelve363s260G
MQL2v6sIgHmImyzIbv4iBIUahQqvxPxFGp4IOzmgqVEcFIJ4hlAEASBxHZn4h9SOIpTAt0sdVRME
cAGb4oa0dACFpBiFUHyePrOiRN50+yNDginRC/ImIPiFURHJ99Hy7s54Xyju4HNEE0O44kYLnHWx
oPesSmEMElXU2hRLpl8jR4eJkAAb4cFCLaDfQjxvLjG2JcX+2hpegJsCr5jSE8KIzr9HER7Vpnsm
fN7XUhWs0m8G+LVZrf22Ujc2zvUc+8qePlgB7zmoTPPENUoAZgfwQh0ZxBZC2Ew2dXGoXZJtsYqw
79rpP10hYGCjQ5j0vY+1kVCLCil3cd4/EwlZa32Yxp7xn4+4HK12YWgRKM2pu86++2kvAwRQsU9F
eSd8oNl4hRckdPMt+LMmC6lICsRgP4P7A29W121f+37cUNxYhvQ474xDCJYOd9KWSYN9P2AZ7CRZ
yZ9DBg//6bDfKWAByE7sX8gpRj39kqNJT4HFyVOKt5Eo4mIm2ubGkWxvDv80RsDNfKHxkGfFYnvv
6uHca8lbJtAPkHALXkybLK44D01mGMf8OygpHPLiVrZknAg9Y4ad1S+bdXGsgJAiFPL42HoQ/3rr
ox+5TuP/V6v4xO6qO7fet0yEDGQ2xpMfXOAHwxTlCWIzY+5J6Db5bgh0QhwEzbVySQySwRAb2Kdh
izXG6JaHbaBXFHP48mJYd0Xozq9DgEwUyXx+iW65g+gpnCu9SLbiVtQo4WV4zHnySn2woQy5GMJv
9ifEkJtVeJUnH/ugwtIpe77Smc1Cwz9f214ax8xZwORhIIy/8VDa6yuLpHdmA/14PmLitDw5vCOL
4wJQXZZIo6L6HE6wz6DzdbrmdDj/4H7ZhBE0MYut7tpvF95oEFmWE9I1RIw70GUzeaCbsG/UoMoe
ZJJovESOkXhLDiNTePjJGRG0CQxkvmxvSmQcGhw5Sphi5knZmpixi3SF3SkS2Ueubs5qSlJJcgdm
3oorKiwM3TiNAzpdEUDaiqVSVUpDwjZbRsWPYzaE2usKla7ojpYJVnfp4vI5SufXxDx3l9mEqQN5
TV05ATBKlEV5MVVGayJDFfxmTf1n5g2PuZFVYw72dAmqG7q6q7xKqoIu68/o6VMO7oxJ0HsZO5b5
2Vb1RQa02iVQGk+cEGxYv9jrIbO3kV+/EGhVgy49f16fKLoZF5nPuDXICSc9QMLT8guoRFS5swCf
wCtq3yn7SbqVqSiV/XpKfnB3sMTrINXB/v8HqOQBNevMVaKa0TShS3Ha8cAgougHYC2fX/aA0MOK
wjPPNnwIMWvfCRSCcRoeZeOqdyAIgg6D+sQQwz/1g+olhIsPvBo3KQ6GHxftSDG1WjF4m8avJWq4
CpqyspCN0iaed6m4TNtNZZzVBHsIskSV1xdA9aUoLNwe60j3XLmyU18bxekSDROxOdJ+uDPVffyr
4apyp3THyTe4umbWSXFE9T6i5uD3bcfI0/MHZKRA4Jhvq5sNDobDCAMTwXP+MghRSS2EyiXfRbMV
LsiDiDmnbzDU3vfZRhbXpYEnKvrOQk2fSesoNti36w602QCO15IqWjt28Z3C20KnSmBQ1dp4UyEu
URGSg35hKxFzYahth8wVTpz+kaSOdmIfDVz6FFwQAy4W//3ldgpS5iBaQUcP4VMDiWm6/iWCbbOG
G31SnTV+lfioII0VfUt6hFVSzcCYufjj/uD+psbX4ae0PxhXX+tmKGBlGtxwGBbYN79zpj8Ti6Ck
sGatX2wfgz3UC1vOiPFhOB0kgNQoQUk8fuAo/nEdShOpoCaCrEnXE+syHQvUMtgdhv+tEWvLJjOZ
XlJrWbBW2a6St8ynN3mm/S6/5FCWzLdOQZ8kw/p//nf7Y+SopUbFXvSPTrjiX/p9mx2V0bLOkP4M
/NwrRSTOIYacsl5akiOo1p03J6Ue3xRMyrD1CdvwawEVpzG/1kj6a6uLgezLGTAj6Qgssys+eDeV
e0Dm0uxLjZN3yH8QZiDLykH1h+ssLT/Ov4G2Mm4pye7tkvq9Br/ZPuUkt/oqXT5G2A0wEMP9zRmY
oIYdCIqHpUIJrftC24RXWCNlCUiqddzXPOcaE/VzXEo43kDsXh7tpJi4tLkQ1yLxFTTKdWO/4cd3
ylrfqVotVKa8k3rWN1X1VUpKETusaiJ0OnoDRAkr9qdsnELZZz6iKZJKGsAbXK/mhWue8GRmHElJ
k2AHOTG2WptMeSiQDKFDooe+aWD37L/unyoBjQZyxJP3UanInw0DisHBfEQcT3ik5s+y53CTvU3p
q5zzeyerxY/giu3J1XjDu+lVgcBrx9XVtDf2dvfRZTrMSJu71d8EPZL0Irtz9+sUMVQxf/YcLT+0
+3cG8FHVEL56lK7b+H7e706+ylFXHHPv1zyYAOtRDDwAgvNrrGj+4TAxaiGd/kfeViKPa83hhnvQ
8rj4aEWyPOkxyZmhyhDb7RuxXFsiISQKRa9DRwVznRGz9I63VsiXlsGOMw5Q59LcZJo2pAOJCXRe
e0pdbO1egtKrxFFXLn7lxWAbpFC2ZNIf3w4pBy5YXXz8OkvUDaTigOqdAj3vz8rACiW6ubOkOoX9
X1YnNU9+M02gEy5ILP58tEjcIzd0fE1Ki885OZCLy0qcfDIP5Mi6RYmWnu5rePyW4GcSWwfxflXq
imM+CW42jxyqxMPXrvwwQZPQnEuG8dPtJz4d+D8bBpPi246HNK/LMfa3hkUar99iALW4zI+t00Qq
DpsfgX+ReQBqFHdW5AflQJW8YU1lO2vYoD9fZNmrmGypDoFLYsPbwX44uIrX8NCTrq+O2m3m6re/
jgzpjQmY2byOCGiMXvDD04M+zBSYgipPzJHUYxHbaXKqYlmgJYGMY6WLSxAO8IxohFaIV4QrYGzD
9jE6e6sMGJR1qe89CMlQfHikGJN7Lu/SCVMbvbmByVgWb+qreG2QYtk1yPrA8VaIWxVpvo4mJf4e
Q2j+JYFQ1MccR2MN1TezF4wY2nmnawfFboBSw3UwSDjjASpX+tgCtW3l4HMQYQ5RtuXpzPfBiDCZ
w2EgEwhmC5c76m7+5KK5sRTtaWiNf1ZiL6LYM/No8u6B3t3LmMIh+p5yeZJ0InPSmduVsgZDiBpn
BZEZQy9MER0BOQI9Rgc2TwsnRGpqfjz08HpStKvtsfXzjkZn+GdJ6RiUyIXsZZKUFyESRujG+gOA
4KXYBopf6Td3W/hN1drHLKg3WdyHdMJpdhFWikyXrOApXVAbzvAajoK4CBqOZuWypMlXgjeyAlwB
SJmqDd4TPK0MDozJSqT/cUaXzvq68seGusvQqK8J4GDl0nuwHejOw0nCJ3hK+un/6Fd0/WwChQgR
7Pg6PzfCdTeIK6SusLs1fqp5nLA6h6Gq6t/bXtSp53EnXIt3dzRaXiKX51Uv0y9OYv9oMyzk0keM
bW3KkxHIvmx0cFdvPLkS1CUQ7beqUw9ZZ8NtCh3tZnmm21U+lBTar070Y2vvYkSDm+C78L3P2f/5
PpbZG8xLAFq3V/kJS+i3R9ivdsdDHMptY2zFg3n5CgoeWjzuiJfJBb5bgKjXkMHhIw3gsGadxUmV
aYQfKSy/09TIfWPxscuVN5YGuTSElmu5F7Kibw44p9nAczlktX49G+7AC9kZ3MXUDWNn4maTj8z9
wlasAP7UaugFUze9FXRbdO+YSoRxL4xLXeaLIEwfsKnYj/VL1PsFj2UNji2urGvBFjDPx09/FZ7m
5raFlXwU9joM9PEAVDsRy01mk0aTEGIR8VHzhYRV0VsaVYL8epK5mP1w+K+N8PbmDy0kPqdGtKnr
WQeAN4y+oYy6le3YmsyRpz/iL56ITwdCUaUvU+m1tKozbJrq4aIYgPL4jHAjP7Qm4+Dpek5TPsVU
Jyf+y6U52ynAhhGt1pOEoyw9sL9JMes9DlYLeYAO7D2IlXg6OHuIsJEgyA/CxBTGwHvKQyqb10YW
lIRmuOPI+peGkdLDzOhGV+C6V+bsIOQeotegXajT0PQ0fZb0OAPUu1NuD0+b4eZtuIgnTzOTY/NR
CRsYLxso1pwORqwReWHG7HlChp2tkMdMJSA8GJP0rKpBCfwwI99PuE3KkN0tbfNk5PuAWX1RyyNe
LB67NIAM24ThESHsuUXc64B+OwUM78/4FQ4J2DsA6SIAs0IrcOkXJ1xv7kaCJSO4OR/7eYyWcQ4l
cu0THUE4Yc8T4bT2cLXmSi2HXn8odKu9RyOkfyYAjq+Z/ILvVSyMDh+yLhM5PqvOQpGZB2lt1DdV
jiSjA/wOQMb+vcpop3Hs4OZiTWuYU77R+bwi+R5oBfwiljWilXErJpMTKo/IphH58hEoYgMr0jo1
lJ+QH8ErGkD7AOIKpZW2O+hB98lTWcO/DInwzMNhGBaeJzBNCQ2EjPJAqSTMF6RkvoYFoK06j2ad
LUCtSf8UL7QpwXcJJbE2P3o0salhn0kV0h+n7ZPzFfedfVkekp1XJ54iTrDZ5SIkfalPE5nDLVSL
/FU4QOUcUKjfR8eHMEnFpTGFpiRmdvf/v8t760OdSZILEGShUtlxE/4spROh2JHru8xpNmVl3Cuf
pmf1pZ3uuKjcxWpEGiZ5xfhLVhyAlZEK8JWr10xuQMEOu0dcemato2mNibWnd19VHnUXse1eXabs
vtiE+bbMrFH/LdvxL1UuCcnQvmYG9+XjLlUVnswBYXaK0L7djPYt/p4PsjUs7R1thoVvpOQuIPJ/
QKuk9ZZ9fMKvsP4TioINwxSMnbDEbel7xXJvP3uU7nRpjPSbRuaKupNViMQ9Qw2Q0noXTnqabiCk
+b11ERelwkX1hSvFLj5fQvBGdBVOkVZDzsYIDkYNWFreQ15xhVlmY5d20Rg4wlSuudB+Bnwlkkxl
voPtQxa+czABTBhs/5goo1+S10YnaTsCsL834cyybSbYeAOPAlLNDbaoNbaRfmKlCpaONqioFqTB
8M/14U/OCiQogHtVYf2lfRv5CCkhaY3fV1sJORl01qcmtFH+MaDrFUGFFUTa61+ynRINsTQIC7tq
uoLl3zCAmsJFHK0px1qzZ7usO/0yhEDoz26ylVHsRSIOrpnYdCFhKfviDY/pZsvw3FoR48jJ2QUR
6/boUK9RYvFyFhe8zxXvSLkqZa26wWW28VBb7dLBagHz19SsbBGpGL6EStLSxVHninKNRqJcb+Ch
85eyQg7ShYqzgz6hCeVmPEEv82CdD8qzTc1WJlvuXJsGc/3aaDNRIdp3YsS2RO6oQD3vXtjMVYKy
DdhsMQRNlTEh+YCGWeV1ca38a2FuP72FX+azNGmDD6teC+fTYUc4vJCaxPi6wPKbF5G2hc0E8xUz
mVG89MG92GxFzdrVJLbQdseUCX/sys8kUWk27cJMF6I+PmwVDS+JlJGALJu0LFJQx59Y/Oa2BCfo
YTfnRtne0vxModFNxaQ9nl1w7wKrF2hNpcjUoD3krem/2hPfhZk3ivWQY7eWl/Ecf63AAGxowxvY
nYiSD7wjJ1RktnVHqKmgV4+3bD/p0fLz36DMQ/iZkYQHrrBj22C+XrzlXxHgmmiyFF100cBha0kK
1YZWEBGbqlkODchoYjG9swiRCl0z8wCbmZ5Ms4XBSeErbwsP8ytTCxnfNuTh3r0B2Q8CDENYWzya
J87ufbNAxTXdGvnBiVPsuw+BkHapqCnE5O6bTkTwlzGQeK40jpdXZqJzVthxHzADEbTFHw3v90So
Ts/kINJ0nZUzdlzoBnDYHJl+tKLZ5nsozgXL67ZDl+N4EbsgSimHE2kfXQCfBoQKlzcho5fWOYpl
Md+3J6JO9s3j19PZiN/XfuNA44/ZNs3kSSnCQdocd5Jx9v6cyMDBp88vujDDRM8T1fdArHbDu0k2
o0y1uJ6hp/EYXlW0YCJLDVRO6C8nwl4w7atNkQsFquAAnDEycSVf+4SvGBg/uKTcPvVRr2HzHaJd
F78nlL66HtoubyXfax9tVGZupH+u8829sGHcKA+PzF5nDvMGReEnzFdfGPbxizOFqoCWVS0gQQlP
ERfWQp/oAxU49D00OfrgrQXN2gqzc2xg7qMvLKpqrhB+qHfy3oPG2OmkUYLlKK3tgBPwfCJYZUcU
UHA+uDfN5Yn0uMtRbb/Usay05jsaucsMSCtA/V1sTrBKDucOGeIpqE91AEHdIEs2WjDdN2kL/+F+
vBCtV7zarFXbic3iIQaKyN281R2HBRPN625+vbiQYCOaaPAi3jNvWipJ/m3da5P/mRkZFKo1RId/
y+baN5d1eitMwyIt+ILnmWn5GPjFgt87qAXP3XjOzGc0U7j/Ij9LkdEAvaxoaXG3ozXWt3ItySnI
qM/j7bzKWZrulXUfGSLipg5RCmuWHpBH0Xxqld4lUi0hQgVSJyxgy8W49bXDRjsy+yjxvQiXFyZT
fsFN/ZbPKW+4ATSWHVZWlARurs1/mBkD/LtAbc8F6vdunn3cMftjuPxu4JzmveHkYvRe7VcoPRbG
7PVkRmMts07EymtBxM5HJCnhh5D/lG2XlzQ4jxvnmEtFzvM9Z27cKZfr0tScgKr2O+zBehxgDB1p
GwaEjkcYqHGkARGIZ4+CrXf1SSQny1L5Zsmkf5lK596XHCm+LUdLFwTVq8pDkEYgCEqyjQGl53dE
YxD+loaLZW14BPjl9j8HFtieOm+aaArN2XyLCIa8c/UPDRDdQrktzwzZq23qtGZ1f8Lr/gKq7p5X
wA4SQOwzeBzCmnj5VbAREG+yS7H4pjfsvzcrxFLXryNie3LjbRIcXBDEZThHIktCatSpzHHvAm9G
M9HxuSbBJy/dP4bJozuPe2m3G0Vh1AoMA1+wTPWGf7xwC9YxhH0qcCmJiCRsDS9/uklW3vdfjP71
sMQozlOOVI6g7/z5FEPi/k1Pp17ETpl2NYhjGC+tXP/zZQb9pHw+Fq1V9Xz3I94zrWA5rvUt4lok
M+alUFx7wcSrCs85J6Nm9K4qFH9ne5RvJhXlV9YMAQMwQ9EbkRGbDBKQFgMX9CCcm3B2S/W5f2Bo
LtKMnKYEs45kYOWKKbFF/5PYsCwwcn65tbUQeyWqbCl2h7nosb2XQDDC07KVS+/cwn+HD3hu2FI/
ryG2x3AbRhL3+bI5n8yGJ6p9xmy5gUpSUKR3dU2hM8n+g0Z33ZnC0wIEYNw299VDGeFT0xqQ113V
9+YTDOiYuABwHWGlQxpW1nOluhbSQJlgI7fut2nXNoVoe5V9Gafb9rjddpdHjTeYmCrnUOzI6PBl
gL12Vco6Y6Pe3+ahOgiI5xX16VvRC5RttDqvpJtgOS/fm0r/72oy/l4SwN+HMknD0C88fTJzAdQH
3oZAfNXr2/AJfzT1saCRAndYgvkdg2nhB8H3J+QyKIX/c2DUTPPMjGALgjR/BfWE9ghf2UoidPib
uvNwPvp1B7ef+5CuIM/18h1DUskwvMxuSWrs9Gg4xYQjr/8CbkYrhkd0N4+TD/w3eiKzytOJIysL
aFbBWIyIh/B+40/+xVHmuXVRkY5c4h+2WwwYut4mBHebTiPQxTKTRcD2HjiRi5vUDL8BQnWTUa/H
h6oYaGgejt1ypw4GDHkw9N5hL7ZenTFDKmH4LssPl94OBcUICQDr3KqAhg38qnml27vnXEIV4Iqq
t2Nyo3Iz9o6Q6XdUVykW1I4nA006l2s6kqd5BH7G2jk4rjagzcj1hVxHXD+e1I/Cjogpu7Rf4vU5
8Gvd0PIKnNCRyI6CgyvsXMrtQXFSLfiY/93N5xZq4zmBWApTuP/NmBHxcVUD0M51Tl+PnaEUCPij
A+V5kI7FC4Y+Fm71jERRTtm+8xNd8S+zHZAkJ6v34Z4wbmxefeK1zwLlE1wiKGAoe4PD7tEBwC2/
TBABX2jti9lpLgqPCVXBi1QyDdZVXn300ZjXl7q2AP0/BQmeyuGabt9Df2StFMT9LMgI2rA92zRa
jx+FZuV2JnKFMj8v+PrN+glE6wtdJvWg5J/URvWNvaNAO+4VEmEzaMD+HCOOhMkNDSdGLwGExY5h
3bRymkD0aarlMkWOm9pfjyto/O/5kBqGx/KdFzUkBSlOylWBI6dEuxDoY1YViXf1v/2WHV9NBpvZ
fN4b8lc0PJHdCojKhHVetuGxLQebhsxZ1XtSS9tS+gbfhJOT90zDjDMhk8Pg5OOjosoP6RGOkHFH
HkuJwK1kmAj+xGotFz9O6cgQGfbH4C46QP8smFkINvFo7u11HGnGHowDo4AolRNQEC5Iy9gcqjE5
hC8S2yMuzF88NtvsT8/djqe6kEENsRxcby2i7aF4abWSQYvVaVXhsM/OCicypjmk4OpKjlcovYAl
1j8Fle7XeBxrKsDu/GX0sN4Jt17+Hlfxep4fblolk9rEW75A7FoY6N15VlLpRZhq30cnjXgHXy9V
p/aae9xpuCk7TIJp4DzVCp5sL7qef0VnBQVb19SRPFinv1YewpdVrL2/ZDgEayoklzfbvhCNXTu9
BrCXjfWES8lSr7c0FcAej9RVx5eyTYFSYGuEC3Oxgdm9M75kAudFEP6edLgeDH7nVsczWtv3CLFd
T8Kj5523j/do3jXs271KQ1Ep8c+SrN0rnWWQDzg/jXlErLRX3MYsfxz+xDJlNyDbjWy07EzS2j8F
qY5skSsiLSXSKlC0h5C8+8Kwxkd4Md5ex/c09LdnqasMp++SRgJt6Izaqese9O4hb1lxmXxl3PoL
MYUZ4lA6OKQHacvBX+HzZ3Mwqh05M4Pi5kf0yMiHAGvH66TNGtWtSM5iNRWq28EP28AzPnS4V0xt
ztv9XngmsB4+vwkl8wVUadsWjMmjAJ0XDXvfsEews4Kcs34KVwNHXfGrwnQh48qLS5JQRttd5lSl
1+WY0kmkGODYSvys3JgwYFuWES1Zd3CHg5e/FiYcpxcaMrbo3A5jnJpqzzLmfIxV9TnOcqCPjqWv
tHkRCiKnWPqw4tONt/cTDgA586yG6w8RT13sAjklu9kwxhsd1csYPXxYP4J2yVpbgC0OtAsWmjId
27ldGgGzXqnghoyOzRjbV4gpXJbzoWa8a3qQX+n4HQ8dPA6mtwRSBWLyVwt4XkOkr91dudFgJ7/e
CVY3TO/jVWZc4yEEPhWqDoVZU9k/iqcjy+ycuLPM9bcAxtLGp82PZAtYynBkGOMMzJ1ArDXrJNXl
/Xd1vqRpD0vUWyHlhigraVHyoDokIpAT5+rP0vRsP3DqqRoLjMKbUSuPrAqIeL17sf/7fnXtYqQ2
3ShuiHKnTekcm3aW4+m/bllvN0Kk+6bJbhXrfwkyRDxIo0bDTC9/BS3U+Y0g7NiQ0MIjyvw0u1BO
ZidCKcCjdoiIZnXl1q/LmIYUHsthsrY61wH306MCCoBp5emuTHa/O1NbnxhHa0vYsvF69nPDw5GQ
BhwbHaPgKCTQDmkrE0kAZyvCP9e8Oixi4LzOqyzwYJq7GVkye62qEJZAR3JhErugvaizgMuARk2O
CF/RTm8bNroVudHiDKf5rh8zolUC6/Ad+tSBL0zR4Sld6E93j9H84Fm1FIhwrTWGpxaUX/i01tnV
vNjqKrBY9d7//we6PJoDFhdsrWCqEXbyBtdb9xoy/RPzcjY43MsZ+X5NSUpE2DU7iqAex6wX3Byr
yxF79qVxRl6yXkmktEpJv29jIZzJ/uQWfstQRRNN0pdNB5xURiIEdKgR1v2BBoTRLgj1pOuvKNm7
VJXE9o8Ng6ZFEiSqq9EXKb4VWc6R/2ZWqHzhhGtrDLHs70YtCD6xtL5B177lrI75czSWh+npYFZ4
9lq5qr3EmSVpPalz4oTKqim8ir6GH+ZRXdMB1nVDdLgiAve4BGriWPg331Xg9GRLeFanbCjPTUNW
LNFwVU9xMVY8f2+mHHH4CKew/qj7KtbUU4P3r8yWgho4jy6vKIfZzux9qtAeopR63NVrS/K4qB1z
gSWB1idZbyqoFsKG8JX68HbgjExLLGHB8Zbb8rWIdfdSpxrMxl1sB5MDulGdhwowwrrwyzI8LVGQ
iQjyOSkDC/nwnD6AqgKtc67P+k0dm2uqMOUCAmyJ8mHKnAeIhuITSSbxlJ2+xTql9u/7r+fsL1kA
63IiJlsCZoYxaVboraLEkxVfkFeHqDi/IS1MlkQfiPYnc8Pgks06NW2a3vaK4uZH8JqWVfExY6mL
SB0MWW+T0zBj4FDUa2ocWw4J/m4RaKlK353IScYLkAW4isFXJKJK5xFDZE2eP3OBC04L6AyOSwJV
8n4ubtlzMQf2UtmL/U3nvWtow5Cm+P/3WlHRDXgfh6MxSgKBMXFAaqeatodBIoWD59bmstOQ1KlD
IewjVZa+lIUWLanW++4tnibCNg/vH35YKXHlvzsazKU9ImoWL/J7R+mtwvhrRNqSpI9mxuv2X0os
xx2xWO2Nqv5jZf5AU/X+artub6gnq1X9eCB8XaFwk46wRrCcumqKVPVGgDHkcRAvXufUKZx5sFD+
jISczcAFt73y31jR1I4T6iCVSDd/Lc6/HYE7vkN4F3/ES0fHRYK030Rh3STekictKs7MTlb6XWhb
R2u4b3iuSCOnTQ1K8iUDYCG28AwwRvhNFdp5EvHor0WwmC2z0oOR/ZvWFDJmVGXM1EcHlGLXvzsA
MO5E0KVTmW8EDOXHV+uXMMsEFW5SiGp2Qzt4dIcELkllImUJN2yEPTkIavNjG7ErpuFaY7wgk0uz
fMFKhyiKpK3bPT0bgQv3GqqdR7Ob4BbczfydgFcS7vOOjxw1o7G1O1NyL9icNCtAvjjS7F56Vos9
4On3HCcrtD7hcCIiMYcFbJgnOv5LPUmtaW+9lfAIN9U00CB/V+e8jJPD0e8qmowgmilkpnnSEee0
oOmnu104pGPJ5asPYIJ+iuNP2HqKeW7+7dPSQeWhLvKPtaNInnZ0PfudpZK+IP7g5SOkZI1plClE
u4vnnWsphzEV4rnFalp9ZA0iq+DWsbUDnzdSa1eGSR8CNwU/FzjElNmBkZ1+HGXu/METwaSvqPgH
MIzRLPAfYU5DYEnn1wrs6aKXXZx9bqFNKWH0eazgvQCbzDHnrOfBwomnuqCEmp/TRcjIZw9buW3X
E/0SeHTyz850bEaPDTMUNSPis41V/UdCerIvBnfqrmTj7788XEOJ1LwjpeIo+HcK7QLlSR+VK+Os
Sx0L5Rb7SC2CD25K6vbgrktMxxthqPYrR/ziAXTqe+y1cAi6T1KiuIIX6H67CBwibah4CVRhJXca
5Dn6ugCwotRRa54+9fCi2M0KgA5WCj11EsYDU3Isf0FrwI7NNSyCH3AIBVt/BtONzYaFEPH7PVzZ
fJQmlsdNbblGHelAUSQ3dXebG17UI028HPsndFGk540ji4EbwMubt3HLZeo+jnQ6QhMZKZsMxXyV
EEpuBrDgergubrrIWlpRncsSzEhGOOtgo5OGDx0N4HUHfDrJB2mCjgcwdpArreofgqCHXIh7tPjN
XSTRvEFIPnSyoJoOUHB5aKtS8Ypz5cow06C9MKZcwDWp1MDi6fd+I1esTYxIyDPOxt4h9c/cWfZf
g63AB3s9qcKSJ3nzP79hwr/6ij+uUF8Dy9HsJOzUCAq84AQ40yKMLU1RfFrX2mhm7BV3kwaPJVSl
KQlYDGehvVLWUU38+bljrDDd1dXkw9yZ4jGNcRE84Mo0Bkbb2g8ekomSNh5mEvN+gTH35nASBiFR
Trq0wNu0enYYnKP3DyqdUwa50owi9QdBdqerWlZ/txL/m2rADq9FfDLkb2sLrnNMY15tzNJhEm6a
2F4w3Kugnnw8lGSE7DLoCiTSw/t2EsqtbjlF5jEjCQTf10MfzHz+YzC9bzg815HpATCpFITST0qi
vqSFjHsEXOCR2CmOqDTgW2zN1zeMcLrCssuIdL2pezKrylTwvL5snLOlDcEoza9janU+ZPzmjaWW
eUjjmNFezdrkWmeFItQ8ELzOuUQnLyyybbA3k//PGbzD86GH4AqQtz2TD9UVLq90+dzB8k2Xsfqd
C+QJLZmlUrEmoOsFBlxUzt0tyz9tnvp1/g3ogGc5J4IIWVVLXR9eRAc/aQs43WeqKmKw1VBSEptS
KISUBqiCI3kZL7EFplgmgKOJJZKSvM+exOpjoLsgdeiomE5gu1CyXwo0xI9miM0hhsA0zEbTrB9U
fmLvl98Pu4UrDVFXsNiAisYfVrOa+YYNvp9+CalNWhjHH0gyTWFMhRNMmAmZFRUu3KtSnhw31ZeF
cAYqIwqNMs769h2xnv5lzLVDAZwpGYSUzhwyQT2YBxUCz1ZQZv31M0+Q9i5IZb9+ucTLQwugjDco
JQjxMv+lewosPH/CVmAcJ9q7pFnLNX+6xmjItF3wERRUO/J41h/BEowZDe7egCTCu7PZ9bttMNRt
444npXzFa+ePtdzjtsNtTR8/aeSBvdLtWDz0tR3zuHrt2C9sQiUXhvXERIYkqj41IhurxomecJYk
Opqk6w7BkAv52yj3MLyzpiDt+cfbq0GV97xNg1IxFnezbkNIm3pOTJ4f1iWjGeZzWqSxcouDWe2d
Z8OK7Ylto8SbBMdDIDz8I2J0DE/+0zo5chcAHV78YNQJPVPQQCTaFFLy2YKsReQK221zPwFMd/+i
fHRpyKanh+OMgZke9at/YrGt82ydL/rsZ54doXar5x6xyTjWqlK9slB1oI6cV1MdnJlpgihAFDXX
6ioZzOd7mzOtHyTZTM9A6NE+l2HjRCdmVGDeuYXVmqBu5yrn2LZ5C0eBGkllMox9x6kKM0EQvYO3
5M+9vxPibVaSDluHADIkkJaLgdsdObSJGwcLAyO1YUnNtlwbGBSy2AHO8A5noFdj2BMxDsTvFyvK
ItR99IOvYm1/Tx9IYGBekOmeynmbqNjRc7hESCRXcZgRYjd1eWGEffhDk08sF65ypzx8i9THwavG
uC++0Pif3TSuqhn8ubjEePQWF7ZWyM7DeF9KFEQq6Gpp5oQtrN/xBSAfvrFrMopb5Ah2rSW3v+2R
7JIc9WINI5OKevKS5DDWOcTdL360e9KioyEVgPz0QPe7pm7Rv3DCo8r9Gv0n/Rs04NTDl5y5HV5Y
8C9veKHEsbx1ual08k7Mp/lTShT1Q7JkeVWbgPj2XXBCxQDTRNlWCqjcEI93Hj38E0VZEhGFPhGy
0LyUfM2kJkUve00G3kVPQA96ttZYh8p+TxH2EiUEtpIxXjgUO/qn7sey5u42I97WpqVuI/Di21Jr
SSDYr4tNniFBnP5FFrBTxr/UXyU4TjRoSdDMcfrDjTuIzs63DzdHSuealtYq83lhEOuYMdVn9u62
V+5L4FCHXn5nZG9O8A1Mg4jCKINs2QtjTU5c5C36Nn6UmEGP3uu24IeisaHFZry0hbInI0QOxvxQ
Ees6srTzS5tHx0zZ8F2l/2pBh5qo+rrJ15rkUMc8fZ5JoxHh6/QGaaL/QjYDrssDJWh8KOvv1Zh9
fEh7UJMUNVb3qiBu5hQXbjr+d/7XFGjIpf65SjWXO97coS6n2x2miiyWXFVhX1RnscR/Om9q6Btd
wZIC3m+HA+XEA0yNV/kXRytI3QfmLpLqAkl0kchnN8TZ5vi5KTIY3L3uNBSuzm8cx6teIVz4nthP
ShAFtQUhA2hrml2IqVw6Nl6oh93yAj+FyJovmrjitLFEux5qi+dSKFBDgwHK0/FUAxv+BYR0b3mS
SmkhWdrXtBwe6Yd/oUlBxfzXl1xAE9UtzE7iVPX6IzT3wZeVw0bfssTkWeuW9hAVDG8CUGhvTN0n
IYgSeaBiSRlpwwSZRymZJrK0njBkhkI3MjTNE8f0v8T9+aBtAol7O28WjI0Z0C1UFfNp0QUiazyH
GGe0AKuFRqjESokMVyS7XjllKodnsSOGwOQuLZrL5X52vrPDgD68jliRkG5CtIsUb9my+K3vTmdy
GplbX4nDK8rrvwhg9kH5/uHJkV/ngdd3+oDfj23cM4rPuEaa4ez3Hu87QX5J1IV5wlpP4O9kc/cL
cE4UbvdXI6dw+OorvZPeqoax7AzEyR7qClFYvj1vUL0HGb5Glp2TsIy5L6TZM0yKfHKi5wxAPaLI
PDVV7y7FmWHvyjmSzvy/5FrTjVWZIa3FFY8sAmj5MoL2AyF36n7pIS1gUME8njODkbRWuw/YpbDA
N38X9xmOk0twKo3tNz/QWLHj9ERM7rrVgibW42uYiP8ubM19Eihuqq1Ua6PnCPeXMHS/mZGEfeLi
Ytdy1BdSmFyB1l+cJNvooRVFPLtWDV/RiPRA9C2B+AYV8oIHhEhpWr5qBTleMpzB+mG8UBC5i8w0
l1X5zLG73c6Y3+mH0JKvq8fFDCPIRDPG21kRceOWS6csMPc4ylLVcXS+sbXNbGc5e5YVnOHdS7Fu
52+Jn5T78UbP4jY6c4BWcMDWmhDaqO6wvRtyIMfwRQPb4MVZgcVoSlf0QS/CYW0dOjQb3aSkAszw
ocRTIspGtzaHXamnRveen089bnq2cPCwfEzDxVVxueAirDqLZKCWhdUykGzQWbS9V3Ev9rpblY9a
BP8gVn7FuC3S9gWd8aP8cOrkzsrpY3tf3S7VzDh51clHYdkHwQ5zC9yGBvqUgztWDiCSgASgkQ2/
a+/2rLvxkEi0EYzhIZScl0luGhCpoBROAaxFakIOk/zqiSpdz8+eUBegGwXIjuhRbrmD417QRhxD
f9PJAYulDke5jD4XGFOt69QQ997kUz+A9bOM91d5XY31qYla4SYQt4WFW+bf4dUpe+DsN4qRI0B1
w178oGXqf2FNIYOJBdsMeCkhBjABqPpGMk/Q1t6sKdFvD215eVhfsLcua66DgCSYu/Q0sImgtTDh
vPa4kEMPxf3dt8lmcowSNDWFluFiAljxOaAteqcVZVYgZfaJx7trCpl9A5Ee2V4BUa1fHeB3g9P8
XPabcR/k4BtbFqJ0MJD1xZf168yqIDs3MOSj7rBSuD7E82DK3XCTNkf0jxkQxJGA8/mXNoXDWXvt
otSNd3TGjeEzPrX2e62HWAVmZ34zAWPdMCFtt+Pv7WdoNw6KtabpySJ+GoIQj9QeJE1O5DFh+M5/
K53UjIgHBZitPqMOCfLCW4jo68Z8Q4fZYJKURVJByJfhps+ZDAcp2/fUHLI3977ATZrqcAxvSo5N
K5zu/HLq9oHw45iVmt+OXu0twa9Y1UGAY9gT8GTWMEm0W9DDdAGdRku/P4rYu7cCOgPWRaTyoqFx
X4jqFhYgia0xLu9lL7KaEG4TqlCrDnJNIiPdGByDp+2OAo449crUVvhpRSJcrdHZu9YHeNv1hE2t
8Lf12xEkFObUa6pxjstE5h1sGwbM1llpf3DZe4o8EdJTxEcF7cKXafzx21HVIkbu+e0TRVrnkSqt
B2HXbDAZ75dDUF81uFb+uVLBUFBLScdQ/WklVeW6ZhWe05kYrKiK3GfelHXqOTk5WTllU3tMAn3p
OxPivXdk37vGGtYq1jhLqbAxo9xxzlW2S5EXFraRmNErLdPZbpvMTfJjIhJ4tE1/1dPExqbAV9k2
gak+l/to2N+X/yy0CUHo2nEFURmT6zy4DXFxuuWnI534ehPPB3gv7N2tWJJdhOGkKl/Fne9U2xjN
ez+1Ieeccy4SyHDa0YArILL7e2XouVwQf/soJkW8xBWhTDbHJHXrTA5kWlaPFEBuyaSi5ijQWJzv
vlZn6D4ierQmNi7OTiSBQeXmWkKDA2GTHxGkMYGv4PgEnX6ICVSKaxeVJT58CvZ0WVp9WWWnHRbN
0U2TPQooKb/Urt3+GpdYXHVRJZdG3LFTinbqMvw1qYgLxo1t3roUn1ZJaEQISBCLvssutk9RreqG
m8SphQoEg9zBbNm8P4H1w/eoKkeQHM7U8k9OhxOG6CcbDaJ06duc654WAB1HEeXftghwwVwBU9wu
Ch8ZPOPwRWDXgheuZDe2b8i2/Up4r4RCKezMWtESYEreHdCNBLNQ0MKvPszrNALgZhEBnYW3QO06
2/hJ9sC8x9C7LTHELdZaCBc5oUuh5XvSXOPOGp6zr/Hyo686gpC5K/xKDRzFJRQ+myK+dygIP+8r
nHz23lEITmHjDQFj/q90JHWhpYcmTt/e+cKfBfuKbFDHjUKIi9srOKeV6/gXSDf+GD0s7heBl9Ls
AdaXXurpqUlgMWOc5iK3mwPmIvqRkx4d55B8U2Xutlm3mDjgOwwAHc4uF+8JJ9ULOo47MdyZ/DF2
c67pmnip9O1lHix3OhVbKmx067un29T11l76mZskLuNqP5QM1Z+WlmVYSK+NFyCxOV+2dJ6aXokG
OAbJzz86DUs9/58TBYXMahEy3XqVaN/UDlS253qmXd7Ihq9Cdayh/cZO0hBILrAYnaYlbH1vRN5Y
NlH1s22iMGBG5EQAOd8wBxFAweO0XQZRreZ4XPE7WD2bgsCTu8iWmYrq1q5IoqjYq8KrvWh9tcrN
/6OGGEH9KYzfbyO+cmB5QQCkyygMv45TxEgv+YLpdqyqhJST6MsZyCbbs8749iB1I4qaQehOCVwO
goYGZVHcSWB1kjBjTiz32YxlQIaurXnvO9n9rpJ7hNUKBw3PSNfed2sZUBJhMnIva97Z0ixgsRSI
Kniu9rKq1Uw10hHu/9DGZMgYulIm0kmvwJBBsWmGrXse2jUQA2L59m2imRd9vSJPJf+LpuH+3etR
zkpV/7KMdKd6GMUuKeUSVLqMkZXggUjKagnLfYoaOsaJqJqNBT56NKCWvpxmDG+2CYyTf9GwaEHC
h4QSYnIGNgp4o5Pqqdq/ijAaccQ0cHkllLC0raw8H8Y+MvqoUr7m4Z/xUw94LCkaN6NXtTHyDiGf
tgld9CqM49uHh755cK4glPu3+SNjFmX5eNpr622tT6UE5ZoOcYUa3JVAc5vrNGQ5YRFtup4K4tES
qizoAqWPv6sVZZRYcqexJ/Dj3k2rv/3A3RR58nxM8HBAG35i2KecLTRD619uRb1g+YQ4q+27ZYrF
mIW7CS/DddGX4GWi8+8tbqJX1hF9y/yqUDplWcEKLIY3ohvLVvtbW5y5Z+idpQLixn5JVfa1BAlS
HaZfH+Q+kW57DLDANC1yMnsfus4mc7be0XIG8jzx0yXU+EKDdiMYBykRznxncpJF1LwfdNY8KU03
BBH6PUwf6Kj8BT6ldeM+xi52f8wdB5ONP8QTPbYL2llQsVs2dyN2wIsLDHsheT8PqB9u/p+IsJfi
CjUaUyF5bJhuQKXAx/PVTOuqWqSEqvH/fAb44azV2kEsTlKOJcn2DycliWnXmHIfxEgjcjct8Cjo
PKmPkGlEOxQrXnNIrYSUa3R2qmc/lQ0kb+LiDs1pbU9GSvxE4ZBoNVneio2TJClcXWuf1Bj+kj/G
Ms5bLqnnyHyfunEQkgi0LQF11Ze+QuhamBY5CJ/wppPsncxo/zJd4/kgKGtdcfQWcTy5ePPAKhBX
i0wxxbFsSinwIteAMqsy3DvN1sFDtz0ykwrGxu/EN/wDsR8ziTO5W78KKMGNzPyUr1sj8g/5a04p
iczo6MAx7jOEmQzMpcy7pgdh97wY3C+IK9pmYCg1/S469qCIn7bcQi33UP6PbCVRlIOy1eq40LnG
IW5UE3BaFKcmtChhfy6JT9eQ4jHAbhm82i3YC+iIeWMRl/T3yDWyuD0UTGSqi/0aHK2kRTT7k/y2
grIZlfxITisgF4Z9FJNduTTzs+/iZq2bIpG0+vSHNjBzuJJuJFzmdfX9RXv68qJHu3Or+Ae21kc/
MPrsOhRq1p53m6ke1zLM+7KhI+yAAgCiKblYe1W79WyAV28Ir7Ww/7fZelGfxluKToQHEqOMjqrV
s1QN9TTc8Vf9SoqpaoXPTkmeKilgJHZIRWHrLslcnZnOjUgsJVHc5sIvFGium14SkYweCIPXvqUs
YJDMk3SPpgLg+nHeuGHUbtyJp+EoE5SJJnTzttPOmIOPmXrTxzvR//PPBOctcdyeFx0qVp16pTvf
ry1rB377W+N/totbvkSQfPRGZMpdgbBrYfY9pVR5xFaRAse3NlENbOkCJ5wjy5FEvuE65w1j3Yu8
g7sMd1yec0KMRSb8KFIMUf8nLmTP7TrUk2IviwNFfMrbknPJ3CnLsTQdOKfKR7/SrYir+v//tzlJ
IlPig1EGS/67p00dWBw4NhCt/79mXwkyic4tuLQaOP7WLkxrCBIpCtOUhBvMRy2laaf4cZR3wNUi
FZQB57BVVT/jUt5i9QCQBOP0hhk/X2HkEyxyUNl4zEk+fN5Sf+cNsOhxvlOEL+XsWB/IvrKCrkjB
Gd/MmDCXWDQIw4YH1I12jxoLn+9/3KjcO0qboIlSDkagqaIKYUY2gyxF4Cw37dMGjMDHR8fbM9eW
TX+hDONkdKwtoybijsGrcjgHZGaHAW6Ho7C4Sa02AZpw1hANbA/swXe55l7lxOujsXOQ8I3+fAJj
7YzKyCla9dLdZ6xyHdtMPLVquMMDvK6Jhxn+jb3KGtdTcXuDU+1Pb8Si2P6W6oszGV5BHdt6Mfzx
zOIEMWRShmn/5FsKGA/vke/gxircbHvWn5nDhYC/PC4W5/EU1WT/D2sekx0qciPE+xURLs6dGTNf
eNMJV4O9g+N7blo7Ir0WrUX52ahHDvHwYg5NKHZ0OJS8+0V3/1TlqdRmIn4pOinY5C9ETHiw5p4K
W1b/eNzq4iOLv023smwJ14FmGtmqJUx8ChB5hW6qBdxgXzhbmddle59+IBDbDkFhciFuqiMmTBDf
pzP9Ue8A6NgI6lxDHYrHnpWylu7GZsx+Sl+irJk33PGDw36XVR75aS0r3PEPPQUgrrksrcw01DkP
yG28qWAWlFXSAaCoUskTFsOcrJiNzYBdprrOgp1JXpbIwC6j2a6P4HJ3iXgB+CD/HgcQx8+GEaqw
zXGtYfjyuJLyqEc+tJ6UpxGjQp+QAbg8zrTE6RNSDByMhCgqwlJbY21z3DgSTVRbxld55Ri7RxKy
9ZlW/JjxD2kDvzvDPJZ7WnI+sF4EXKsdPKWhqDEmAoMHau+WqfEr7ZA67wJ6cpujJtMQt3XMuPPd
neq/vFaSkOezm7f0GB0lWTmQO5qx3sV/6eRMUJ3rlfBfWZbduwQ0Y+SZVlFtn1VlK/HeOYAT5Di9
XhXf1tyagJelRqO60rACpoSv880nG5Qz+80zg///Wax3tX+A++qXCV1gOSoKikpcVfPvG5gUteNQ
6xFC8xvrzE2aFkIrAdJ+wLbaPodlOBoA7VdNkXyNRMTejs82KcHLsHr5vGqWnJdA42JNTnKMasfO
MTrT9DOnOa67FxXvSKVnrTYWgbhfHImJW34WmrbRMuNUky4NCJvND6TcbXa7Z0+4BXDViX5t4zSq
KkZGlRtNAQdzAxoZ4ufwr60bbditykvQdPO9x2rogUqRruf1hXh1hh8RJfCDW21kayH8Z8PvYja4
52xhKtblo+Z0jXlY0cPs53LoO0OlJcWT20mB3Talj6QwFEtkO1KIZYF1/+ggqc2+m8gS5ftKyFGU
hyS10HKmjgSIMNCoUsLIdHCbNAuOUPCDL0+Q8XCtCoPaB7E+TcJyshfQnMhiZJJvRI9+UzCgTKb3
nmTnmcqq7jiAXFWvFgG4+aSRfj2bBL10wV4Nb9mFnWfqfKVb2hIPcNF88IYyp9nA5FI07oGo44OW
YT46yLV80qfONL5+J8BW32f5th5/cjUmk9nPrBySwESUVcbzHHtO5Z774/uIPaHUSRVHddeO+uAO
/3GXc0aXg83hnXhFuiIm8JjCd159WZ/8vrxngYSgDpa3nHsG0K/bwRRVtanwilkj0FPE10hw/sUg
Brf7+RQ0k7mVjLzAyTfrfkv2cR82G32s8PJ9wvs9k42UG3uBHP4hPVoDotgsydJ7dhnozQEUadu9
AF+WBMy1Ye6owGcZrMkjNByu7Im5VD2yCG5HgBJ1vtUtCYhD9u+bw9WwJxUvzZgaoCJF9LEO062c
TPRKD9egDlFDBm+Py5N7YvLpvpHyZm537Od3pAZoLrWIcs39lzIfNlg9+jcmV4KmhR6TiHoObu7C
oPh/ZYUW4Fhj++Iy1bbEbI1NzgEAI6WbpbY9YL58OWGW9BKWE+h41BnTnzuZ+x9m+So//73Y7VRL
LZ6AUKM8cz+7XqKBu3vTNc7nQCx4MvhSuvPLfPO2e3ITYlOwgporN7ubNGM5MIgJvKEhP5PfrNyf
eaDtC2kW3e6i7hOsEOU3pNOObTpNafAp2H4sBYbHh9BN48MSPsI9CcjIgyUp60zuUYMSAS4K6lar
YybWpq6pyvNtgFJHR/9p5DwoZzzk/asCGFv0cjTTpd7vzR4G7qIHSsv603mDjYVnyWHHGoMmv4hc
KhJQ1QlyooMLdoQ4wFioqzss6KkHfyjD2mOnIjEg/sBOJZsSIgQ1wXDGp3UYbMtZeLBUdjxSoT28
1RgMXJ/IvDYIKTqLINW6XG2JDauWN0M1DIkUHJrpGRjZOilcJTAUN5M4VTrP9hwewL9WWr7eihlw
dLyD1/ioGxZ+MKnX6K13urAQXhTEYvuNMKzDUzPVMdA1pclj0WcpNoR2CO6bQEXfhu5aRB/Yf8qj
nAbvcQ1/C9hY3yp8x3txS6Ho/yWG/3CTaf4u3mxibABWa7zK+xH/zi57Q8QnH7l+xw1EL3ToSSjn
4neoxZShzCF0T8RVR/ZDZHjnv8H8WXdn3wDR0sv+BoQ4GoMnzQCWcgie1EtX9LnpcQr7j/iu1+yX
BVYO381omc466uFU6JRV+0XYfHbBpAdnuJJSSD0Yj63ayqc5RWa+PA/z2VptageX0SMkSNSn7KtX
EarWLcOEK2kCeVZeylWlYfvRWTFNtnlEjfhFbY2Ve4c8GfA61s1oPvrENXWb3TiSoJFKRfQkDiog
ylJoycaVXxMmNhonOQzgQdHCTB+kE1DgS4etBwPyZKB/tKRdtv8pWKFVdxUOKWN1m5J+V7TLXtjN
QReSOcz6J+MfkJnQzv4ZKDaTJSO5ytisXx6XCc0ZxfW5XXAK14UrhzP8NEznhc1g7VwuXrapnwO2
dq5pY+JDOh9c8KniBprlWocyZ8BO9yxAjxGamqN4RYJEK292GZUcm6UCLn39pEc+ZNtoCYq7ZGd7
Nsn+TDHn3rMuVxoXFlZz/eWL6zdbTUV0c1PhrrUvtvadN0Bu5EEcnI7hc/VVQzWy8pDgYMc/P+m9
sq47Gph1wA9fgargXs4/HrkI16FgRoRttTmi4OHFBxLohLzKvQtjr0UXrP4UzCCd989PURFHPCsG
iHZf+13HL8o2LmyrRwfVltvcCe3YJZTc7B7vgPWQ3dI2axHEvj6ApA11qeeVdvwNTZAly61kfFkO
exnGsVXYpfaoHzxe+K7EGwulXB74jxbw84s7ogFC1j5AowXYJA3msuA77o7ruDz8+0oX9N5IROdo
Kqim7FZPGYhBphAyIG1jJit88FfEBAl+AM3CxDRqD/kDl9eHQjSE+0UFVFLEt8azBqKaZOG9DhzF
NDwrynAfnhNxHbsc9lEX5rr2esQ7nVXyCcOcFoqlGudJoi3oxuTljUdb2WxzBStD8vJ51XQc83LW
Q85X6Y+DM7zuXWrdpfva84noj3lFBBauogfUaYsOzTHNbSshDp7Eqza6zk4Hqdwyn4iL/hZDPV08
yDcl1S7hiBeFS38v5WRS08WEEhr2fjHZMvKK1Pg2bS+IHE4boyReBmjgFed2MKkEDZ3ZTj4y3U+U
4819+VroR3Y4d75YRtZKOeQIq+uobSs1kkj1eJi/tpwK8cI4c8gpmEprZsquwyCC+DbjZcy7DoFw
hnGvOg3qRhn9rgsx1hh1AaqpZhX/Ic0Ms8hYObd3i1Y6prDw8t3IroI22IVd2hAzeLaW6AA3Q3Lm
Uas5QsfabWb6zCPN7pW3kiRk62oEm/qHF7QT9qMOENlPwBjNqvklNanK5T3FDI+/WCmeTsuedI5W
EPjx78OdgP05aRrhVELcGQxwuVy+Rd4GQ8zGa5pxaWlPtgNhN39iaQ3SKmauvwq9cwYXddqIArin
Xy6NRfA0KGPZoWwsjTLKxmniuuI1z73Ov/Wda4Re87qSl1GJEDmZOfaGHbNtKo+/ps0Ic5s83Pgf
mn/jr0JUN61AE/vPggm87ScjzV+asllvHJcC3x+wCqus9AsqHCGRZnvB0PyiEXM92jFA3J0DhQ21
rNcd9yFQ238a9nDuhBcSpzOdN+JS05uSzw6haiY250vFzG2rT/c9BFw1JvA5KLDspVkg3spyTWOl
4Hgp4liA48U+4n7DSeCSvIenN51U81E2EA95WadwCsOHHxJnWx4r5UeizF21cPCc26Q0jlDKoQZz
EY6YT/278QAWRx3fgB2sKhebLwELKitNhVcw5qysO/wLOikthOOQpZafR+RH/h2mPNTzlY6mls6K
Pls6v3YdD4Wt7Ob0Ord7nRAyp79dG8SzH9BknoXAtOkSJfv7Q259B5x3/0CHuzJvBj0mg4Ankb2I
m1uoJ2Mak3AXNVXACUFq7MvsiyZNptY7fbxbxf7Hqe8eZFQIPFus+dsZqIg5MwXHNrxGEFpohWPw
0EzVTFzD0MBd7O4fTYhGTURMBvF/374lS9fBisaik7DLkiQFYy5sdiNEP0KZ46WVGj+Vs5+rwi+1
BsxNc20SiE/EPwareMwc9LrJZ6ctSLHD2ZJg/l7VKEn5U2N0uNawc9KeqCfR2/C/Qnlz8QHQ/CzV
X0u4/eZmQyBwH97uHHqtGnsPiMaiBfxaJoct1truPZOe1lKu8Jtwetuj75i/eJUz7cpJADW1wENp
cjXl/T+OAiIfko/oAbzRpXoPMAM+1b1sxnr3hqAs6MzPC3+VM9Lev+Bd/vP1S3omLF8nVcx2m15E
rejtzb4khtWSLjUHY8ylIVr+uet/DuWWTmskaaSZ50YXpk4KcNAYIV0UwgKCbKE2Kz+sqSBDxJef
AWpfQUhFEWWH63VGDhHGEDq1o2ZX62WMmK0ZGWX6w1vBDhl+1wxFOllPDHQheWZG/UGZZVf775PK
lZyiPEdTU7bR+CvbBLYUCWuWIRQ9aKEA5uk6HuvtiIvWXLeomCMt1LVXY4xmxTM/+k3a1WSdrYrb
wsUorH9iXA1XU3w9uNmosyGyF6im4lrbzHRAbP9uuZnUUXDy0Pm6L9iu+ZbWz8Cq7WggIYEooNu5
fK04W0iSUHxfiC/6KoUBxbCUnndWASCh7xYNEv+U4gw9BDGJqqZmZdw4oP3DdOzl+Vrn1h1WJF2d
vAeLWOA/1h8fVA5D1jJGQhYAny8PiKQ60xUqnBvyDshSVsAGxxt5IeyB8oo6lDyRTykOk1Tx5qTH
MEXMmpafdRaotKfOk45E/NYFbg4WLHsGPefzsfMN9mX8Kdgw2gio/deGPzkPy4B8s+9J5E7Y+ZKk
0QSBFNqlZMwwLmiDiTEMErCjHGOf2HxXwpjGrjkDTHmUGHA6zZblphHOuqBH7jMHpLfpkvNTBZEG
QbXSVgeRpYoUSpHTlijBsyhpsBOSgKcnSaTi8VNEL1XOWdJh2JIz+U9ztDY/9KZbm7ewUynv0o4y
KgdUC/JbfnSE+9InOHm+lHVV9wb6MuhQCiyJ7RxeBLEm0mrWRSQm183LLDbksrjs7F0NZO0ryaGU
9jkyKajIMlDR4T2fwjwn7+lUt2firZ3gwJc5xT1Xlzu6uVUwMC0urA7lEMQoH3SpyzeH3qXeX4UX
dRJ8y1x8xrzaqBiciMZtR/NiYyMTrwB1m2HslJe4FTp9hkTaq97FSE596r/r33mJh0rip+o+yqz7
0OzgNpTGF1PcM7s+4gYrPI/7LkIZHs+Mvt+rZiqKMcTFM4otkc+WykURqh9URPhptdXI1+00KTUy
Mej3D3OBPniVpiNuzW3DZ6rKgjv+st3OeFUstbALk5RK5Fy5gfEuglHd53hmiJR3dm5ZdGDhV5kO
AxgPDxCWJaLbSeG5bk3+DsttQnJzrlbAwEYKfmAT32I87SDmxip1vw2Xe+HpAnJCG1Vilvn2Satd
4/7k7K9NAG/a9TPwpzsT+46Z3gXDS5F46ltrR9tEdXeN+xwZc/Rl8Z12+6FS/p+HW+4vCnSbx5eN
+hoKbOUIL7XMhisyfq2dlewPGYNYOZ5PcvDhHTDfaxvGS/zOtSNEh8i2TMAhK1WImB5mGdldrexA
TabKzh9aihtU3nAl67Uix6//f3+M2ln5cALjlvnIrWxUR2YVYx08ZYzCGi9EDTa1T1N+qpraf5I1
vdT4G4mxvKaEiba/7/V6BoNSV7F5eP35cK5Q6PyDuoZi6yAYlZ/KPM28m1NER82RH5+brCGPGjAP
zG3R7hvJ8JklzjDpPW4lEt1wP9c4q8sGTe0zgQDAWDJd7IBPTJzoFGZVRBIEJFGgU/HdN6qz4wp2
HajZuDHKaDRtl85TIotO5Ke1u+wwQtIeiM8EI1V4qeN0zt8jFhCQs4nVPgRWvZK+yZMIznEExrBg
NLcevXPfLbuJiaxvU1wF/5xHgECv56ij65exax3AioPtlJtDLFtodqCONQmUZ3ZDXQ2qK3Qggoy4
CjkWXwHe2wfZ+0OFEvPmSwQoi7rwlHTICJbWHoO9gvQ/lk1biUeO+LGbn6eE704fvezgFm1Q98vz
359n6xsXndtxMFeBXm3BPeZM4NjUf8Xjxui5oxxZ8GjW/cWpG1o9NPlUSxWCUQost3HhmuxkmpVT
HYhdXQPhVnwCQRr61PSCaBhy5qHQDtSVGkfGO2UEeA1+7GuKfktL0fJqOa5v3F+nE7X87AALUoGg
pVkBzKcdrEnforqVoKN/82obgruaffBcFkWJA3BEME25AdtGmnrDHwLMMZJmyyHIRSbKpwnr1GR+
ixSF6JvGm2xXjBKcjmnyyT1I63j3gfZpNCdrdiJ2iN5QO0HgED9+zTKlb3Ri4IsY9UEzoeTzBTCy
R3mhRMN2WlhPalhCenH3ATz46Y/mVl/SMWqtsX307J5gqzlI+Ek6trmNIaz8Iyj9u7EA5hOLJrkJ
owzM5D2opg+UQ1zMDNvVSIwBCOyoPQhR64sebde4o0mhObzqDq6OdvrN7u6Htdvyp+rC9S31Zrrz
KuNUr0nDFjTS+lBRPDmnbL3MP1SuGi+TRSFzl8Kr04SrsO/WxQ+730r0utSzaCRtLGEkEdkPTNWY
X1e5lF15oBozqbfpbpNEDvfXD5WG/R+W/yvPzC/awf7uCkDNDiwI0qwd7kyAEq0ImSMEvWJBpFIc
JmWo7mnX4PhkMMEokX/9lHAciZPx5ujBs7VBG643iltUVN8dB1tg7gT5XfXJb979al2ObTDookHt
UG+IQ8KGkUg/JTll2SWVZP6E7g7kax1vJA+Ik35c9CxMIavptXJcHC111cQ6K5lf6k1NdIClsIhH
xtfmtEnirMhdoyl78tVue4/NP/10EUS9x+qy0dxNBwmHxEH08AWb46sQdmuuBfNQig+zv1cESHPa
bBZ3p/qwyd70ew5fFbj/XrNdX8jO0TLDxuxDE07GBZz95xZdWGUa7pC3sSfzkRaqoJaUX+mSXr0M
wfMwP2ewX8Izs8DkI0p/J2kVobfaoSScJb4eiwwwaY/xkZ4tVrsfiBJqwDSSOtBuUFAJ7N6H8qCA
LyKiM0qNf4X1+ge5D7oIPJ1BjMYrNrmlO8JKbg37XgajFMszXMYAdzA1ATJ+QQI1NvNAuogXPST0
OMTx23Y5DPk+XSOOv/Qo4ziIzGJN2OsvX2aLWbeL0QnEE5wvsgEQVgpC5OLO5+g3n0TUgtkxTdX3
t1bOdPY9qqe7yNr5wRRi5heFyCQeMTW8vCMTWv6zgwWH3/ERQEKjQHOceX9BOkEIJs0yYLz/js+9
IKQOzWJhW8IGUJHO1Q+fbsg6Kq3yI2FkjVR9ULCeFUpojGjh+J3RQLjKa9nLq9jR1wrpgajeZO7j
jQyq1hv0RQX2kREkicax8VfAlUFNye5+HdNzZKUPK/x1kSSkVu/hmlYTy3XrcNz3ghUDHFGGr7Qv
+nWNa9UYzksSV9UFLmD8/DhAcXk6LFvRZvA+Qpm8gq8fYDhIaTXYkksi7gOjVwth1wfJ5PDlUpz7
4LULHANUjAi0sHlzYvZh7eHNGclvRLUNDoE0TayiR9IxXEmZIFDJb4WPizEVBneHifSJFIZDGPMD
hZvWkCnJMpFFWWzogTMxqY9lq6GFJSTACvFcCWi/7kFdtyNo+KOLvLFv1Wd4YVQPF5d0m334PJIp
gkmDQagLVZa/xWP2f37EXHa/CWj1L/mGKnCFe7r4Nt1zIxwjOMtqE3x4o7GMIbg5oSJihpzaoBqz
gpC7dOH4jOphTBwARP0714tMKgDN203IVe/uAzXLd8ZnHtyFTaV5nnw/SnuAjmaY9TSZZ18A831D
DfoUzaiFASIH8ieKwxapoSLUuzfJKCzIachae9imj5dnP+atNScDCmqaVHyFdOPI0JrfdlgFZMxL
GmD4XVf3QoIdbg+OiOWhHUNtkr483lrtIvKOOG31/q5eir+VijRwdR7D3v1blASKZYmCao/sYTpg
pJckbo3pF+tnFuwaFKvgc6Wo7V1oeKpfMz7XpkpV24a43wd1RTCVMIV2PbC52BV/5XpdgGznbIXn
t8tyo8bG6cPBfAceilW7i+OFuR07VQcIpc0GY+8WTcksgtSPT8zgNwSrXqKK7GM5UIkCaAgmcTJ3
aM8dtSeKM7P1lk04gipTSux0fTM6NNFHUN2GIi2LVXr3s80itOAGORBnZdab22/YunQSZBuxFJw3
Wzq5/k9DskLTsCna4RgApxTOT8jgqrU/tNrP0lO1vANUhOXZvWy6s+NLcRtYcqNGGkr00esQKGEB
4egZwbDcqpp+MRlwOSfaCgbUc1pkc3rZEhZ7ImQCK0Ip3X9htoOs7XS2d/sEmHy7K4bEpTwNs/0d
2LeNAoTPgICeN2i3U2jauJIZ/WfLaHL2wFJvdYgH+PyJCuL+2Cw/FdaFdjY5kO8Ahi0XHUfgeyUL
vWxe4ThYUqPk2KFAfjGklNcMO81ozwIXqX4lRGOLrkyUm6xaMFNqUqF7sYiLvbktpA/78Ez3Bmhu
sbF8Qigb1oBG5ip7edeGDB2UjtzrWSMt6QI8q0RGNZySybMSOFkQu/Vuz77K0qUYLQy98LuvgR0f
Q5u35m+dK9smEK1wQswAIO8taAdb+Su76ar/N14SU6OK1Pf2UUKp8hlKiNYLOrS2Oj5Z2amwYKTN
QM1T1rEdq6+OyKMYeXkoiyvx5ftH8ayLZKxOfHEoDLNZYXgvKpbYI+50H5/0ppeMM7kjqOMnVTKr
iBQOL2DkP/7OU1+YWh8HG0603A5I9HWoM94ZMZ778awwsdrVxxn9xbgmMZIlWNSlLDenbaNFtOi1
t+iPv+YBIfXxD+wmjSgxW9o2QgrOzKcy/+Vt8Mh1fqQMqHVSxSiCEiIq8m16IlmHdlNAzQXl5pL8
U3jRVwZz/QGRohDr3kzwoAVdDf8K/Ij0tW6vl8UgDXoSBIwX08Ry/iTXHxEiAzZvmsA2YhgEkozI
2RgaUj7Nkh/SxQ4BN9LF/mbpimIqaCLSu9y+04BA2hNPEp13oNR0Y3UTwW2EkQRxeW1BK4BKk9rm
np7Zlff14qgTtNlHEe3pWvFymwBE2LZFDCogekBn31AOL6Ab0QvJaWFEE5W1MF0YIec9b9Ity8gs
g94oKYwgpb+OwP14V5KTFErm4hYX1YR8ZT+FzuZHlyPkNAIC5FVEj60BUFGh0mdDoRSlkHjTeINT
/JB+dOPX89eedMsJyklQmaXHC2NL+tWzsMbPUMtye8RAxVcqjQBVFQcc/OcXARkEjFMHxSaCnXIQ
OA8SA5pVc5qWl+p+tCfQvlTwG+i46pt5Hwf7cQy5vgc8mGKXjb3VVJ5xReAS2Hv6qcPTEn6kckWe
Up0Gp5f4cGbZ84/CMsy5lvF89iG1nh3nog/vW9WcU0aFA1s8JQPIrhsQM14D8mS3JJBEvO+HECpq
Br1joQ9NRMsmBHwBo24QSWGRrAWkFp6fM+rsSLxdwArpS11JiSKEWWPO3jTzbEpO850KjEbPessP
+CcsOBe/qiFHyFQHE+58XKlNzSGrLQc9Aj5H8o4hyI9IrhZEWk0uycggl2IvrIDQVQ5La1bEnlGF
RnmfbVi4uvMtgxRuNAZtvjgCS4bUDi8lUq1iyMcWDb4Ak2C5Vbw0PgpCqJj7OTLEpzz25nuGC5eE
0n/Ye1NOmfI5n5ObStqpn5welPkBuu2J8dGOEz7RynBuCDz9Q0oCNKtOKoR2kvoB4BVPyPZDVNW2
HLROd+OG5xtUwYa/B8GoN+DHYCg1WyPSXeX2oZfW8ILUxHRSmRyyAs1ORfKsooR7VCGSu5ztP5nu
bzcksvBuV28VsNTCwQR6TbEXaROrXOkLHL/8D3XLF/iH+2QLJXD8BOwgGfEtVCsy6YX5hMkopLkw
AO/ruJwcSCxum7IusdsGosr5oiYQFfmj9lVZ4SI2Cwc1S6ItfZ47wWOinoVORBL0TsOG5fT8JzDw
lkjsZaWp76ZTjndgaIo3VG2RdkcXxGKtPER493n5RYsbQUp8ZAus+8tvJbc4E0GGMHILKWjtJDRG
Ddmo2GwK78p8YZLXTzLpdMejLZSueLgyxy1h8ZVgCqJ2TZP22XhmEOtCy7TrHDSWDy2HAXK/Y8Bp
Eg4vijJnnrOoh45m5yndzfGrJwr8oz7QTEJtaHwLSUmSytitkgrhsB37Cod4hlW85SoijHOcW+Zv
mUM1dgUB6NSGoYWDgWkFTzrvmzZNPOpf4AsRx0+e9Rl7UntjziafjxisxT3ALEj7GEwATnIqMh4p
pr8xkakmPyM/pNJGgV59CznJeo3fdVuRGDhRNsSuktyg0GwAyiHic7OLaURBvlSDaetzeKDxmQ20
jJ9a/7bZ7DH4kd5zmlAwBhJBSzGKFMbbS8ARZtJBDckjatLxF5KPbNTZwgCIXmEykCqMTbF3Gl/+
07VTVO1F5OwXCYG3MyR6xUO0LKqrphQYZi5fmv9HXYFDU0czEK7/lG6y+7RR3vBvRFj5KeAwTlQ4
M6w8DiaspbKnlIZdV1Zp7kQtKRE/1uriwftUcvxpk963l04zOYuNiHFVMfquLTmdQdAM1Kp6KQ0z
K2O/R8s+v+XeNElyOs8NtJrDu7sYaJNN38r0K2eSlA1ZK2sLfEHQaoQPdUePRaDPVptL/J+yGhH8
JD1lE+/cgUAPV3ce9vqHZvQml/aKtzhCPIMK7kDBDBw1bSLCATnXlojXDr2ZbjtbNE5sIfvsmg5Z
c2U9IgvE2ZinZObYFPvqYOlnG+9yA8SD6pESd0z8WdLb5Z5OnyTsEwmj8S3mv1iuMu7jisivAnoj
iT6HBRRoyR9tLr04wkU6m7cDfzPHGQQqst6r5mfyfQdfiHRmvMwI1SdiDobn+sRiGOy3zC1qXWrT
UXfIe2d4th2ueB0P6i4hD0Crud/omQNrdsUqz1vWdPizdLtKFRzN/BCp6ZoUL0bPeCQYZZlA0Z3C
d70xALFqy1SSqvsG5CTs8nZk7IdXJoBweBt6NAwIIHk8KX6PkzHb+w/fLPtfZaUlfXtIeTYGkIv+
+6gGZZejBgePcq4X3NwKz4GjeEnBL7GkP1j0WayFkT4jesi3kHikL8cPK6FsP2aJ7pn9QQPw6e5G
q7uNk5kzSoCNmy1TNYY9/CACfhD5qB5gzRqlAD6CEUDLswKr+8A9EUnD1qR93xlD7vLPT986N7EB
8KJSlP/tlKmWSK/Vp3rt1uxnAfoukNYFYUGOqYzCrVcPGgV6e9qUIFAFuDg7FWwPna29kBSF7X3M
F4uZQHTYeLm5ebmrgqruLDA6jlta7HmLeSHVfXHuB9dt2o9FKUIQZw8KArQ5dg30yOlEPczYvtqO
zw3gL5fzbSs0wsySYnkTtaQesOV3pYV4kXZ5A7ezmCs46ro6aIpFLWg4Hr3EECEq7GtAPFqDlzLS
XQkqQIfQ30R/kvEMNOVOvHsS8eneYj5PC0tYvoDEVt0OqOSmr+mmIlycMLp1RQYFeqYX2WAvxw/S
16BFIVEfGv2yA84HtjED2rAYzyNInuPTZXZi4X0V2nyoZzJhN+QAjmBCPQlWEmNH6/AjlrUa7kFh
td586qIuBzBz4lGj1f6P0IeqWBikCVavn77ymI/nRsoAIEIHpwCu125jvFBifBF5oJwjY2ytYSkV
xNm/PMSqZGpeF1H5oA04eR8Wa1ctAhKoI5IL5JGBGughpIZjeHdL+DBVAUMn4ovSa17BFzurS023
e9FOZq1Y2SiJ5iPGKeVqZGgFtcXZT7QDmb0Pzq515BRkuNk135lehvlIr/CY55Oomgjae7FkOodM
BbK7Cvs9ZbAZMYQH9dhiITV1QWmnJyG9Ba5FH3n5b+tBIKGP14nI0ljb3mmnSbfmjG6d70hLumVj
zYty0/RRxAzJphklgh5wulTikRwRR2V2q5xFkh2AujB0lQQkM2NDaNp16QQS1//YFbljZwrpAJDa
8PrbyZ6uG94RYanSNwmioO0ZR4lqHZyyNaQaKSRkviS6g/eiXzIJxWk1EpapSIaIgfQwcOr0soMi
xp3ygLYMRaJ1pS+b7Zx6b9GcsBNehfdLd8GrVCVrPuPaZHvljbCBXAmjtVZhYrE6sB5MoTg3ao/K
qliMW51ZpubPYXzY6JBtDptxKHp8S7aPDcMMzZ0wc4GiBBzH3tcYzuxmsXkQrURLxoP8QB3rjlpK
dGrfQT/GhGXWLI2mtU7NLAeoUQlFtGwRbb+9hUTr2GZ6MYZzMkSSLqPBVPR8uIxZWIoLP3f4ZID0
34c3+HVw4kuyfsy7aoCZnwC+kLszP2ukrFKJ7a9BwXfGKc3N6j8DRBF+WdbdLB2SiiVN0L4nQ7qU
wh/tWJbiExXjjuHS1Rdn+3k6fABncDOFko2Hjv1afUiiALTiW+KOZIxhPvebMafvzvQp+E4QceeP
vAJfUhcwh0QQz2AQ+Ny+XN3KfkG3qFhBKwi8tdKcfW5gRrC5hjonLYIwplyy8iML840BHNuo58IQ
WKqf8snVuvvhBBw9XLRAFjmuymty+S+TYS8UkuQBK+xaG0M5R6wW7qsDBPCk3ud2zQC1/yab6eLw
Gau0sZKBeJGuAis5D+nI5gza+08DG+MppQXzpY3GrOHz3S3C90huK1yv04h99A83gjBPSXgfdidx
gGgigXda3C6MxFGwPXReV6xBu0/tLhHCDRNOWxF5abp1+ZMWCp3oTVGOPZdhN22zCqy9/6T/zoBx
hJ5QfLN39LsgNtWCVWh9R9KrMtzY1nh9h89DUhdnrVRJphMY3ZnViqT9K6dbkCjVsi28lZqvmpPQ
1IGxjby/KZhOsAwzHmzlHoctOg0GR1kgst/mGXm3aUcp68cWlF/XBAndXE147Iacukv9CqWsRHyG
tfN71z4zVMk8K2vuYckqCfOPtKkTiDYmbssk4+Bk6sBUJa/nKuhAeBe8X3aAwULqKSNtDAnxr/cM
tFVeR4OOW99wQljUOhcOn44I5ejID7Xn3qzYvxrcavJQVVeFV6com/lt/LkKkB/ciCHg2Cu84/+M
h68DFNAgguCcyomnTsRqBwi92ZzqtDKnWIHfoEsViTfDwpzJda6l0C+tkuT51J9FJ9fIdHsjHTuU
80pcnCUD1ms3jU38cRaVpO5gj8WUPJgY7HLFWAacPfeMm2Ls0L0Vyp085qpdVo6KnfPzy7iJl65h
ZHgo0p3SpryzTXfaJ/GH+wNSP9wmsGV0oS65K7gv0Wk5D0aQQxXFZqYgw8MqqbejPHmfMiAv/DV4
7GCl5w3rfYbWiYPlu3fqztxLCrGkFNGbXtTKZk3gA2HCfvA6o6dF3a5owkvhaUsvNWnNB2JOQJb0
Cb/prfHM85JGETwj5puiHCTIA70dqA7aCpX4WuL9hLsdKviKfY/g4QhDv1IAaKhoXOGsuPmx5aDC
/Sf7JykApAzhzHN5/vwKn8mLCFlBsOWb+q+6iWm/truaFwVl0xQMB9aBo1Lm6EBlR7Z+EcX64APF
flg9XKZ+on9EEBNoyHaKqZzkuIGnTe4lFhXo4KwVLda/5lgrbESNzwm5uTUXnpoeRxGDHcbJjvv1
l5551xNQFZF81QP9mGRiQOjsnrHhUhH778zHhT2c8TVO9xhf+doQTiAwM8Vpn30dLazEsJb5TGnw
gfKi9XIv3HYiUhuZpImLvJtvE0/P+TVFcEwkm4vFKGHZ54p5lcQHFcqVwVpVmqAx/KAVxxCaGgXR
8Kz9PJk0L7AE/2Jq7j1qOVADyjegd9Q1+EWfVyZbu80AMmzO9vpGfSkl9oppcmDKipDax0T+gPuS
BRSiDhhi8hCw8avvCvVbN+C4zKJ9rEJbdf8NcX8/wUBtly/v6mL3wL47Jw9YUOaudFyxwXgqVVhO
RzoSxBmfKfBuEg9I1XQplJJqforfpknz0WX/nEY4WGiwH6C9BjQhtzTKkfKqpuB1+MqMW9zrzL/v
dkVGLtSmjvCAACAU7xXSTH4nFGkKJbCNCQ3JviQgeGWZPMRyWQEmqpiylA4ZgjyWQExX6ehkAFxQ
bjP22tyIO2YmX/EIO/LFvkADFrSCt0rO71M5bNzdP+JBUyk95UYahc5TqQWNLiA+41zGY7cKQoDo
G+fCMxlP0X6R4uv0vRT1BnTRySzTnEWp4EC6+4o4rlVhs011Zh2lqwt0Ndd7pPrgLul7FYC04Yi5
A3kTU9Ecr11kRYBF2gjorxHo7F+dXcoOeV1i/KLTXQZMI08tpmcrIV/zeSmH5PG2+7dDFA6uDiOX
FOs1lO1lipKbmLYT888vAfQCmF6T2c98oMcxI1MeQXO651L8d50xJwjgbCmQlfyES7twknE3npSe
e3bpRrkIbc9vCChcZ02kDF83c80tfB3+zeK0MCFyO08MZ5IUX8SFOsTvEhx/hfanr7u5UM5emxFF
oUpFgqxoJIiD4O+lPIJNAaWAa3qocybu4gyZ+Q7bSieD764I5G/OTy9l1SdnePXDpJRkcdeVn6ZR
J3nRBCxw/2U0ejFEh2B6jpnh4rVlKcMVZBBuavBaHlTzEpRt5aYO5R/l49I1WtmMHWLfgZbNqcH/
Ugq+6r3LPhynQ/D8P4j98d0P9yRIzwOPSpXsxefIWU98OU5FbXuy6qxKb2+vRvLjt/Jjs7sCQkc8
d8DfizVCltynaH4DYRPEemdrxTVQDsVWSQvXL9UHW7qYRla6NY6Ra9aEToPunyQiDoK0aj8FC6uI
+HKyHmBsAlDfkCEPnnBpJCSZgsQyIDwKAV/ti0CHFQaUj86SiQm/W9yXxoBevp4FXypmDj9EOXGP
ee3ubXaAEiIbO+6H5PIm2/0CtjwaeqMQLqwfa8K46rQD4QjHGXP+K4mTWCzDG/Z3oedC96QbrDHz
QOpyfFdqYaNxYHjNahrKNsvuQV1STdBE9vjSCJr3x5/R1evhsXv2w0sxVt4QTEXMv1eCOVEuWjv5
/yeXSv7b2afJ0+8gWSUdTnFwjCY7mdCfHgIO27YMpEzWh5kDWP/qQ+U1lZOM5oxKqbZR3b5aYVl4
7ajQORSg64uJeH4mMD6tkps9EZROm20UZ3FzPxLaEBrOU0YRVrD8FC4ZBE9awXPoTA9Yreuf191O
zCLV113aEsZ0omFF30RS0SWdHbUXpC9EVkyb0QX6f16nWV2i2UckcUI60tmpfrT8+ze3bNQv430d
eMaPv+WmHBmdwLZQ1nJbcVtBn8V6CrFEYXO9XUAMW+SLes3zbtYbHsh9IdUdSx8UI1CiBd3J9PKi
YqauH8p44lnVapfpJNuJPrrXbe5tzg5pUEXPkAytJKbthlouZRtXdzshkjv0JNnNUu+psnEYBsJ+
0XFK/lbVj+iM2UaN+mjMyLHcIWcoDiNBvl6DtTYgWYDGd3HmnkMj+cJscQDNhq9S5O9li4AB9gJ7
87UzKTd+kjUQCfDIf+1ml+ZPyecZX5PVopKuxMaW0xX9B6CbtZe7cyjBkl5+7IEB9uZoF6UtDxJJ
Axi3VvRA2R52GaZa4ZdDoLIORmm2300P0pfve6buUWuKDCrweN7sEP223I6N2Re+IQBwUjLlM5bI
YaYlEFDsciuqtL4Vj6ZD+kV5bZWwHabNVk4zgQnYdPBf0EPRkDxXSP0teltDz8Yb9Zu5+c50isHR
8UxLjgRUeWOvqUEMdczmWkYf24PInvag6YQab8StjHPW+SYeJQln7Y2HoQhTAreQQo9o+hYtB0Jv
tAwLBUUWCiS7q5/fW3MLfF+UmLRwUJd0+zRbcs/+JvbpudIu/RQuJqPN6L3Peq6rilIktB7sOnws
5ySy+W/Mw+LipGotQebEPdPoYhUpr6Ova2RJkts4MTfS/dfnQWWbsUd7DO9U/GteySJeFgfLX6di
MyMBV4AFJGvfi6N2wX0dFQOXuqdntfpLq3tWHNHDbpQ4CsgKUJqxy04LEMpvLYimYIemwxGVEDjX
kLofDynJbHazbh63jSelrrAWnDeNCMQBP33cHUF146d0V1od5iWi6Ra2LwYvWEOoGfEODxysATi9
Er/8w2tvG1pXoUOmno8C1hq25Bl7VKnOr97DYf1kCi1bAh1kM1gwh4XZHyPAw74xLNGYho6KJyNW
Py3Xcu+J5bI6AthDRUiNT4Tcxecmw09SQMaqLfe7WI4AFIGnxLBpkYm2wJL95330KCKYj+7y0xmW
dNnq/6R3zK8xDIpgZ8WaIUcnJMv4EGqLAdQ/wnJf9X77GX1UgCau2m5uWBiS+ArG/5aupJ8ZuS61
MRv3MlR+0ZvKa2yXFT8NiR09VCUW2zFLpLzy6Vk4onTtT/EL+9D74H4mzpatlaXnm/JZjvScmMiw
YiiwND+AxHcOI/qKY81OLbuukr1shFS0WtAVVbZq4+hL1rJKoORwD15EFxPUIeQq/Dy7+RWj0MNt
AvLqpTK7Z7M+jJZVBFadaIyET4TB6lkKrKX6J0eI4pFDe62obiVAuLUPpCuCQA3YjJuCWITKfcgP
zTEMy4yIaqtCDE1bGfKsHS1Zp5ZzrZf7Ue4nkl3feGwVnhQbXb3IKq0FY08uuB+3q4u/3+oIIYPh
/D+feDlVjlSqHy3CTbVaciK8iFSGTnDGfA+7HTnn9YPZszXYRI+xGRnf43JxNOlct1WVmhdFdPat
sLW4aILX7F0uRUYwLPeDSJQklJdDiLV18bwFWsuJAAZLVoJ/TZLRCgOe5GTNzoUaV63Dyc29+rZ0
7QjCnlev1EpjyR8asBsfEOI4xtlZSW2oXiJ765jsZxt4YcSzCX5xTF3pYWlfS9y+FHwG3CmPT/a5
qsPGhHxz3Tw/wbVWJlIsEanh+z+zwOBCiki2pczUUHTn9TinQVedz8WJ/0taFEj+9tp7tbwgIMAa
rB/UEhXQyTE2gZNXRdWWUPQr/chBdGC1/zHCTc7tm42Qq1lh9QlKyY5oMGodONeO4tUEx+S47m27
SBKeTXMd5uNuxRLkZkwD+x/Ni5jhsTict3zLs95bfbfyzCTkJ/dHHVp86TX68j+SajynvSD52JrA
LRqNGBKj3qCbPys7XcfSimi/aUKHZpJubKIkEu4o3xiZmwuvryWveFGBKxxxB1mZkKFjfaXe0lB1
s55BvWN2oBFNSCHkoM7GK6RgEGv8SSLFZMvdhozsB4IOqYa6VT+GUzDzSTBDRkCsgV3DDLLSysf4
HvT60MFdADhLTyTo7ZPzgCLztzdT7Rc7kFatWhhkx2HTM2Ygcan8x7Q1KHmkPlIsqA775m8gEYUA
yTZrazceLmjMaYfSjgvBavXbRjkqd49jMZPnx7YkxFKbk6zxvCDyuSsuzys3CQFfeclXZr4clrbK
QbaEgLPxURI31rZy6GXjvuIBy3BW2CVd5U6py4wCR72Z9EXx95Yt/fV9NR90k53n309YChs1X/7f
iFiRoGIdkr2YZpxrOytRJgHcUwbsnvVS5kExqCE1/XZ3G8V0LVMpa6JlUzz3Atpa1qKl7LYOo8Br
OVcu48FXJlrkf3QhEy+iI2sQaOl/VjaSj4kt0Jod8IWNxofgwds4z7Vibv+hTVokltey4KLq3bE+
uSqLcbacuTRIEXazpIGwM7KhLGHzDnBYwiqH0tOd2zX8tufi0tWRUWDuqo9ReHSOXPRFMtnGQl+4
VZ+6bv77YubljMAAs2fYMW5tRXgXdmiLtxCLTYySeVAbu4S9vaNwUOUKZ6MHH/bTVObaC2S87wfK
g6An8YhZ1OYv3JikmK44xW/NWkqkZD6sX49esakjnM8kY65AEoTusrbxerf7Im5hcqgncAo1YJPL
u3o9vLCgnLKaSbSNxb8mdMUHkcGli3brFSxi/BNP7CJbxTJQRr+aVH7cYAK8zVnF1KQwsJF/PfRC
6Nalb3aLl9eZvLUdoOZYAmPEB74JPmWIfAoiE75jeLfEFywk/XFXeE9mSBujuVXYiE7pDfCwr1um
Lp5sFOxTO8gZl4BtZ9BeP1s+sslqjhXgQ6Wy2vp+PtIo58Par/xQGqZTaMv14DLbXP1RirXWjEGE
UtBAulEsq3ECCj2EkREGrOMiV3TBBUkD44meMMBGUq8OflQTTLrJoC73b+q6uJxGzOUIIQcVIXjg
3dzpLt9/X3S9gNfc+wyF+IFoc4+DauZpBrbDptmMYVC0IOBEvMr/f4j+dfTeRVrHsppr2kcNaw7Q
y3i+fhsxSGz6a3KXUkryouT8YfDF2HeF4XfpK6RYCUBWxKXW2jg1G+bADULdOGesncQYr1xYvUtW
DKITtHJQtfgWBHfHU8T4jgxz2rJ+Wdzy80H2BXqlWxLvICeVrh3TQRhpVs87Od3ilhqgt8qNH/ew
shpawAf1nUkj4iOvhw6gh0kFupaYVBm5NfBX65BuOiKSGzRSrVYszWYUIfLXucOj09t1ODHznwmq
tkQtO5v++2ynr7uocKeJdyQUeol4CLTHNelPyQTKn55RaHSkSxPIVxDc0N9uQOy19Qqs3UEq1H7s
lm9i1F5OEDf/jZZGbsaIY16czVZAK296VHKGdnqS02i7EnsGFylycqK9w2QJLGosRbGrVfMplQpC
nS+I6c7lRGrxF1jW3oN5nL3I6bRVimjJRaiGD+rvrxIwlvyD7GQahTvU7X4KLGYMrqglqfAFEO+C
UXzF8XcJ8jrNvYAl4x2wo1RjelVz2cz0DG8R+bDJkQLj0dQu1x1QhIx6IE9oXCVp5wUnRStceRv5
0wdxdjtA5xsCuk6DqvpPLP1QWwAT0XdeX34/eqHBrIrNim37u3bTOIM9u1DioBqioSspkV5W+Wd3
znsk7aRXeAH2okh16p/AG2waQ7yOFFvNwVlMq+431e+tIR4AzMvMqGzgJw5X7CHGl/PewkQuPCWk
ZK1iYVHTbDnx/a18NOQ6v9qomesTdBoFLTTEX8iaTqvB8+/Hn7VwGUebKESdlcWKsojb/y6MdyWy
q6l3c1GP8T4Cpf75NQYoz9o/lohUPZKPSmwQwvOUrQUs2EkB7Nq4XB0MkcOU8+wRjPMLF8FUVYyE
xdey3WoTqd/zQazkp3yeQAFZJRC5PPpREg3Qv3spHvWSWgoOnhhT6U1HpCQqWwi+c5p1f4p7YEKw
mSpEVA008O/4YCvo8a4pf8Cr+hozy3hOKBr466Rx1hGxTPlJJhsYlEXw/FhfMWl+a367e/FvUlP8
rCFujRwdDLyNMNqIAwdFlW9/d9HLVznJoCK5LPR43xjNePcL30Qb4lOQJbZl6d+3B8rvLju6/fwu
2mL5PkdddLwnm7VUazzJFkkrIKPgxzShOC/OucIF5Lg3dtag2DDounpqnViC/AS3YZdyh8g6gaUW
4FvNMZXNEzqDLuZzYbF9wFPjO/ta6gQAvtCbRh5ibmlARr2/Oj2o7JPLTq3sbHu2rlultWypuC8c
2KZwEddfRT56rZFF9QilrkOd42U2npB8Jh1mDbSa17vtds6KFltkGUyhHSYghaj2UkL1y5pPlk5x
YSmvx/XkgTZmAnVYvAJGDV9sl7qtXk8EkObkf7ILkm+rgQLeayyRpdGtgwMMD4QUvZwTbk5rEihz
QZW5XOvoY/qQ5ABcKLqqxGOrRvNCMMCw6nNcmKOZKwUvKX/Rc54HBHQrHfScS5B2DnsfUMj0JIBU
OMGs5zIbDK6HNTwrH/wCzAPVzxSHookkwJLYXY8US4uk2ojJUFwqwFtz+WNH5oZCty+dz6aZq+11
phy9DED2GNbtgkjZA+QlavlUJicVY2UjOsHnFxYvr4vqS2h3hoxBRUHCklj9D4Q1T67BM49d+FOK
p6Nr5Uncv3sOYdECcBLjK3g3gIYKhRfY696BLXzLyMdqsW9tmKwpzH8P1hJnhdWb0uXDaX9zyjc8
sDhREM+zaFITQCX7X6iIvCV430lRMCWCl0R33W4vSxeVUxZhnqRFY53rNJCHjqd/OVfvOJ4es3vW
dTw375oPG5TV8XUzgF8HcfJWIoObZx2HlQ4P7W5J87SI7BauCLxDMSTlpa4wifDQRs2/JJj2U1kR
UhjVTB+l4oVqo9UNWIZQ035eVpBWbF7UBesandBc8ObfRBSH3WVUV84l8I80h3eEreXWTFep9k6F
F6NTBL7JGEO2UltzldoZN6MVxrw3Ht5Ca1HbdzbIcgjvh1YLNMqEFAe7zoLnPiOnUpki2RtD3scR
6xJKovZillioJMZtTNOWrBTFY6ArsvPVGsDjNzttRkGajXNNm5TVD43d1oLcwuWgx3VRgBxXuORT
kdsvudaSjiOzGtCMEi4JdqHon/cApvc2VViBLlB7Ta4P3onBbvTc2gFiScOJ/aOYTItE6kPXBZbL
x8qkcw5o+tByEEhZFyoDTQ3TxgOtDTvAdq9yOkqtrF77QrzuvEvQnfEZJxeCEvLqTdVZFcRneanj
2Htjzaro9XAtkDh5mBNABAXWdwk1DBlv1QTkJ5VUgCXGIkPlmxSRTbmSS3ouJtw68ozzyW7kI3bH
iyxMMLHd18iUNovIXLQ7N4HbIp0/KL7RQKxLYazUEAViWzuOHW5cAlk19mNP2h1WrRESXyceulxL
ETL6oFhy7YYV5L/eIfAMDeZPGTTVlUCdXYZah8geZEWcSMYYQvaiQepNubPmG4lOCuAFm9ZnFe47
UCE1h+WB/w4QQfkC2OAUcgBVqETKaUX8TOML1IcdOpPeOJQd3CgXwSsQwrEU/6dDmUdiqMVKQJeX
MjAzxZJUDiYiTvUZoq9u1zarGwaXu7nNZnSWTaRSPV3P9pO+xDaed55Ao7ILMnmuCu3zMa1wrriQ
9wYeuUq29lI6i0U6s3GZOO8WlM6VF0sWga81l2+jJ8qwD6TV43rXLMCxEe9UACoLAUpUaTNBs7dI
kJcsSKTdoBBHO24dtTv13TkW7ewTBivPDG9ToOqKw1NGKzILvQcrgsgD/m0R8e+VV5HjRRf8bFto
wmaLRaykUWxZGym+c1oj9+GKffOg6UXsse+joRNIGycCduJ8gHEarVGXua23mQ6frpJwowkox0hp
KBuz+uAWTfQJ5xgRxZGmpU83qyoj+IGXmp+PR4lrkXZGssRjoHeB4yFQe5pmLgFd6GdMe8UPy4Ku
PARfP9XBK3nAa6XOSW1OzgSy2GXSbyIrKnNTC2+2iZoLWo6hnXStDD9ZBicnnu/MBPzBGveaXeqm
B2NRWGS7r+CPIXGz0IY9Yl4NDrrZ8HIv59rNg9jWraB9TTyVTvXLSkYVIT7iflLDRmkW+QQ6FnR7
VAmYvdDL2s0Z+01JC8mxa4ly6JzfDPEs9FlIVXchoI0yKzZTt37RLiK+6u4MSyN7HEEtlsKQxnc/
h168xOxDqeai3LF3MfpVsIC/pnvYvVvaaqY93QAEuqo4KSM0APoS8TR26ERkaD/zQ8i1so4rtfC8
vqJGFKRCj+f8co90M3NnXBGDvtRDkI+d+vyrYzZ3ptQX4Qi9TWnYdODX2ibvzWN1Mk6DXKX+yYHy
qOfC39kggwHVAHuGPk41Cveq5iPVpZ9q1UQfdSMfacH2PhuSTfRRa33xDz9PZMbNr2M+6wixJlB0
+mnnHa1Y0ZW+yL5EJOEFrJ1Vm5033t5EyKFw0bts2Kg5efUGX+mQrr5IilyanrhMQqUj+BIhopgN
I5tOyau84oIHlnlp2EyhArtwwe4nrVFWAqnuYSUJRNCix06aKSo6L+y/4EfEIsSk2Xta29tbqO5X
U0u9LSnpsjtg+ybIclmuBWJhw/kv1PFBYkRCfU7VTs9oel0dWNgVSFh7t7ebiEPHZ8wpl5ZYE/ql
YV4xbksEnyxnULcj0sQZznfZ2iunuYqY0t8B0ySw5/gyuB+THb972ReR+/07rjN0nqsTgd+TTh3c
0O1HthpObb4Kj2GDBe2jIIIsehsqQr6deIwh8asM0681v6nzm0EUZfQIMqhGSxlCsFNCSlPSzxi1
mFwVmcDNBFUsjrQZvmnXc8/qT9VTbh16f5tHur+mroLpuZCEVdc/L5AXXRvWLFuF1SQKp9BxJb10
XO0hg401SI6f3LlA64i8QA5+jTaqwJ8X5vHWQD26FHDlh2s+lIt33DRl8hU5B7U9RDghP3hJmYOI
cQCksJLkYzvj9u9phX26iAB9so5kPX1W8McIdYRujohuJ6Av9sAUI5mczupErl60/BicZDsyL3OL
LkRR9eyfCdNTEWcQwkpVxKXZJMgr//SpiFtSt66GoVuKGu1pETT+iVKuLr5h/6ivDMZEbqq2QV9t
RWRVMAzR8rVNWWL7S8EJhsxQqB4pfANgbcnITJCrgpnANV29O3/UAIuK0coJz5eqZh1bc6kKI6qi
HcN1VU0PAPE3uHFoAmk7iz3BKSxtqWnhOhxEZj2/a+kXZcW2o1awsTShFd/MpcWY5yNkQ970nOLE
B+3RrUhXS4+xUnW+6w0kaeKKRaRoigCNQLHb1QBhBnXFvoTi51Nas5rfIwwIW40CAeKyeBifmxnU
0f8Piw71Qn9uKHs7I8SF3M5ivw/ELevLi2GsAQMpP5d2cho9z67O9eeCbAzyAtLdoOdr9T59fMqp
d+ihTB3wb/1mNGALsDBFX0OSH8Ypp8QhQ+dpdb+oZfhh0xKTLPpv4QO9tilgzJ3MftnNvcYIWF+P
60ktduSuZyomz1o++7rWGKE/irlH9sQSRhhxUR+oXBWiFb6N6jZXOcSxYQIFj8JrECvQNVmuZYXv
SCIlb4SVWmHJodoYtSuzrHBdF3lnHyAsnodEltMRsQvhdD7UTQQA+qGpMivX1WaA9CTVTrhVvTwu
W808XjoodJi/hIZK1Idya/3TA/id5L7gsnHSbh7q8NGC3RHnfDcW4qO0YfZS6kA0gQHQ2xaGrTSg
L50tiShFeIFBDhC9AqC0D8iudr9VfNBo9WAV8eCgmWxqcgyHOu3nhQ/hfOwqUdZ9qpU8ffX+4XvX
ytebjTKnLwKeQWlpY2jZJHSb3N7381DVq/684tycta5dzrTKeTNXHNSAz+BsKwIozXBoCjkcEjyz
iQZOrXOViUyVJgS3QSnY1Ntx0z/LEWvsU7KEe9IZ01Ww/BuXItoGvi9A/2RFbaj6L+dn8ectw45j
TGT/ww7OLT4YIbfgyFMKQKVUgZ4Zb3kXjdJPhwik5bgWVNDMreQiWPT63SVMLNi4SaAtTYZx/Q2p
nu1VZHbU8P7kG5R5iZElNSnXfj6DKECPEwAh4gXDLpZ6cgxJaJU1jZWjGuK9AVSBlm1JeoVFlea5
w+iVRMw/P/OXOoPoME30hICB4W2DV0LQLsF+E3hnjQdKkVQhFbNZ8CcewSYuZ29ymkotjKh9HulJ
qMQ2QCdYv0zZLoI1HlUlMhA4twagn2wCGd6ha5nCS6EAxBZsdcLME13TNLaW/9+u4WcC+phaFwmS
89NQzs8VifhVPJ8WqwRuFSaaKrFhYVgX9j+uQi0kesnZzuJhptM3cbPWKw+H8QG4uDRZ6X5opFH+
TNnyzq0TWlKp79cFuHFnjm/4e0oAdZGYKgEYA/m8gz453WpVR1S1gwfVFM9OeixHPfhWADgGn01v
HUG8eVc6Ll1xQjxHZaXR2tDuHy/KVyoFKgtRWYOh7h7Y1zxnzHSZJRWxiR/+WZvXOK+q8oSlKiwu
1145nEkAxFT3LL5FnQ2+NdrTFwfb2HduY6rk2sWimW8TNyk4Kij881ACdlTe5kKhjgf9w0iOnZcS
CAEH7Y+NycH+0eV47MjtTwTfkRWAKZkIoeWz3HcAm7q9M+sXJv/KMLLGCuIGZc5GxxH8bsGTjmsv
9KYwLP8TdctiIJtPgL6dHLmX77chc7gBr/PkjXXulB0AaKPqOKAfY7fP/rlg+Aw20REyrpd/T+Yt
rzA8OUnJ97qg1+MA3BMkv68DUd7ERDVGqAYLWq2kHsn3xP37hkdDrWeQI3mVIZoIWxI8O+oUkybV
rASkhRSdlQtLbP4J3Gil7+IVymrh//3jWjmin2bcaBZDDQMjcU4PAFUgK+JbkJDOgtHHwSwTXgUY
CFeAiRS8cRKax5dUHS1MgJDyklZ2TFjf5aj8PfVnoxQBEdV0v4h8lrSCNyD3X/Whj8OizbUWxRrm
YE+Y8zY2/q48vaF6uDNUHCsRW9nnKaiTCE0HQL2mzJeUfPZ54t7X2gySAKbzMaousZsbsaBd8rnS
uvWF3mcf7gvZXF6fUPQuLSydtx4Ax5kSJgme//U/6w6Zr4YbzcjXsPJYMfjfr3QEc+IIi0yFVhys
Ada69hOGHJ5ZuXAbInqPwO0Zzx6yqblYCGG+yFkDnGiPIG7IKmhCu+RsjZ/isPuYf9JNwyZvc1bk
sgg6NyHozCSl0DJgTYSlivsxo4i7SP5Vs2kmMSlFr37WyplkZSDFZDl5RdGRnDyNswtmrV9NwPNP
M1c+m1mA/JDpTp44UtTjJwlm/sxrO7ZQozTeFQLTc6x1IiML9zcOgdNqP2ndQyddvk7kWx38DNqF
9z0kwIcM3G58jFfVVqYsrKqq7xhol6gJMZBoDFqre/naMGOzPhaO1tSZIK/6CNNLuppkVfkszJEF
4dEdRBB7IKfZOnnWF3AO+dSXKH/bvo5rzrfTw1iZIlEbk3YR5s+VLhbXMhawPLWqRnGTLcawXEqi
B9YdjnPcO5brQcizB80mpzSm0goeGm3SbKUYQDr6hTZwrBngx7TG87w88nu5vAt6zJduPsoethl2
vTiVeeF+psdThWR/XSY36kqaDgeM4IYhzMpRZPk6hrL0Exi0PPlhHuV59M76IO/dF9wytlkJ42np
UZVnm2dfxvWcIf7doImNfLmixC0OL9kqNV8lLtoMWYkKeIy3mU6UVu4i3EVT7dQTdSrEyIChvKDd
ahJdA+VJoSlM8tGuKP/Y0r8seV8YAiqJ29WQO4EYj2lkszMaXhUVXPa4t2yCBfmE7bkeGep57Z2o
0h0dUL6gCKVVdYo4ZQmS9fR/fi/YjLEKZbUNKK4m2y0ipqMIqqzpPKxchCjHf4sn3jJiyGPH7hh8
lFIeeujEVZARalPcpYP8ugiqeSsmpu0S8JL7SQ5/4bs41im6kUuy99LEf1MR/FvWqAMuVTGUDobG
Tq1N3juj1NTD8UObUEI3Bz+jHp0vsZEwETvHhKXQvHEmNdQlw1jGj0o5cETH9FRLnGAbSgdMyM+1
l4uw8G50DNeE3WmT8NdFaGTzJV9F+eeHPKlrnh85mts0Eak/vupuYVGNldtOUfXJbKnk1fmXi45z
2+wcg5qgM/FuDpQ6N4xZ7yYaAdOyUo73cwBTt9rBux7Wha+hUPFKazU4TxEKCiXsZ+e/hIGFCxfC
Y8/GxyubKVT/S5NGfeYAfyNc4sfVbt/eCQCqiSartm0iG6LZq4Htw4fXBz31JPi4PBODFvwM1gt9
dtios9EvmKKPZh0HuzJYT09lDp5o/UOhYoAyMa0RO8tov3XmsVbK6HkGb74M/HCdSyfQ8Na96Qn1
pNAc/mwq4ABrYhU0lQeGdW+uq6sdhLWQlVh4cN18/odIUb0giAvexkw5OYUvjf6PC/OQy/Mpc4CK
7eWzAW0OhGP7OvSx1UC2zQ9mM/qxy7rvfvvKt7O6Iil6+K7SN77j3BbF20Dma6xRU674DzF4YYl+
ECR6MufbTxQqF4WAd7n6tRquVBmHHHHE6MalSA/md2zvMxxVumzGmc4oRxP2bN0N8TNd/QpCNF+6
6TF7dJauXVpyKJnPBGK+/RYJeHkGKoxMLQ8SKkaYV7F//SYWeeL10dt4b7uikHA/yEgq3kKva+Km
EY2XAu7ltRqOEVGGeIDOU+3yygxeuF2fiW8N+mhWG7uSEf1wQJHSvzkVyARP4TTJmASjX7gc16eq
QRNuunN0wJcCh4yhb5++kiiX4iaexyss5YyDFcoWpcY5N5Oq7EAc2q5E+a3k/yberMCBHCvCdvPJ
BIpJF5zbVUiSmtZARVKTkOiFiJ/hPb6O9CTRCL1WVGCLNbJYUEFDZRd7MTl6tz3APo1rH+cam18V
UKhTyHbhkfHXYRN/4O/7QucFIiwGAT0nkL4ok1CQ++NbyPTSKifk7QNtGliJfZKpyhbP7ytUsd13
BefpsC+UQGrxbByfpyxxxiSX42JUObVY40laU04WK/m7HwU/X2wjAJNwEzbURSMAV07maWdMkjmU
YnhEaAubpL+DQdKhByGxrEIQrLcYbQz2bfENNK9W7XPQ9kuBNr9bI9/D6QbOO1bAb0Ojgx1Gx2cY
3f35NDCHGqnWkk2TCmvSK2Fc7T0ouBcOfU17k6g33TZB2IxmJmdxLxh2G7dFnWypd53iX6Fi4DmS
vj/BpWmk5TARAoEu7tWdS/Et3IP5U/+xXMUjpbJkWhEElLQKUvpIgNTx37w17w9mpjzGqwg115s6
Xz5GFsFVSa/00G22onDZA+k4zugXS45hAcJLjjABFJV+YwyKkTjcD0OieuCxumS7vlI8xHR/o1LS
f3irrosglUYVEh+BKU6yD8IZH2XD4aQTBSUn9OmylKXdqCFZB6CXQV8lMIdNgAtErwAl3PMk0OXw
7tV4xY32PKutdXih1v4+H6xSIk1E398PDn/MAsN43lFAup9GpOiwkUpmCgVEG3NQyoIfIx7hBzBc
AoOa24UyfeTHkaq8SLuPjqyzHKnhaeKib67ovMnncQxdGFZl1z++JML8BtUB4AJlEn1BB37EmA2Y
DsbFbJ6FzMN+LC9opoeUEleELBFyFIxJWLiz7Is//8TBrBmP97LKeUJKoLcUcqPf70qR5vN5lT8L
jpyBu+k7VOj8BSYEkOlnOymidDQNhCdC6VcU4AgDT51B9JMt8yGpG80cd4TWORI/fXI1Mps4XD4P
QHl4nbvTp3nfZsx2IE0gfjAsu/S6hPiNrH38q7GpLQshz9wxHk1xSvrfFxwF3bP13CWSoSuMelzZ
VbC4wVCUh8OpSnB6E6bvceVTCHSuVQmxv1896lz56kJJnscQpMCyLcFs7qSnHYej0kGOFnEbqTFw
tvbPKuUA+ZsiTL5W50POsA0Tus1HYju5xk6cLj7otQCDk265o7rWTNroKCJUpKWNxaIx75KAbVsz
Ohlmk7Ss/NdH0YTQkhOmjqj28sSbrC4gWoaXnSlfzB00ZSukWkUexe/M/hK+HKkCK7a1xWZHu5IN
lp6PjiHooc3Rl5gWTOZDWs3mteih+sPFFAtox68jU/ycVgI33B5dU/N9BU7exeFMKs81mdjJtXHW
C6zRxJ3IIlzVEIC05mmWmi7ehsc9jdWTFSDuHEl+limP/FVnnkvtDGNWnyLYzSS7cdMZC8/QZNnp
+uH7lI8FmZjKcvuGH0y+MvsnzHmhg3KGFIlAoMTj2dlR3bO2JQgWDeHCfds+fyZpuVVaEtVVlVPp
f9+J2F+s7OruE/xiPuAujdtYhgsUaiOgQVidoumHKwKgKaI2KIuwLsLkot13NY4zJDdQMfXjcXZq
F9l3tjS3qwcssAasAB7P6wLVDE7kDuaCs/ILksTy1Li8xxSbV5wBkwRmLaNV7WOxEy7Gpb5xa6/c
zOV2vPbgW9c1jDyX5GkFkPBQGLyiFUkIR5Gq+Zke6GZnGcbKkTFEeGV7bGjRDpReGiclJK1pD4Ao
pTHREOg1pzIxIzjnBojibegF3kJeA1UIq5Zi6evyxshY11L/p+XMCRtkiIn2STgztoCLFfF9SuRN
/wy1L7Ms3ufhRd9AquICpiDOuFsEY2Uze1YFYeAenJuZgk3x48gMvkhl4wQfzl0avXb2uc5P+XIE
Ohdh27vLXqwBVBZSZPu53mFXenqqUNEgK91g+QuKXXeMNIO7dCv1o0qs5ubMKst1xZDRz0iMimY+
uiOpKICTzsqI4gH9v6pjiWKNSpryie0uRYjElPS3QjBlJO2DMtpLg1PPnBu3jViVPGEKFsH86A75
UstJc+SnZ6a1xuXbxIryKwDf9p52V7U0c6HQ2LQOIFmruYyZeRuCcFZ0g8NPyC93F4vyy8pCQnDS
2qYxjgR3Zemhv7HFa8dF4MSkJZJCt7M4VTLpZqnfvs1geX5NYdjlcWZksrRZ+1klOJ9GY9YUppG6
YPOGrj/ZgGbTl3UcJcD4OTmuBTtIRgIH3CNe2Fn7IS9R1bgwPfDpnuSYPyTV3tXcuABdTpZVEUXC
zwVyqR1cI5f5+YEyZYgDzubWoDiknmjQPw/jkJFZHSXiybAHpjkuF/hSH0exacThXPDNPcq56aPq
PED85xiaCvQFX0CbQl8m8j6xzJ7BRSpvoPL30qGviu9F/IyELcgbF0W/jOLUzgj8/F4+XeRtV3qc
/ZkdCk8cwWMfCgdmuTK0QDeJFsGcPZdiA3AfjwiLmukgeDgZjpnqFEBwLET8aiKQ48fLxpJqI6cj
xb7VDb5mCp4VBDxbdeWxd+ASs1UIXvmnX02cc//K58zpG3d2T3FHB2ZhmuqpkvgBzqVRqCpoHbGv
zJMwhRnXGmmhg04L2O84EdLQh0XHVo4Lv5f9mMUX5FHx9hK4WbBaiy4dniEBLSU0AG9DZZaWQo6I
kEwSw87iG+dPkMAL/WCNIpBVLXeY1vqdoUv+K84Bkh8FCRbj/oj4RtzSrp/mkJXonBB77JLgqHIm
svR8pCFYahSam2zJZcIxyEiQzeF4Iqv3EEXBHP9sN8zUmGIPxLv+ad8jFZrQ77rSO19uVVpgD7zg
ZkNVrJOFigTO6HuxSWG0JhUGkAhBg6ayYP0dL/wzT10mRN/nWcSLxuguL9lg5BHT5/9Mdf2qXxuY
U/Sa7beLGXZJHE+BTRInyMKgPaR7O+4S6iI4CHmrHDjEwSJ/U3Q22KErT4LBNSSvPvExzC/lN1D2
dv1LI6BpXnAtviAhDDOD61z9DoitjyE5xae65dIAFHMGLevut3khlOnlDlzcyQ5wlV/2WECnlpG0
kToi2OqQj9HT+hOGSOiw9EaNvlU0DtXXjTAmio/c7Ak54hspXQMXgukgjKLjz1+M6A1ZMPYzs/L8
+/wgUAhkJY6BqofvnvFqQLo/eQhLXFCJJuBvjDxjAQGJRsGK8/uWqvXXkrT6sCr+Oc4TdgPPMyQK
rE3vRmNMz0Z/VgrW+gRQAnj5IU4GZ6vGVt+VXnoer64EkUa0XMgoj5sxHEuI24A4N3phGpcOtZ/R
W+cVAEMV7Zbbih6hOVj/2+OcMntT2LbpDGoIlEDhZhmzUAk1SSISCaeT0lL73GI3qbXW9gH5QpZZ
ySZIuwzqjJxv8sZuPNpt6ezQlCJSGc9lnzn690AOPL92jS10BFHr2o6AoxzF63LudKkf5DpWzgJV
7JArXh6Re4jowKyQlHdy6ygElusUS8NrW7x7pPE+uzLIKW4tX7oKHKWfNRaQErXhr+H3jO7vO9oW
na65Z7298fsW25dnh/RYFteBJG/O93m5tkcHHNHu9DRFAmUfQz3liGgg91Qyqj+1GntSR1HqctRB
Doko/rrPAZ+7KE77MYClFFrysNEwbz0GyhKBe2u4Im/vgDfvIHPi0LoRsrhS5tuEqK0Llms41lTK
vMOp8cpE3dBLifGX669noOzvXSTU6Tll+oGXNAmVGaFhbK7ycrXifwOHgypVoR4i9atMv6mDMPbX
opcDRwpDHdkOe/Nr119rUzjUixpoBZnXAN7Fas9gbJwtFvQvnQx7sor4E2fjfm+lF6QqwPelEWf9
P+magBlOuEEVXzmr2dZHxfnwKg8TLiohQCVuEXZ6/R+6Sm4hDW5m8/pfPiDa9SQEuSM0bZp6aLup
YRMxejv4IfHW3y3ljMjaUNkGjUApI0GXFfuuR0o9hPUlUiqrTTb0+zy977dDkpZo+JuZDLIBTF0T
yyFTbhh9eil1cfmPe0GTKhMwlqz1bv2/+bzeNXJmTILSbBk5Y8TKWqM6BI3c1y5kqXWYNRlA7voe
JlavVXenTdMmEqn8xfy1tLt2ZXOILN8sFWu0DQQioR9yodMlrEaaZGtxi/WGVYndLz04cL37zCoK
adVMCwq616EUW1qwCLb/MnH8KtT0T8tMwWbTClzYOMWbyfsOqYDz7JhRjFkqr0rkUV15IJG8BZEx
JyoLn0hTf6rRE6ny5pEpODdCSR9DXCiHpN5xIg17yO9KrZP2+lxr9gyHKXH0tQQLZuxZJy7O95R2
zt6aGH8DPK0QAlw/EmVRyFbO/t41fKm29/XrMcesA7muJmVb7v/1VI2fwSsaA8m3fKrRpUOwsaC0
wLohCGwsyL8uZr3fuTirvV5SgiulrXNl/g7HaCDDbbDCzVDIjcxVxmJ12HcMpxmzYphFtuXv00Vz
gu1g6Dv+LkWcYRPtpDg0EjM9UZzJE15qQs78p5n5Xim/RyeGi0dVr/02BVmaRMpztXacHZwDwRXw
RoGlLUT8mz32mS9yaKoP3YYA4Qcq4Tu+bIcwQsdcG7ksO6B8e3Jo7l6ux9ifbQoXC5cnoNG3qOgS
ShYaRzLzv2OXLvII4vsZd4OjstcnTGGzv3oMTc6azttp+ALDY6+Qz4SDLXjIrxBQml2Dmr6om2m9
4fWSbghpx/T4yDPPbDaiZGvUUdwgx5MkhVaCvh5wfxoHYXS7Dnl4/1BxB3nUoH7wSrIdsWtONOgZ
bpD+xPGUC08ngv7Dj7Ml7cHazeUoCyw6+LEDhgi9BS1GnJobceXTnOnsckFzwAsFDI68XXMREny0
66g+5jFVgGzVyz/JNFKAJiQN87HG2sM651GpNoKZGW+ry0DXTVNFoWha40v9mspvj/dl1PR/oEqV
YXBT1r6G4ZV6fg+O0SDg4q1B9LoJiPnxzdmljHw/U7HboNNuTzq+Z0WEUf+GpFDvUSZDhp4bLJzr
mF+/uwD3Tem5qbQTnjZy3lYhEu4fBRVsOIdenug9VKEeGnDdpiDKXK8Bk4ngFXw/bCmyteDLD+sQ
4K4wOs4LCHIsOXVP/A+gGPpyISadCH8JSzCphmeD5xbl0pDIChsBaVBdY84OYIVG01QrSK0YuVx0
Lytxzw91WYg4i4kdzGVPastdqlfq4wNnz+iLmVlgfZeNceXlhootQ6r/ZvWJ0hC1khSloY2Fr5B1
XreBrjajRRBeI8Y1riceIJMdP84JjP5hs5UPdujn2FF2e98lhSJplUF/r9XsMQm8Vc3GZGNxVzYc
XTAHLCRxGZUQDE160Qrd/rczYBRhJgRWRWCahLDapUGeNcDvnvgds21CHqaTS9JABuvpc2/WUTvF
O/fgV6etlVPrcSaD2oOsyvJND/PcRgdcKiLNX5dVSKfHL1SWYP3hEXvI+z0B+/Dni6fJldWxfEe/
2/2sGPJbCQkm6uURYI0CJpZ4/DkpO+Svk9bpKejwS8EQTAPaM8wrtTW78md7g7znIXzrUWVj71lT
E48+s4jSdawnyMjHUvSjprdXmrmLeX/4FBnUS7zowZZZAHDbYEHPJi7he9m2qe9stAeLqdR10Igj
+v1zhK9hYV3laiKsdUKtv6nX4RstmwrT3K4aO4AKLS/l2k9aE0UZ87q9KlCrPJSESKeWoQfz/iSn
oFQ1hsQQ+36Uy8gMegrq+GByc7BSxguMYx3vBH+CpuK2DOFA8SA9j67SzFlI4uiGTvBhj5GaWWTB
N4g0FVEzQfA+R51dEdqAM5UafHZgPmDOsPVPUIRAsTUHWzpmGO98Xxf7tB8whAgHBFadbmBLUfhC
VAYbOlXPAmz5HLqgSV682+mDwKviudNws0v417WgWAJyckKVzdTsIC7WdO1k6i62NRSqrQeiePyA
V8XH48IfPCQAet7EO2/BXK+hKvC3bt3h7qyGFpmM1a+SOSmr+yZ8gmz3F9GLnd90mBu48+FzlCuc
QFv3iTyEC1sO2RfUZYFzQ7Lw/P+Oa30aikKsCPIJbOa69uJdQx/akQRfGuV21aq9Rfrqnw8OgB7B
LUP1zIPdaQOsDPOrpHM8vG5xtLN29K9plBuc0EHZSh+hcYZ/m+4Adble7oiqdk2YaVi/nMdoF/RD
NeE52FCLxj0iZPGr9TsdiH2VPOQ1AdeJWdAKlzYIzbBWU6y2rjq001rzwnZ6vYP+a1BK9rjp/J4j
ig8EZu5dg70wwKQECpvr+nxq8s3cVLaEmTn//FYJUGxfb1o8INrxAM7rvdB3s3xxwZLGFdCYZIlB
VVun9aFP/1JLl7qSx8A5sjxwSexkTJkU38/reAHaEu56LkC1zr5m6BGKjsRghfg5HI6FJOsz7J5g
NDmjfvK8UVBUCRuiY1FTh/9aK+Jb+UfCTxtSJybRNy/jciBEPabM1+J3gWHKizNsM6VxekoCMXvJ
8XfAsAshwD6t8VLtuQK5zLE5cSNGnu87gs1cHmcmg3gaziZ4uWOAyCJ4c90hHHOPrmdrADmh36v/
9mZFTCZoCj+vly6Eh1dMTH34iUMHNhnvlKPZZZT+1i3PlckLLGh+gEXQVQjam4eXdNnsYClNIKHh
+UBs+DkRflQCWVdRSnje33vQb0X4iCsJX4mOBxwLpX9DlMVGZ+1tUxS0NwBFo0DHd5kMYOuNgxLG
8NBHHtTjIuUPn7yJwD4JBp6zVCY7/O5CR6q2M0Uqcly/Ls66N1HEyJT96bCydZZ4tYrDyTiCMvqt
jniRF+1IYF8qearrwkdXlQplYn5wvegYJ2+huw1y2+Hw7AYTJNWqutLI4VwkD598vkicM4n2QH7S
jV/7rzUuN/RzorGS9V9VTxlXVDO9SRFL+YFsD2B+RVk9UydPC4lA3fFdJFScinK7ITq5CYoTcvCD
KPDBZ9hbfp4wAM5GN59b98n7nnmZgSXTH/IPxPxHHi+GNdEoemv7xUh1s6WomwpkaUO8PDJNRKht
QOEjQNGHb7VPH4l1phhAZrSHwoIHH97Lw9W59Q+PDjixVahQyiv+8hb8KABXt69MezTb1C/Ca48w
VuW8zcfEkJoqqg8pdKeDiw+udvGQunN0bZt+I8G+e+3f4Y24vC62EzKAcpZJDNG9FIs2FQgaxiXD
W8zESteN/ZHICugyK67PjULrrKBE/WcmeUrMFQR/3TKD+kot85y2ta+kGkBkskz414y/3hT4Errv
48YEDJBkRNLHmxkUlJfFwDH/lLKDry7WSzg69HZQL5k8WXBMzLPAUSM2K+TmsW/6wBx23mMvIKnx
SB4mR8rvoMELyN7mGManRgonFaJWBs/l2BInZDUuiH0jSMkL8++dNDAXsYhQ9gWfjD28R7/qO4n1
U2PJC3Oji7z36FnyAtT3pQe/Y1YXA3KcK2qRPxU8iNz+d+/jv+5VrqE30rIL5FqIkZycTon9lYlk
ATEJzXJ5WuJtT+qTSHzu5N11SO3/0rfpDw9cfysYHIr+7nCWxU88qHkP1tdwLDD8CRegVzWEq+Hj
kDSE5VwsDtFRLO3mAsKiM6Gch6+u1IU1O4bqeqf0Ff5L+X5ksTHF5MOBQpCgW57qW8B6Z0ZeEdE1
nMmYUKswCoLnZQMYrbl2EbuZqA4vrmP/xgDkJ8BDOzL9sp0OHC5NPfiOY108WQb+qGRm7iHwOz6x
2fizcW5eb/6FqyjdEv4v22Hyk6QRnV86wmlHl1GektN7DQ+DsfnHrzZU4/LRtf54/vZh+cWfxDm7
+LUVCVaUF3eu9bOH06U4U4DIKsCno02yoZBZRflHIFAqevN/AkKsY9ntalYAiZEQryfFD8XyHs24
5lEVkrcw+TkGIh+uXxywJ1WscQErGeQipCQLy9vYmd0jEknRYdghFDtWmuO1yRbqyHfdzinWN9E2
iAoZWhIATbTpdu9+GM4wKB/7rHDkwmoEbWPq/gPNPfGdNo4LMrVe/sBAiM0h+9+pl395plIVHmmH
k/d5n6J8HDS26K1IjdCn3jDuosTndqX1ZxX9kY3KHGNUeo0kHDrI2gbg1OKExMlr/1e2AA/PAUL+
k14AmAcvFEF5bnF4J8E9QaifO0D9rCNuGR6WpHzq1fGBIpcGAFW+IgnNYiPXn9mDD7cn8BWXyAMP
8Y52VCuF7qE4NqTMwObCVQDyRr9Ez98z1R58ScfYyuSYOEjaDGAdlTGHiGkq/yZYfPrcGmYltQru
Tm+mFK2jMhCd9LcsPxx2FqigrAYSsCJhdTEREZl7XcJDB7ulaWIMu64otxWcaHX50iF2OjYds7Yd
H2ChpEzk7pKbAwG/cV/W1HWi4yPrEjH0ljPZmb2ioqXO16y7Jy/vEtRaSWUN5EmAur5YKJn380p+
gAaAGjUng56nz0Skkqbx/lL1yCIopA0zFMC/LT9860wxodm4x4zDR4SZHz+cpzQ+umU+bkoprEu9
wpYl6VAI3d/SzZAWrrP3HzPCkPiG6IJkTzJcq5LC2wn9Ysw+DSBH8ZJUr4oKuj0wU05KzsahgKfy
xY57xNvCAClCLJjJwCui/Iz6CdkTqLaon9YRiAzA+4xrydl4SViycEODOUePylOC060wdPah28Pa
RaVf6w8lviaBP4Z2XAFgXvB8pLeKren4xFfP04IvbN2SXkwTkRNJGtqlOSfeboxN7VoHImUCTgYy
KtX4XESebtJx9sWc3nlCHKZhUmHyZG5AwbyafLKa0HiwaxaxXyUIjavYMevkUfSAmAnen/kg0yXG
Yb2U3HEoEh8fGSOSIcgt9zRRKX5pf+jCwBB9BHt0WzQYoiGVjANTEIx9NaiEJaIzOgV0IOoxsHXQ
IBMvDVNRpzQVnzRksIn+ARFGNH/vo6124RfLUkxcH6dQu2wN/N7pVThJybjtbNh2a6I3Slr65WUV
yPOow6NdAVN2mXRUaqo0k/AH2/+C4ErJBlE+Ve23iMLslE0Qmac02zZsS+fAT060I3FPvYzQTays
6gHA+1ItcIjAwDh9+UzyNbFWx/8POFX00otC6yBqcMRqS+EOGL2pkaFNUnt3+4Gp9I+D7cOdM3D2
/dETkW1SZQ9xTCYWnW0lOorxhD7cYrAcKHkmdCVtKOggif2VsaaRie9DWNuOcvMrZdOlllQ7WH/k
QrDyDnl5mp8ZC/Q/pSUGIFLUsOSRvGCO1uNWqEjjLt/eBLTtwpUshAlk0B8ry/J89y1cBWXkVHU5
qcpBA4TLlIqWLvij/wku99VM1HMJ1AsW1pu0L3H28j9Zw4RTrZJiRKYgYWVnqP5DVGPypQgey577
QC9npe75j+CerRjZwr+yyiFjWC6kNeIieiqLZFz14YUCaPzB+ocwjow9al0qs6ukznNWtMIVQZR1
YM6CgTw/F7gZeKkoLKT+n4SztDW2DLjs2Rfxfxyh8D4AgfueUa+lUjB9697G680hyf4rvwyEhZEj
O8rT0j38Eghlskd85gRnMaiMCPPfd7BzDsHd0cBUBYVwCS7NJIUmr4Dd9pj0nBV384k92+qnSDws
LgiXwdeOQwgXB0535bp0+bI5HoXhbIfurGXkziwIeWrbvtjg6iG3B0qz30lUxLKp3ywrmB5FIQcf
K644QX24MamleR9UXUQ9vRGWrPTRPT0Z4MsFP1X6wZIBkkvwjHl4odIQboOgywjImRlTVE9xiS5S
F07qk7QdanwOB31aGFRrunurtUmVWBdCEjdmPQTWss80JP2+691twrXqnBSFSKFdmc5uI1HkqtpW
QZoJB9LOYsElaky/wm+Pw1uPCa9or3dXhHie0WO2/2fgLqFmRpylvEkydQUeqRfJkYzGWxrU7WGT
0Vw68XUEGSv28jP1fY4s0uI9nTfUJaB4FsQz8EHG7NpMfTk6GBBLyj6Bh5p5xIoWTpXftMoimohK
GKemk07IQq4V4rl0WkLBCQnwlZCeyXDkMWWwVc6yvNbAFvNrpdNH64G8gFUbAgPvXQc2llHjSSJj
PCfzYSHd98B+6drdjl784TrRKaL6w89Rmptl09WVFzxZQ5Gtc0UcoPeIkhwLXXuDh2RIhxMoXkIW
Cq1k6YA7X7Bib2nd9ZRJhEdJ0N8ctSLw4EyIvQlwfxKjXiHrcXjCY884lrtvMkmOz56LEYkwBtf7
wzQlFgeDJAdFhun+TsSWWB7XR/4l0CdebLVD07l3SU/oZ8K3JZoe1BJWbyEZfTzT54bJSG48dlPI
3JngpuETdvZsOnGMNMn39e9JznedgoylN/nAjZZWLKfOxZh6Uba5Ad9zmE3PXCAwa1fbwQf1Tam4
b5ovRwLj1zvLwsvzAq+TunzIXvuehswznxtykrNrEcJps0TkrQSIwvABLl/RvX6MSFf1+m+FIEtI
1rKVrnOc4nNW2mn38BZ445FXjDvxEJzP2u4NUsj1VSmlDIRZz1y6dIY7tX0g1z1RUqOy5fdUasrT
PMgfFHPkuEVj+x7/5kYHXu8J1F39vc13nmFK09ntq/ub3VKx1JmHSUeNkLur2o/I0C3cxYJM55FL
xRgGsRw0CiKzsREfAvwssYCRvt3aB0RrA9Mz7PHP5svVpovNUqZSy8PLCGgAM3oDQTQQ0eFcr57y
GG135fYxtSicdidfI9EsDY/7ZwVVC5RS8HZ+NZlMYkM5QJEfxeR/1ne1824PXSHAttCFiaqOZWKt
nDsGEa15wKujndEc4ZgQYGukwgR8aTlANr0jRCNhpWNQrIU6c6tlIihqYfflMBZ9an+3nFgS+VEK
TsO9WEMlhGMuMIUNio/47CmvKg4rwuDrvIuZ5KUA5yhqQCv+LsxxK+WNVdo0QLjfS09k5mbNtcjH
FDezF0G9VtEoRI10PzkzDTXRsGxdd44NdtewKO4XdiHQVmOWXggUYJm4yB8ocscphTmWnBpyrIHO
0g4sQaigqaZXJ+nUsFOZxCT1IlNnsxAADh0AZoe0Hozv9PLBSJxi8I36iRL6FKDSHbauE4cRIMlq
WAku4ij3+4GGYCFTns+RjWb6q5U7eqgeeN8kicBoYEpyFIg5b8JukxvCWS7X8Rq6mNbPHfdt30Hm
enA4w1jwFTs7vrOEscjobFNpoYOuWMfDXjijfLjWgoTLsEyDYCgK+PbJaYcsFvsc2u8jXN7yxGm2
rsziJZKqqiWJIWDI1exYDZO+2QsYZ4FqVKt8faRuLwr5vvCsf5bpzf8WIzXdgHqYk3NLkeXJWHXy
7QLYNPFbCWem/7AjwTHuJPsBfj+9Txy/H4C+QkRQi99QiXcmKHl23opYtHcyIoC/Qd7RANhaoyj3
O/iW+qenXu9uC1N26Nf8UHD95Rn02WYSHtNuxHIgEtmPBYV5+KaiZFMXHJElPbdx5AaShV0ik+45
6mp0eNREPnaRoA+Q5rvjPY4UExkJY+n5W1qaFmV8u9evQrOxr1pN5B9sxyFDT21y1m2aeuICkNUA
8ikaBoTcRpRY9z4E52yaStHTZ+KI/xOgbiny3pYSQ1XKFGCP45LEMNdvtJbs1X+1xxnadhuTabGM
q+XBaccqpqrjqiZeDaTuA3ykbNSpBoFr523uILDRCU8LO8Nlb4hrXodIwsMMEP5QdGh8Gc2u3vIV
OG9NDgu+iPQmv1yF+pI3uD6PvDNcEXnMsB9TNa5lN1G74qK+/gtSwZF5JlVPQMnJqZI/IPXPsIEC
1+fVG5TVjrKaGOZOUnthGfEoJPuA667aufMXdkSpeCzWrsDuDRbs07YKT2XeBeNoRoEXfp2MpDwL
aVv6d8vNyi1g9NbMrgtnhO/3S4KPMRuymHQrBzD3R5XjycfuasH5nczQHBnLV7ORGj6gQYkxmEPs
3VPcWuV2wjjPtdwk+cRuChQmLAzf34a7ZAY6fEdwcdulTlB03KznJd506pYWQJ3JIoVbAMBB9Xt5
e6buDs45fozmfnuC6BUZX9aMRjospLe+cNffnlUakYkZnp18nrVLLhiotYgt70VatRNIdJje3OQh
KwOS3fXfwYVckhVKUU9iaMYqzQ2wumIHd2xCJr0gppYMggjNlV4YPxfKdL4A6geZL7sHYJ3WMKZp
4BqfIyfCuBdVZ2oAWQB+YmlNIJ46JipfkKsVPIhV5+94HL6gSBRrUWs97Sos9hMvD8kxaSyqkwnR
7JF4TaKfT+IL5PtYMRkYQB/Z5pJ6ZYPEWQkUYodiaOCBiHBTrGmBf0fbZz+ZRS0AjSdcj201HmTB
s1t53us70UaK3BsaHmbwoliW9tGlFhRwJhAxVlupMfQ6mtjUXfbXlNDzjf3OxT9BiUC73SbKGoqT
vtVKb6WSyxZ/u6sqR9zGOx4hwmp2nQv/JJdRE72qSQ9I/SGDXTs1IlwvJNajVvgeJsOB87i++l9p
NGUYPzPXNDM2nf7U119JvLjMZEQ/nl6CUV8mjv7tbqmLH4neykONoPvwCmDgDLLfmOYwLUw+RXnR
nhZ+6thSRmbIlu+HNxMhQQk037VVZXvq4EBbUQWRBKSkH1NwsZuL4NecySUgMWSh1rQY0/0GEEve
/1UErA1sDkzvVnVdoK2r5E138fLnM0RQEE0eY2kgEdoGCMCpzukzv0GFJ2N5CEPW/Djg3iv4pqPr
o2p/JpfWiSf2enXbdM+QzxazSuhwMwPr0UWyint15vT5gSguOG9EgbhJ/hDH21kg8mYawWRGHN1+
glN7wJDinErGSx1wmHYQbCwnxwQUD+xmOihy/7KoB3eGXSWNmEddz6lEw4bxJR4ZtuoL51vYOfNs
j1UWQTfv90wgF9YWceT9n1YXQENGC0RJF4vJ2TnUjImrpQhFTKDoTStaQ2drUvtVFi+/fqCBtTIO
6X2l2JRF2s/Muxf2jxggtE8AxIVQ1nchoEihA0VmN61K1ITuYrvxCgGchys2hyskZv9r4YfGvGfY
83U1TIhkRFTg1yemHJSy/ZgSaGtJa+4qBgpZnFTsAipgpH4j3Ymu7+aVAlOLuBCC+UR9mWYxrm3L
EuG4K2lBtoBg+2ghpoCQgKwX+TiSzqh15E7+EjnpU5hc2XquravhnylmlDLrgp39nOSCl8BaKm3A
Hn+gOJ/Apdo2TqcabSmzjZKD4yejV7gyM1imSzx40eCL5TsWpC9lpuByibP9JQIZDfhzqJg1XlJd
TvS6LGdynLSo5QdNZv4/abnb/DKRXGeztP0qoDE54CAVtKvmJcaY23BIFP2SmN0Xb0NE3srSed1l
Bv2uopLLwtO2P/KnkPshn5spHFisEyRQfM7l3RE/ZR1jycH8i0HTTw8IQIoCT6nIAEFsl/7O5d53
BrSWwJg10LzK1OBrGKOpeFfFXqq2W+cuSl4/TEUWs5VcbkMxfwGDk0iUAGZNvevZtZFxI854J+AW
ESZOCsypBN+1jji3DhUQiktKkdTXkAEOkd1rCDg4XmCzRcKinGQ5sghxR8xkswix1NyRjVQsw7Ug
1az+185eTWuuYY8npj4gcGUzwy08wX2P6AMMSgVV9XTgfI6qAzHnW/orzXM1qK0lqEozzBNQl/VK
3mpK5GDbQmh3LL2cKCiDUrY6qQoe8mQ+guw6YmH+qIMdvW0EphTJ0Q22i2QCl8mp88VeF4QAgVhr
/VUMi5s7gO/1BmVda8l3I8oGLox8WMMjjepoFdVo+2airbzvqR2IrLFxKKimKWnzqIQ0TcalZKVw
ePqQjBzGjxavwKMj9Ei2jbJL/BunM3lz9I0iZgwqxPjplEP8FHVoI5dZuf7Nj+OlYL77suQw3Lnm
3v+cDvbtHjiVhym/N1OKQ8uSbISuCru9qGCLW4IKAuMar3LbfsJJu+Rak5x/m+m92dBdp6nPqrO+
FR/CAFrNCKx+FAYKYGC7SvOMdJwLvVF6U1WGJO5zrL4bd5iZNxpW/Ev24NaL3h/MEf/i0wVqt0Qx
6HVWPLzW7JzO46XYYdifHxDGHtPnSZpOul0uJmgoLYKMU4K++6AynZ3q7KibAvAjLB+1UG9nW2/n
dYpjpTbkl7KnWf+fcwYcn2aTKfGgFRoBQNMLkpB5Po+tvwVU6Ufs3Gjqy3RHPeoeouokxd+KPLbg
7O3QgYZXYkMm1aV8jrbgK1ZOqg3wpmn+CO7mMg/5g7HY+AKQEwGb98UM72DJLrxmUBjSDbOx3MvZ
4MRqdttMg3pJY0atF07Iwjzl9l+dggv4F863Jq6uunA4fv0umIU0jSD5P85/JjRcskrIcbbCjzxT
d89YcjzY8oAddrw5i/kJQyVRZGCNvCM8Npj17Y1pU/hHMgsUaaiRtSuD2crfMIeHVtPrjzmJXvz/
IM16pTN4sAb1fcUOe2cXASRxDRi6QgQSNL8p0yFRM+OC0BKI1gQxTqCToJTb5K6DHUSp7mApS90i
TJefwxz55mg3DNwqa9d1d9ZY+8MjSIPmRrMJ6ZpLZAI51A9XY7voMvsyCMCE++DrjRG1e9j/Rmun
zyiQwGZOJHRt3FknJ2JmhuKrXZf5s8vrQw3ciyKmM64y9Q0ANHqN5yDs8fX5ylWDUAwm+lcP8yNX
E5aWvyMFWXDhuehra+jlEBsCjjCGKoXObzbM8rfBzxLzSuRm539kGPBBiXXOOgpy4PtGG2cpX1rd
FPbWGZ5dI476kZKV8U2drh/q041nCAK1vN5IvmbodS2cYZmwG7WssfrmZKedsWvbUMjwTwCM73XS
t/tFHs4kQ0vHckH9kJEgW0DrZoZ3trxlrGBuAQq55Z5gJfY1EaNyqnPO3nWvPiN/N5XCsxqn06Nv
nnOha9AgrFsQwZqSqN0iK+rXBGdUucjxcCoG0eczSw3eXEaU0yLJL+cHWAl2PuYv5f+N7GmMUPKO
/2UXMwDnzpHCRyRvn7K8GdiRlk69G025tD081sTgxfaGoZGYzWV5uK011bLEYnx0q8P6gc302EXW
U9Tk+zihtU2gVVT+xg+co7CGIL8cJvEzNwOow3vnOJUpThuAZ3aHV1EHFGxRR6cqkTNIFNHasJve
iEKK8G58Vm6/gU/ppmw9yaC2cN6xysJQWosxUAvZbk+WypUk+yX9WYhdCwGnVohxclPkra5XCu+/
mIzmukKxqTRjmbn1wbSEiCOz0tbfeSoQorIpfiOYvtMOmadS7TF0Y4ZrLhQwC7bJZNvLoe6KY/XH
rwTqh5tfbUV77o1sYxissZG9inGNC+S6Heg1uBjaa1c+SKOI+ed08BVJhv80eNWiFn6sVQMAvwCu
2FZ2MJhuSrjw5tQQVoLFMFYREkYLhW3SS56sQk7YnJhQznCo1iMXkjDaouhkNuVeSyTRllsxq96O
ImN8ETzofyn2ZtpL5Vgy5nF54UJXopirgLYG6g5BAY264g3Kz7oKkmvW4wSzGtMMp9O0Y4g764e0
3dae4XSfFciqlJBicY/xfA9K/z9qyyMjPJWqn7rpub7NSWZVezllenrR0THSTO5U/gskAhXJ8jNX
wZdb1XniTm82iAx8pHX2YMlHWTYd46iB3LHdOaUo/rwPC+BOUKmz8BLtIBPDuknW7akrScXjJ78h
y6MqFBzDPg9C1ZjUu0E8jhMCAbBNZH/j0JsQPjqM1F5Cd02lpnSLUUTpcS6GscQtSulncM9kp0lZ
gVh/M2saRoIvx9GYsUoOCKNzgCQuNVRZOoaEf6laI/8Hdcu6w9usRaVvx6fTNzVkMB1Y5FV3nXU7
sCUcJY0J4N/HgtNZRYcwIS4q8dk+fr/So44TzWzou0pCOcGVNOOBL2ULZbDykdI/iFejhX3CdixQ
jABCCo3aHKPh8ZO6uUyoc6BtAL2FhD9Y+LAOLO13+4r00xiGM5D3AoWb8aA4V8vBshdqnW9lNpif
4a8ut3916RJJ63XwsnlJIze+zfXCPZ2fhnwhzDCzUz8xE+fo1keqLEn4RwRboNVaNMez6ceBjOkv
hJx/r6KepWJk9Yv+zIxROvxEtRvydIQ8cSsrTDU8A3ABYoc0D2WoSxO+wcE/0X7gLnJwtTnaenrq
n5NFJrWd/5VE8DHchdqruQZfIPzRWdjcGHxHZW1p8ooZCpKrMTSphGm+yGabTvI5XlXsPdI2cOtC
f9rhFfSmUaQV1U0WOH7H8gWfbue4jZRJW7F/EtQ2vagcuol5Mo5mGtRNgrXCJ+IHeQRKmw/XzuMS
psdOJ723CRBKJlG+tAUdyjEiYaIs4c5rmcMmKvrVLTdIK6UivflpbwYPdMb42o+DWoq8emYHVC6D
493LbVdwPV7Sxm71aFXkZRfdCIIDmS74AAEKib23YUUt7Hmp3v5+MhOqOL4CsNvs69E3RgRhfdDm
wYtx1fEnGXACkkKnvtyXaIZrQHQ/ab9DwUwz6FcLiSsgH0ZkbB7FDUGZFzn2pidhfBMru3Qq4zw5
ZPiSxZpDMuxn0CGNJqWa2RU0nS25vytS/UxYLIDgk3uxafrZC7Y1ZdRMi7gLG65VJu6ZWp9WfILm
AX2ixU288KV4OrvGlrLbM5ch/1H6puetielb936ltqSIVy6WkmnjbkLnJbqzjzzPJnJDaOD7r675
jaaUJ31z7Bam3/XFS7YdU06g3MdER16B1vm0mivk568BbSbkqNHyglqOBFKqBZYLzbG3WA5GyFAB
jQ5V2E8Wkz5FmEhsEtomh2xrBTn4V7RSiiE+ssWU6/24uRSPtkVkf8ZW+NwDELD+m1PF8sE43afn
U6W6N/hy1MPlW0Ddg2BiDXM6Ly1Rdm4hqygVE0ge8tHpeAJ2ixpTWCRWkGF2q9gfwwAgmD9p/cl+
d7/Gsss4cV1/7OrqFDn6cJ48lfMac1kes9VmMkerA9mwiziTUN0fVpfr+KHkNP5ZNw/76Rj2pban
mo8pW4Muqskts6waLYpu0LyCh0RryP1zkWwH6pzgtTIaZAiIcpg/g6P4H5jtZVsL0YuuNceWoWRd
PN3tdZk4ZDfPuDptjt7RiH5vchrdZz4gRa6ucngyQKxNc69NyyErE5GBc6uQ3/y6zOVVtdlglBMn
6MqUxpDFhKXcJmpohIXGjUwJvJfCOaK1s3WQRRG2n02W5AG/lKFMwWetEuPyRkFcPFAdvF7hRiBR
awLYSU8vQWMC+NjvuqaiDAmKyP2bI7ekPWiY7wp5DKHR7CHpLhOkiwrhZBR/VneGR9WSFElALcm8
N9e+qgIf8nhs2JQg71APbw+SKeSLfTqm0W5I27jmEuRu2V2NUdfpTVMGNph6X4pSVApRd/4a4YMy
6pFz/EqBABK+R8Z0Z2genwYyF+herkmqU50T+gly9VVExPQCbyZXznrgRtbbZUxqt+JxRksUdoHP
jEYmUo3voHddaoDqxeUW4d0GZ2v4VQovvLOT9WomVRu4RLDC3HuHvyGF/87UHzSjC+wispg8qTn6
K7RYaxdCrLdSN3S1cby+GtsMSi9g3XSHwmpCYOrUhzbBx+3MHuSA0MlDUK5EHr2AENhpKmTfA4nL
I/KTIOvBAk8yiT//PQQTd8KUk+h73KSmnYTX5U0k9dU3LpdcCYuv7N+9yshBGNT5yATGwldxN8sy
DkSHRrmyCMp8Gxt3dy/u1l9WBmMWIpFjjEzGiCG07ktDb/ta7yn4iDv+Xa8/Ih6uC6yQArq3vh07
fzWVNI0ciqpMp+FzAAwwbI6W3scrJOZAugmBxTjPBZ5O+4MxWA11xjBS7DA0RvU+e4Hq35FAP70o
JqPvblHali1U8D18+tPMOwtvUzW5hWFHO1vKhqPkPcyexwNTqqYYi2USi1/ps2qW/l6rTOJHTC8p
0rW2BiWh8bWjBakJo1gPy/KTP+2cExpmphwbXpBUimiRD2V8/eqZMgLO+p2kFEej46AJs5pQSOm/
AVwy8vA3LPJvU8R7z6p1smS565UTUikJPZadJ4K+V01OaCkk+D7+QuhjrAGOdLtrSz9RtokOnVf9
jyA1VtXlm5trTDsjlIx8SFnBNFrq4PZ86D+YqkUpU9UDsiIYAiPU1RgzjGjHeYZmUdtpSdP+BwVK
5nKNzsAlZU2WBTzbGaAT/oDWWTagOVS8t7mCnb/h5w3y1rKMMxjiElBFM1kkeaGQ9lHtGskHbzrX
vW2GQJpVs7LzUpb6npOwA0QnR23O2OkrgZRKoI4HyyEI1jis1iw8wFKcsxW19F8/AH8dA7xOGrIi
xL2iNnXMUGVpx9uOlDaKMsYhFmkr8IWg73aQNTpln/w4/ueJXCQcY/TGQTTkCwdCiEtDChiFVpVF
re6ZIDb4N85D9BvcbaXUh2kgykoa+dW+m3/QpYCinvZfZx4QaeVzACZiTxt07F//vL2E/7FPTZkT
97EnX1o4GQJI0jgStsCtn5y1bOtv78WQn6ghYg8fDVJ+BvHm0C46M3NH0jrg+kdzWRdVcR65AiTi
8G0OKBeTJqnJkj1CcGyv5s32PNKLXn3F36zTip+XGvRxevmySY4Z8JHi793GUVRpVYMXPLFBa6Oo
61fZNFvI8WmcY0Y+8jwZN9+meE9Zi+kDq+ehon8rtzmfg0efgNbbmnfvUc4tw/qgjR4c7sH2sRk1
BtsyyoIl7folhAvGgKGztlHtZpCQo1tBsXMK8lhGV3OxkeuTUOlkjfSIo6vbMscryMB+mLn5K7L0
sWuO07HRjbatb6xmn/lbOe3i265wyDDbSCkGD0JeR3fM0i77lrBpf92k8Za3//lf9mgj4rXl2P4x
f8eflwP7XBupXGH28z8Lyk2Fvp3h+WVoshnFnT4VKEl/5Skt+3luGzSjOKwZKWuEPhaui8tLPSN3
ElTNxeiyO0Ob40uQMEbWRioltR8lRSUV3WxysaJ62ffZfpf+Awqq2Q66r601UXTbHzPR7W07+WWZ
UrATJXd96KYVmdwzfQuyc2c6O9W2CdCt6jFzW+kVJ6IulQNE5AuXy6f9uxKPYgeX1ryUGaCByEI4
EYnQN5MWnjP8Gw5xtEeAdEvDPwLxyGt71rNOUxMeLydRMqz0JirOXR0n9EYs+J9kCCVrgOFUxqiR
NrwdknWUhRKzQZfjE8D1C9XIvQEZ6zLQu8tHhJ+1yOKpqvpeuOTCO2l1QWnOAFEDmiAJmPRelbBv
r38tnMtJz17VOG3H5avCi5targYApgTDFPiS6N/CxIpQ0MP/wnjb+WKhTrDkoUjjGBUA00rohFcG
R2WC/V/ID0EXLTi7jCjT3+s4ruLvQ84Ut34lL4wljnj8jG/mmSo0FC6dE8jQVeioNBV6nXA1T8RV
PGz8OsSkInvYS7GQAEnrced+ZxPewoDFrQbgFeWmSQWcgbdQ3RQXwiIdrHptvXo1dD6AcpQySIHp
Whwrj2wKyRji6/yp/QtMDSMrnzlBhkYem2zGqTLpB6mHj1eF8KPAAGU8xuYKbP8d1ZXBbAJiLsy3
qX7dtQJoTV7i1/mjy7JUUx24GSs9tY1dV900yMbM69o9phf0bio1c6L3/3TJyANxmS797A1AK52o
tqzl0H4PIn8hyePvcVYD5Uadeb1Gqv7DmueuubxSTJ/jFkuBUMtn/I4C26LWaFSzUddadR4qI7uf
XTeQo52AYF/XNzdzF3Ew1mcrHAa/A0Yddm7+qkebp68uofrx5+IHH43Lv34a/b/WD/Kgy1EnHVls
Vq8XIStv5aRu2NfF6sd1E1zz53sBsHbwz6Gb56vn+IlKkO4ZwoB+RWRGTwi1BKHdxt9qNFIYQY2G
cQ7QfErpNz3ASauXTnyoYW2dq+0OBpiXc+FtuUbjb8oCXcoGK7IQNa1miY7xkgsnfW3OiVs06TG0
rQcBuggo/TfAzdHzyjnRUQZFpPn+7oVaOLLjhR2jHyIwsS9j5DLRfx0jSjfcI0VsFvhmYmFdjD9A
VtT2IJI3jZW1BQ6PMZPXOBIEAsRN2yqBhqBjjlyjl1NZxw2j/xyybWfC+kuzsbE1XGhmkjPmK5ZH
anIGFh8oDebfcwCWH1oztGb+FjFq9vs5yq43PIoWQOi7joOtPar8Id8Jdm4MpyO6u5InJc7HB8Ks
adpy8TN5eDmTGrEgLR/fGZuYpjV0QEoVPiI5joqRu7250Q/l3iTKTC9uVkmCYhG8EKP0OxL0Drv0
+t8dkz28QImSdMV3XG6rt9d3/PH8lE4nBJNLrjwmpgf6ogBaMhTftOBYr/pJbHSECt4KFmNP2A1W
Bhp4ucpK+Tvavuv1+jMi9AP0wKsO7YRztKRcehZQEl+7cSm2o8roZYBH2j91w58ZcS7g9gxpMnOI
LEVfMhjEfvGAOltINJvhGn4CIiSc91vBJEzL+w48IwOSNYxxT9aj4STvjm+TRqqyAylpiVWj9d6U
8Jf2gsppdQ9ElKjrzuiwf/QBAN6ooh3qlfWOY3AgnYKJYoXZro93ZGQKgH1pWxsZPscPIgYbfkvo
nV22rZfT59MaLZFOXpgtkU8sGIVA53HypB1CM/MkqFC0LR8kIbyKW81V9a47Fy0pIamelEiPSKg3
tlZs1lpHx8fT4Uy8hXqOe0pzpIGIdsXam/4K7qMDeYHe327JqLwv1pabA3X979VNuJwCU262PC7J
MT66lr+hGUDjgM0DlQIb245NptHAsEh8PTGLQeHmeQTQ/WHFCgtTSTnaY4RnGj89EobAOsbQABRi
qGOQofZZVPMzt48BvkHAZsuKweH2ggax3/VtbxwCoiZoni5nR1mc/6EQvaehcJouf/9y1L/Hdhgm
MgiDW0FxFVkCwsN3J5GlOXRZFbvoa62jJyd7Kg0uFQiunO5QZ9zPZZmn51tb46+A0uxkVZnM/F/6
tyMOD4b6shTuNqgLKYJ8jjNY/rcXGQ3F2/+W4cOuyCTEc4uQkMcPUrs0s4lKtmv8YnEXZi+TyHlD
MEZwmsat/z42GpP8hlHtyZtmcVsehhflqGQW93BFrpmDe/wkTPaUQExiNExB+b57sltZv/zBiRv4
N2Oibm69nvLEygGUg7PA6hc1NF0v+tL8gakjgcalqQXMHMl8k3vVzVpTrgEHqKTpAUvQRrx2tvvC
6v0hyArkqgI+K/J5UYMwZ6YmWtC7UA6g9AbcKBZik7gTDaMWoUj7DbCmNWqFIPCc7KduG7QmnHbQ
nH8H+hB5ymyIZ25ndRfELinzLtfDtonVXsUcKqiarbXfINJgePI3Eus7Pu/r/KJon30KB2+UxllD
h3LHEB06sM4/rzEs4h+58SbR00okiriMhyb1EcQouKmyiJzye9MrZh/VEziCCk3u2ed7eANxg/Fl
r5DX9aymFGahciGuPVuhiDwevnbCmmlOtPmTzytSZyoGqEwC7kWb3cSIBP654Vk+CKEdUQX/poSq
JuYb9j1zDCkMFutlqxWlZfAzLFPhCztT8kcDZJqRYcAI454D2+NuGzemItu2KuCr4jOqj0pWQS9y
OaBwHsp1rigchVnaVHFN0CWcD8sTZH5xiCW38WUYGjvpvw0XDvnFxN0PElFFtWTBCih4Mr4kHOtL
9wajkxQU92CyWJSBuh0l/GEwl9y2a+hWBQlvTYtNNS7kORYoQ39MOMf9/0g4jHdAoFeotqO2Twq/
jK4GuyFhQriyajC45/oeac9vD9Ake+1TcuRVNov1ecNAI8LzzMOGjEPBWpmjWRQikSXmaskcrSrs
VhHEtNccLbTiVUz4/SDrWZ0oztTfkE6J1hL+oBJr+hP04yu4/YhhJTohDDUgSLnp4NIYUp+wsq42
UQs2Mb849DNgfNUJh9JHyECsi2fv/X+wg/v2iCHUXTJnV63KjrjQYgW+5zKPPgilYQJh/Y3xMyv+
Ut4JFx66QQpjOD8M6WRWuNDXoJ1tfoxt+I6/79HBAqe5LitPnhGNN9O32+bjxfyFRMxJH84uo1u5
OvgzYHyjQFgG87iaSfRmXslwqJaH8qqkdkMSGprHJZNeFc6Y7ZTvUJhRWYMXvN4uud0USu0j6y1p
LbndJ75nTVQesvVE/595s4WLbVwXJGYYUDZO8SKhL5OoPOnfpgFkpr2BEjhfvIGFUFEiG9s0JAi/
3+sS3+ju5zlC2117N0+qen1yDD3ZPpnE3ZYKvxQQrQi+jA2wgQYGLbUpmr6b0NGv4NKEnMg+RReq
4HObcoCw5ruP+fxb6JQJoDRabpEnQWezVvXUJdEVVYvtTEDUV1DuayYwyug8bPH3vrJlGZUcZuHt
pUoAfkUdapVAOOnv6gDlTpqRrae4TMz2XdJ3IiW9Y4dgAQcwWDlcpphitpPTwmx6OdB1kJitGIIe
bLtrB1WyoBf5rmAGcl7roKOdOGqVT/+bXoeV6mcqlF1k5WpNecjZ84AQwRoncA0Z6cWaV7iChL8O
B0hBQjXHatHqTN+Op5J/UXkNGv4/mJouJTxrNjox/M9WNsRhRSA7dA27STQ38aatK+Eb4S01U2+K
ucEFOAW6OCZQA7bNNJbICEqT/gLR2Id2NsnCby3mbEtsiS8SIOWbdmKL6ZPq7ThN+S+/Dw0FOGYm
G3WblN1yKDymp2WWQZsE3Xx4jCxSptnGPZyMho2cDSYcyowXb9QNPhfvI+ZkaxH/Pc66+XmONaSx
UFictDxxC/DR/ZOsyxPOVNATGoVEp/rZdg58mYLtwuEuCdwEeF0L46dLHcf6Gcc27/ynNYRmCDot
lq0Fr/LjEmF+N2rg1f7DLDRggP3GX5RYRWSiuXzBQnyfp5piH1Tk0HT2pmnkeis8IyAuSqQ+Nx3z
ocOnUEMAMTQVW0hz3J7zGtuPkujX/B86QQXkzHOgcL21iRDIz4GxSEhFe92FQPA7p2//ODCHaUtf
OGejsEeyHwN5s1TwCCQc5VWmsSer/mt84jQzp78Io8gprwVtJGWVJI9xvv5flJvXmE+L/mPygWiV
lXKMcxBScQZceu7wTsPLSB/uP1WGsLMg0mXxSeKsjUipZAXJ5tGTHQtwrUrIDEB8i9pp0Ej155B0
Hj28YqkQMTu6gId/jVt1EC91frDfdFdgXFvLZYyFPfcN4KfSwybVo5VKtSD2ox+gi0UsbTK3kHDH
HsAF8bqVhBfSwIOTuRTrKHzhhZVpXcMytmgDnP5PCsMWPjFd1Zi7lCbll9qC186r8/XG00TwLWx0
pGiym8uzccrPwxCEvzRW6oVSHR2d6lD3MBV1Ri6cBsRqZKe07UgWyqXSrP4J4AF7VvkMUdTziALO
Rl7wt7zKhhH71WRDU7AZNfw2l4fojnDTfBauO3jaZElYtUJVJTCz1RvoTA4h65d5n6xiYBsMMJfI
1CaI6sQJv0FplGQ5wRj2BT3+cAWV7KncW8BcGjK/9Q7vNU0z4jYTJZ5XDZaf190rqAsO+WbCjFRx
aeDmLDg38cxszOeF40ElXwUvhnHCTL3vE2huFFznqNmBLgccC3/jaix7suViqwKySGTnmZSmhku8
yhQY4b7YjJGFg5jwf9TCDZovF96kGAzoLPtKHnvCPAm0T/+4zicmBc+w0s4US41dzrmXgnj33Ny+
gC45A/brUSeHGpsPN0cPCkS5dGoQpk2uwCfY8NAQyUV0wed35Q/vub1ZOODQBmJ8oa9IkAni+4CE
f4UVxBx++JwFSJKKKRXmOET+1XImPHmJxtMfOoXzyDtHEeB5od7EBhWq/TE1a54tL6A6UexElAWT
vOCdmZ3KRlk9ZpIGiJmi3Iyo/tBzUQ4bs2eSd3hb2WngULoPG2uiZbgrbT0VXMTbstf3i5EB+n03
erwCyP7p1iCpwYYmrBW6n1/U6BXmvKLXyfQshHQCMIvdaRIypnDV4TiFBrJ6UajtYVJ8+06ReTLm
4qJhbFycUSyMD/Jy0ljei0ZrsAiObTrhCVa+xVZgsGp8aTbXGHkGfuKJ70yZu+8OHsGSMQmo3g9M
sNhntmXUg7ePQozjkROywhC4Rzwqhhpc/Umw6IEo+WL2Dd5qGqWylzzM1MxomxuELxO63QLnycPm
xd4nkZATCuj5+fPXxgdtJm1vQl4AQq8081k0r4e5wmoXIC/7J8Iu1z32h7ZYILzzeWJXtUQHdr+4
6CfPCe49GU+1UBLxTJoUOvn4kI62cYBeF66Dz+ZswJXWhF7GzJyakX2as4DtXJLBdDqCqMHpB4HM
YPe01Q/P+RcnrLlUWYHCCE+k8KkRn/0gkqEarfTynApu81ny5CilPmdxdq4O+wu6Yq7CSWRH+lPM
hs09jn27dj/djtRoB/CUOAudgulP5FyImTpC/X/WDK2NWTlEDoS+syohMCWIotddkswVJ1zWHghg
/Jg3ePvIvmK5XXEAF8mWv3yVd5+BJKYgvrWzD1vsA+q4ARhsylSS579HVLweCdvV2vMnHKVnBMX6
eto9Xffjfx2SlRxRRYIMWtRMasWeSMiiECxUjav2Tu1Hcrbk5VayRqY0vHt4r9zTq+Keq0wU8eb8
1T4C50XTqDZAlSqOqIOzKSeAYFovf/un/+JLBcIchsD1ZPR60yBCgSnxpMVUO6PTZ0M+S97yA2oR
yfkiY7QWCdLg37/PTvCn9Ze3cTLShAL4kor3gOO/e5AwpN6ATyF3GNrVFUaS8MtHHC1JDmcfM6vn
9wvdpuHST8CHc6n38WaGZVAjnXnYo94oR7pmMRSz5SCH43/ZQPTdor/1Ahps1SGu/2lT4anecSs1
FtHxx7ZLwpN+ywh8YVs36iqpeD8Yw0JsgiWrscSCLwPy7SUZx1tpM8pLbYydbTczoW5ttk+ndKtG
PKPVsC9jc233b1y177ilF+VOWJGEq4zPGkDZug0iSUCCwo3BljLiN6JHlVu7ev9Nclj21QD/nbx0
eoucQqwfZKoKOsRo1CkGyVJ/4/K8jDRJ9m32fJ4X1LPM6zgCcyRNasAgY5nRp5WLtE1RaSM9iP+2
k5Vl+JQk46+kf5955b5dW0sH+ZYDM64kypRs2CId2VHFbDDMUPJeOsC4ZdmipMl25assU8f1fGSS
R88MzzsT0F+uuS0lYdVyKH+WT0bPKddhGpVzb/oViyjEd4HYFqClAIw37uVwXXfueQUFptOtquGJ
X6R7IeIYWlC5phr4UoIV1DsWg+0oZXQT+sc7YzYbk22/VU6fHyrPoyffcKuJINl9h4RXYTgyXU84
491xrvaecUv/CIF2Ja648/uQMkcLFKGjtLyic9n1/wOvgo7tTsxFOJs6CB2V63tDRVNGLpA2IGOl
3riaCCjMW9l+Bf15fG5lhNVn2LFsvgZ7eStkJc8lcDK96ayZpBryYyxksQlCfvblddjMSi+g7/fY
eApqelKJtsP9BT1RoPcVfkExWJm03J4Ikld7D7tbzCDk84b+J+S/T3yweHLbsrpNwhpNQgp0CMrq
AMuZ4Ciup2ZHHmLbZpgVn207yU5NR3nfTJXr6IVtExy63JGcsmaSGbSM+FuVXpdRMspLk6ooghdR
F77v9/uEJ0tKGxNNju8SJ1Z2esXCHupQYqWavmVE4sBnLtcvTBONBtsBaAdMnAWKxIz5xjNZk0xg
dtw9cVapEZB/rpFKg9mRLL6/Dvtmr+dIlITxvF55XNY9T6OSBR/OYz7oe7UGjIrsoyt5T8FRvNJH
jXdP8ptxtOvzwCuMJdcHIzSsA9UuXTxn0z2OPxMyBam5eWytuUSFW4n+XaKZ8/AGDnouhhISnNRM
o6vtxJlCCNbLhvHuXuUiI/uHs+hJfDG3QnT8LxV3B+FW9gqO9nNvo19QKkXXNSe2j4HXSDkzXz4c
gLL8WOBCjwqsyCoCdL8F0zOfeDgc208p5SrcTL5g3RwgLSxi8h5DWoPTMi8347zWAxg+q8O+jtzh
0MAzrXxA6gIgsqEZ2/r608LMoyRMQBJS0XfHpP4bg8KEe5E0qzr6HHrWPXG3CsJx42zD6mIlDvbd
/9WTM9GcRK7ygbG0Sjo0fvInVXJdtRLwSK6k0gWPTzKUI4Agr3Mzr0hPSXfod67g59n1PszRwhyo
bH8uEJ9RQlvm/IH2zZ9rcUMDgO17aEkwReOgIYYv1GJgCx7LBARYEofKrbLScOmBTSS5CyiEaMxf
iv96L/s0Vu+1wPjB9jCCofhnOy1i/1QP3AP+I7i/Ok+tW7ADHXHguQG//RlK0USEZFxrKPrMmJmW
x4KrnotZQkVZS6/nKDp28ZG54zCXPJqu+niLax81viA2+JCZ3J9xa+lh5zKTCIrIj7SQ21BvSkrD
PElvR4FTKKdqfMFshgSXZCS7eqcoJXQcS4yhaoFKhyDPHwLKy05NMgHqVItWkGah0MO3cGDOm3oF
bNFER+KjRXaXyUS2DAM3+syyuolAKlXCCRA05P1yniz3ynGb3NpuqYMCCNJI6lBxjpcVPZkguBT9
pEm+AgBfqJvXO0UgSX0/oaTLNnXMCbD/VCPyuf3GbmmPWCAwbSvSPOvHBH4T2Ud+Qq0z4cyzQm6Z
ZeXOB766DnsK1z4a1/2+aTRgxGgzIU5k8n0GE5eBWifEfI4xesohRTkEyxPXv/nbiIr3vPIhpXbx
VsS0U8TEIZM+/nSCrfSM/fgzTpVtaPb7J4zLDjfrqfMn7qofbY5Z/uQO2Rf+pztLBSeKoKDxPkhV
odUbHhjJAHyJVUc4+UwqCf7Wg1LIMogZxr5w2FXeFZWmA+2Zo4lhMyoRgNF7rmwrcma0q9lyLt8s
4QgAqAQBTiGOuVCjzWO27DAMvRtmYSlG7yLskoPxFiyt07lUs8MINvwcZ5alk6Kz3Kju93Xy+32d
dogxwq9N48svws8DgRAbOm72aaJ/KPr1d2gsV7zxcYbYonh9BZEM31uZ1vbMotweNotT/PPvHGYM
oT4e9soh5PoDpNZiQgVEgkKXGrLMN4YKGE2VQrh+TRFnw9x5k8BCc6dYp+O8xVX9DqyEH4r+auJ4
vZtsqogbHEzxQeFXhAZkP0dm/vC1t84d8cFGXHyjyrN96n+8hTWLHkiHrjv4ukRd92EeADh4Xu7l
fQGR53xz9NzvORj5GroXtWApia6+HDVGd3L1JqpNxfo8xKfIKMCermsZZ7qJX4KL3LlnuP9RWoNs
g3XxtuK//WsiMeXueRl78OBemdR/e+nkzAdHSpoR/BeTQoYHE2R0XU2xBHK65yNmiNuGbVMYKlhv
CDl4OKmHIVMk89l9pbbnJsMerlrvknCcIkI7QU1DD7xdCRppO19a9xTk1lNYLEdeNeIv8KrMMQgM
UMVmWUT6y13l0hH8YZYcAw60KRWFpUNHADZQXsS/RdppH/oew6CptXs4PuC+lNr+1e5m/U0O6oct
WXMlPO/nFJXZ53LqtqOzu4PGYYagDAFYS7mh1GDQD/zpUzUtD1PEt48QsZ8f+6eIwjN/oA2frBi+
6/AdRpfVdSv47L0YXbVvAMlzqWW/5Y/nuF7M9FsOJjpUIJqOFnjrjTIw9cNaw/mOOJ+qGKtiegB/
CNBAO3m1F18BrAAMEA573mMHX79CbEveD9xdJMfZoqDwXMwhWdzsWtyIgUJoit+EDE5h9119/dCj
2VmS4BekG5bmwKhK7tBheDDm9sUTTmiHTO1o0w++FvXbnTM0oT/YKflZUrQmZvHDOLpCdtc04WWy
owCIWMzQcvnlN2c+ou+PgvQjEfJ4sLTPvIpEkyHIWwAC0dQDSCeLeysJAhY8oIvUaz/6jkUlZvby
iSSF4OFKwCtDkuw7W5zMvcX/2IqTqCUOLtosVZfDrDyOTLRngE1u3uwyPkQlohXSf9OuLKLegiMM
mo2H+UYjP50nJ3Do8gIZgdpfi+o6ZeohaTOHPM6J4IjFTsU0jiB87wtoQMcdbAc7Y2oeFg1OIfL2
j7Pd2aPEvZXHtR0lZrAZBOARtBjxlTEo5/wwIMp9rT9eUIG2ORwP8GA8SA6tSmq1kXPA066o9Uwk
rOE7yp9DLlnLmR15ZHOld6e6Z+i/9p78WxxcMlW9mrEipfzove1ZFvlEAvBEqd1BsoPowoW0hLjc
XAmmMMYpZ+G10OKteNbWJd8AjXuQln2iyG1xGei6WuFLFo/rOTjmJi0bOI2PtC7BNpa8A5mIikni
3kx8oNuWeklVz08H5gHYudgbYdzGoDhin0W3y/qlj21goJyB8CN/2jG6vo2PNqoWh41c5X/cQmmr
asd52jUOZqnxgA+MHoW6JWySSxbng2nQzBb18JiNFkp89LQjCeE3QL0OSn8Kjo8kLq2W4q4zjEBt
2Xo3QJy3cMXH0iVIGbBGA04g6QPN251J19v71lYQb5VB22560s4WxPl3oT9LNl9j7S5+DY8bOEjE
ixFGL7JD8HMMB/n9pOG1ykPGadcNg4QgGFQJ7nPISmPiu2UXyiZuO6elJGHiLWsMCMYihIFdxZUI
c4XHQiyYHt1vFtlZ5L3Iuh7coqFTjqdTZEDeANsY1srWnIFiSjSQBgW3ZbUqYyXEdGzGLaypNiSP
77zDjHCwfRhNtFW8yxJ4kXJ2UE1/t6h+qpMzvpA9fN/0ToOODbK52je0nNpl13qOpW5F5kexRmyF
T+jPE7kU+7HPs4feMoPRiAIcXWqtnW3PaY6Bj3LdNMMKQlm2bh22Fk7GcX+yKx1tw2hbd1d140+t
tOpucECAnW5HfUBINlMfNW4kxU1QRMEHvb+U79dWEV5jRiIvufztdC0yl13BoLFbHIpUu8TXly7I
Nvgiv9gzVcqtL5RBvaUFpF3W9n2A7TI3wWHPoLImTfgYj808vLpbTfNwV14dQOzC763cnedtfMaU
4BOAlOnpYvT1r+YKJwdNa7/pRYbLvAcqbFzUF1UUdOB+DA6+9yjr5xjnYZECdMkAsvhcybiI8KZ4
hltM59QuYreHv6yeHPC3RT+0qnchuhmMXAesg4cj5c3DsE5UFx6+59fw7GoogMaYjUQ1Sns0KbsA
89u2921r6MwL9Tj4tFC7/8SwURISo/wfHYskI54EG6iA+VN3hPmHni00FOnhnEOnpcNrrn+W36us
eOZKc3mkiK28aOg54jjGqc8K7Umco15PKwDDm/wXpkCBtE+pGucU2U+kKsCKFsiE4OY61RNY/01j
hKaGl3mewhFoyqNCWMfXAh2H2WGWwkYkpMrLtStGrdaDMmUMRuWBWCmG+KWVs7o6JI4pLLZM8ziE
mNwsI5wBVoa8Hl/NvP03rcKfvTjJ0pv4o61miPetAxi3k4uJGJeTAqskdeo3S92t0iynvPRAw5fw
vEDzy3BzwHxEMkqAiJrymup7dsC942uWTJpl7kvBCF49pI1yb+Qgzp4A1FKLhW5zrI24nnyteBdu
Dxh1WlYhf2mBZmcpns7F/ST5uJOAjDHw/y3DwnrnaTRQTP1UFl7f4gTRPAJWFip9pKmcS37ZCx73
Q8rOHZ3JH6Np0YXUiEs2qYvam6i0zrX3K1xuOkG8Ew6NK8vuhjvlMNF1id0XnrppxgRkr1ps1nV/
VtPrmdadJUWty0HkjUyUnKQ7dey9vO2tCyp971EgwakIncpgmKSJ1zytm25dCP3qdBraJpG5AQT6
XczYFqR2oNmpSUeRAeh0NKF+MHjujxsh2k9B09bxO1K4d59DKLLrmq07BeFMqkCXUYTp8Tzam3y5
9NVvivjuPbPrhZ0H3ZwQ+dRuQilp5B1MOiW3sd4tZcbm7UoFQ+tFni2Z5ZMvRjEYxYQfWAfbTBFR
AVFSZ0QZcIoEQUc3WoFr8vACDD8Mk/q6AU/c5wUgWQFs4TaFzk8ToPEcJb2+0HPt1WR7CTDbvNU0
/uuuvY1NRlNw+DdFtsiuJJXuL54dmmS+7L1DuVJIzXSGfPSu6vaKft15e9Qm8a60RdINdYnt1NgK
WjWAxApVfAuTco6PHu/wO+wV/kkm0Dcmet8xHeMA+GkqUEeMH/suoRn0pMb7sE2LOQt7B9Lde6Qr
UodUnKm52re8IGQZLsxXXOtqZmCgqwLYd+T+YExmVwisgWf0KfbR6hDOvHTerARcBLIv1FdUpgBu
cfXNQNnLN1MV4Y1+NBE0SM3IBZckytUPlxaR4eiH74lPbzRKGmTx5zG8hodajd32tQo2mOFF+NZJ
ARVXEGVvKu8JeyvKZjrjX1bHkSd1XLueuSrKNvpDsRBa6EjCXmQIsJRB/JwzlJNnyv49mAr2QXFj
qtKXmO0hhivW0ySYZOUikaRX8BQ0TMHhMpZJGHdHsWNYryPCH/lTglgzNiAOi/deSMCejkqJrY1s
fcfg483XopIg20UfFv0Q+P5oiLfYIW4xntOA+UF3LsfIxfZzKA/AuOgB28e3FjOlUpC3zoWp470V
v2vnuniLn1Y739PBGgGlXkVS75vQbnaJZ4A76OS5zc96UuRFL9AZ1F8fzFGyYGUSvyj4msY72PJh
NYRIXut3tLDqxRkdHSv1rKCpXX6Y9pXv29qfV4IaGM6mCvVfmYoYQKN2OwgSYEW2nB5rOIFBur9s
lUAO1RO0RZneah0PPcihhquEWgY9MyZ4kpmvm8lbfveDOyn37ZNDiEn9mGKBIhNKYVtA7LwueifI
Vhv355Q4muveDT1vjAqrHNciIsSVMH41ASehrBvHDRItv9aLNp6DQ4MHVctz4e5+fdBIB/VGlDkb
xqO4juzlwqGE4uy5aP6i/pSrZTYXGDkY4U5EwD2C0ABvJiDBMDuFy2erwDJ+M3nBv6y4R8GeXm1o
6DB06VIcs6yqfcJ3qciw63z+88UcDOiHJiE6JWPejMqpEwJizEqIJGefsH9ZcxvbzFUCIBcYRtnx
jPbomzeLqT//FRWkm89cUHtsW8LCroMsaTKLNO0z9wxWtWsU6m60fz+IyS5CxTK5cagA0GtlEvhx
NlLbAfy/EomPJ9nocUSmxOEO+BsRIdrkLIBwXZ/XORU9PBM02cHQeA6MJRwK/GNeZSEFH/RhJ7+i
woDWm936hBV/cObCbQV1LdPaqhKoAdb7OI4aISRQZ8Kcjh5wu6AORjBkwI3Gbebu5idY/NGZ87p2
I6fy02Sm9ixyWY99PeFS9nGXT37FyhQ3wH15ekc0z5V59EfGZw4PJKVAQHEWfrLeYhMOyQu1c/Dm
TaZoGggfFYBt8s46Jp6gr3ANzC02k1e3AzKpa2wKV7ycm6iyUQ4THN+c0MHup8j0NtEf6xfGD2uW
+amZFSG7ZPms50PxupEkdw0l5YblexvoSeiGBFZkj9qt2ZdUWZp1wyWhos9JnqEtIaQORQKS+tLh
R4gymeeegerajF8KY2fF9jkLWOuPeeCKPSBA5TFU3Km5NgbodAMIAjDPqdaAQwZPMz/ttvSFEuIl
cjs40t/Di8n8k5Dpe6hQFdQR65sheQx6qDtqpV+4Q4LdpKVrt1rHRnjMaynW78ytjn9JCDur6Wm9
otIsbFX7wmEOJjwtg9B6jDSRNyYFELTIzd57a3UCk1l2ArKstFlW4a+9IKRuIMZExCyyupYt/GNn
DGfJUldGLo2bExO0Uhlt0h51gpyrIJUgjxgyWGrOCi2qAWYApIMshIWrHy0rKkJZySEk/XfIY3do
NjzGwALAgzMyawjE5/DajGUZOdNCqVbG5wwj7PaxAPPi3keyqY5No4Phec9godfcTLWZYRNNAW/I
fjQRACdRi2v4Q7t7coxvBQOdBzv/IBJkZ9ZAgxZWi0I5oHK13LYHVpO3g/3AhDwBKHgpjzZvAlBT
59c1gkDF+iKMgX/G+WB3J2hXiwVzM7/BbZi3YTWg8/pNvL2E0sBCqwO7i4WFP8ALKfq+LRFKgVio
dcUZjREGaNxpWREHJDbej+1zHAt38S4JwHy4IDbpKKfL8zfeLl1fUJjyWbxo4zESrGgyH4mos/lP
0p63sSoVNdVj3vBfBcbMPzpcFJnITwt2lLFCOogzHUY0y2JVeY3Gtuilu7zEdOQQdijEaBoXD+ub
4d1UA8hLtuxkls6CZVdvrtqHt8ZRkcx4nDEN1TWyQuq/xqbbe9UOJUnXjautZ6X20YBilgVuOxh6
zC16edwYEOSZwrtNsXjRcE5xe9mJ1gB4SdanOyRCw+wJ8kCo7nztm2yxfzabwbITHdWu2jjPBeeQ
PAgdwAC/EsccHZ+ApHkMB4P0iIp2xjDuJ4avqaQWxoGhYsDG6x/y0a9Xgumazva5ZfjO8LJZ1Naw
Qe5KHlC7AshFq9KhJ4Mapowwetzb2P1ch6Oy3+XbxORaDRNi4B0xprq/BRIByG+yGLdp1jHmpRoB
yWsK1MP2egCPdxbZ39ngVLuU8U9vueui6lAt24IeJ5ND4K/IYqW+VNsvr9tfSp0Cc1zq5AY6sStL
EllgItTCLgx3XfNCGe0sEo8uDI1RkdFLDAP5qSkmzM6D5E8X/ULeK9UdPXdOaRIoPe1j26YrcT6G
bLwoShGN4Q+FQaf+TEJKWWtDovH0JKhSxh9RitRcMVyIQBBpDZ9tklPT67zh3i+KQMncLfH6llZH
ZGCZnahMEye9CG/A+9YcsoiQkT45qx/X3Mlv3o/qmuvmmoDdL21JpvhePXUBMFZ//tmIAq+e7er+
eHu8Ruf1pNIbOa+WSAG6GVHQbtS7Mq4EvZ+k45hYusMRoeMf7yapK6RD/UxJKwVouT1B4Su+xtwQ
mKmRsImRhuebBuwCD7IfDzr1IR/o9xe73W3/hod2BcmsZkMuMR/b5YmQoxJ2iR6ty5VgYiQ/Y6H9
z00qhcUo0bN36pX/Or1naN7WchGYZaW4lyT+TQV/Ro5CRutQcvvJUUXFKfnvgV73mhA72uUpC0DQ
NbGm5mSoJFx1V1nXzk9VeL4BaXJtqRt8s0ie+D/mIhyJ7a4og1oA3BqBAVwO6v1NDr+P0tUzhz1c
ZoeuyfQ/XET6x+ON/HQ7LgG/Rb4xVfOTZ+Y2tHlX4v04uCMgHella97BBs/hTH1lrg+xQoTucV02
GUiZpDmbjI1cY17Of/YVSgemH6CoPUk4IlGpOtlvnbM2ndoQD2YIeHu9uXkP4eaT+FQRGv7aoTlN
XiMWnnkqJjVbFOMCW/Y/4Hfrm4FlIYkzHUeHzqqnuN2OabK6nRoqj4p2SRwOr99q4hUZ25Orv9cR
ZYdaek8IjOiFuUmPPV04ecVNQFv0To0o+YkCWljX3vUS5//imD58tTZTR5CZ5qX9vPO4pQYfegY3
JLqBgITNJsr4D2ANLOH2BSJMLeNSUheuXBJIV1oqv4avnJNg9gPFvKNz704JrsPrFl0HV/k3FasO
CvuH+U0Am1ICP9xWUlxpNrNydegJDIrtVZF3CJYRmr2jIV8k4hTAfUez8C2FTJLO8hpsXB6Gp2hH
TC2hCti8q+W+JFCsQ+BEBRSMo5qU/gmQVIQNtN57NjLT1BKh/JUwlwmT4V+H3onN1aJLwFSFecSH
MQEKA5hON79y1U1yajDLqys2i9vZfEmja4e3VAvveFmPVjFWsZm743XrOOztlcUCj+2ERMRfQSk1
rZ9l3GOAKdQZ+i6sGlBFN2a23PG27b3lgV7A9R8jAuOIALj6hYEBUmA3n9vUl+TZUCgwEa4xpC2n
NSqvl+7V1gLdzwQiBqAPk8/wobKRJIJJ2sVoqmm+PCtkQjMXcbpNhCpxV2SwLZk7BhaQdJ7IDyeR
LP4oK1ziHZ33jeTI3lvbsinfNEYz1YDPklYb3tRUd3uwvBHLowKN6Zb+UEkyo8HFpTh75rvPwjQ5
1UAwgLwxcIvBreWoeyo2ye3Y/SNupfotf7SJArv2SzxL8O6P/UzQQN7DZhewPdVwUC1a6MjvxL7X
HURVmK81ix0UViHNQuwSC1vEdjXjUi4X9barBGRMeJTcP2+fmc0M3+ucIZ/QqwstUB2tD0/DA9sE
iKfndQMw6R4R1QnK0ivbtMcM2X4rLj/INQuFy8XS49elI/lPRLO9Ku1ik8Yvf/VQD1jWDS7tuq02
VKQuwHotRnY80AT/vE+nZ0W4kF3/O5puLJEJBbvjrGuN13+K1ZFUI9LpdaJKevuhQ5rrHZ/pWoMh
sLpkxPBon2jVCc2m0sAiP544J42SA8r08XGBiDENWY0XAXfIwbW/NvhZo3WaiKl5lvBtX98pnqpq
pW4/pF7oSlALZsK2IUEnM5kdn8B7HiiXTmRyWLQwaRR1Gc06ANGIw3Lj5dT598FJECgS1Fz/bwaw
mN/mzaf/dN8HXc8qksZEALtoRjE4nIX2ITSQWUKiz0kSuFsclruMr83riLiqeli6qUogspLhOA1d
AmJDnDw6+yUc8VuTfcVIwp6kcFz9bQ5U4zymqSsWZARPIg5hdKB6GG0XulW8V2IAaSCOX/DbCabR
oCt89xj8o3tl/IljQcyFzRdmHBTCVDNulG430tFO8r9CIsqT5FDIXcBFvtXk27vbX8Nqk5oi84w/
jLabjTcNxIB0kNAdz1d2Yf/LMMg/MM65jqjdPNhoxNV404b2uj4CPD0gMaw+wQqP7FzlQ+Wsgddq
qLLhY3Tfyg9/1JA97tkPd/PT9GpTC5RYmDMKrDFkrxeR/JihTUxSW5n9EvYe5/6CTSAww26aGMk+
hjTzjxj0U/NjU93PPKowc0kXspr8aQdpewK1T2kzjVPCyxqrw6dGsguBNVQQeWggBosdW2O6Nwq8
T8+eGCgnyedWTRtVuNOBsTWmrb3XUYU3Zo4urODR2pGqco5rwEart6M9JbqgQ2114JOjelpwsaW9
MnRrORy8EjabqQMzU3bS4JShZqQYqQ+x8EsHiJUgRCijYvWQwYFjYDtBpBsQPyiTlzReFvsG9kMY
rwoUhNSFj9uYP9cUViJObwLiptT48bEvKp6mCHDYuaQVNlghNgrx/rNb9qViCvoTDsBsIrs9lMrn
vtDY7BIO4CuZaqDcXbFaCTauziw93Y8P+bkPrtd+MKWOIqs28OHPUUcmRo4n4Af8AB8d1xOZF9IP
DSTpNFNWpqtqrVs72nIheYqqAo1RxiQOEQk66ZCFQqsw9RtZUZJv5X6MkPa4JTZtWa7F63oSorLc
P1QpSP0Becp0ghUohr+fWzZcmonjpaqa1lI2g1ujdP5ImF/ZRS6wB17bhoDPXZChAMCkD2xM6dKL
2gIE3lBuXOOK01wRyGzxpmomxk5sAl2p8hOOgs5n3FQuYq5WnGoBThzyt178tjPNxfr/jEdPrd0L
WkSzybdpqYyYhqC//G0GaSH0l4V+kY/IH2rnrgkyug5jU1xeJgLvovIlojEahBLzbml834aWEWTW
84lvIQxJiuJ6KgsxdpxyW9bNT19RdfoNHepcd9k42PnnnYVxg+HegNNqfNEHRM7QG8BO4074JBQV
OModI+fNEGWsWSpPZGjrGR7JDPBS6pEiiTB+nTtMzurZOQ4z6NOwRLTPqQ8jtMBfdhBYN57xeSIj
71H1CJEvc91l/KDLase18aVRiXV1yFlQn68rRbyYWOhsuCfbjnJQifk9+QHDwsAA0VVW5D5g55Ja
FRKN5KcQBVLj27Nfe4KgQbDql9+1sUT5RWC21CJBVxS7Dj4UgKifdH+its9aE83AqQBtfNnQucSe
BofZ7/b9Zm0dT5gzH4sto1HdAoWav+7UFnJyQSzfAvHqF75OmKfvNslJltxFlDMt63g5+v9Q5tVT
2AUaZqoOav3xVgQjqhWjBbizgexh6UuyXJyn/bWEH+FGvvAs3CfJvbkNlb86z2meMA4FJcPQN9rf
/Y+NebCCqimd7Lft7K8st9SRKjxSz4J9RrgNiJ4DIhotktt4bBb458WgIAZ75oU7lFrgtkCGtXPs
GBt55iuKtfUTifP9sgUPSeXMOYl0exz6e+1tLt8FeddM6erbPB60ZvtgV2OVI0xI2So1bAka3dPh
2nLn78rPf0iK+P0wPg2Uf1uWLVdvN0V0pi3eyaJpyDK4rln5bN49TvN4tFT+Lk8dTXYesAqadBY2
ur3XL1Ocec3Nr9w1rArU5Ugu9LCGlzbeemsr9aAxXoV4aSfhTdsoiFuoj65FFehzql0SDclCTVC/
yiQF1egau041dlaKGPriaNDuIhFr/JHjGBHcr06sIGdJ2UZFPH76C9Wi6+nJK3qjK4mFsjB+tiqq
Ph1lvCmHq5X3KtuKTUJZk4BiOc6BegcqcmrYGbM5/HgFvXZNlPUyJX/ReB13M3sstlhkHqXyPK+j
UcQpuApCah9WMMwiQUtcmAuDBTERrC54V29NZ2hXWa+3wa+BwhQc+nzq6PnHaslhzpiNsavUMbni
rL6V2bwGTBx+JgmjQ0IjkmjMB14Gm85L91oe2t7w47UxwGhJILGBWXqJNVzaytYPSgxdqOpytpDs
ato7m8slxZgb+WEhRdTDSp2KHndWxOhxeyhaVm0PL/R7GFRy5MCmbRoL6rwCLclrieSyx0pCSVD7
UNrFwHHuVuidcDK4lnjK9ziXjN2JhE8xPV7H2yw+eLZUw10whhmmuffmCjpROCzjjc1LJwNAYj1T
Bo5Aj3qeBJcnu46ZBbiWfv8E5AGkQvQdqWh2boguol8dYK5y8c7iLGjYvSeSWtwlkb7ctpapnSRO
A49HI0Cqq5UNkzrRQF+3XpLQkiZeOhpd5p5686jb4JpwwQ51LvjEpjaQj2vjD67VEwAMjmsOoHHX
6AiLoHfPVznHILKfzLpdgBhECzHcya97e98fJEPPu1HEP87JharEH/2V2kaFJnOxohFaPxhaebi/
Ez/MOGnLt00xEKxHOqAFlGPfsFktrLyx0qp31Q+PN1EMHPHWCy/Y51cVa3MdFNam9zVdquImaN4f
ofRTusIsTjUmm+BZeyvHmxUr5A+IyWG2dWylhIyqdTAiSGEPtSgyzZ6CN7XhxO+zeYxezpO9WpTk
Ln+tmf+L76/QX/vCR1nSSlRUQtx3SVofXoXJkVo/3HBgULvZGR4mJD3kX16N/u90p4g9G0AaKhmQ
YmW2KRKyB7/DEhHfz8sYm0qgXtshYUvBfWO8VZQQh9/25AGxhndE5ADPYrxhQl03eW5bi31POfM3
g0hQLxDDOhnb0LFH4wGK2+sjR592Yk4fjp/0x+1auVCTUywuwoDxL253UNosMrFQlsi2INXaKJJM
e8+r8ggkHj6nNOoguOLPY2rCTlNjBcbUta1ufxU8F/cu3zbvXE0otGSuRrxTATqatdU4IuklQyWo
G5UAb3s+fdtO0Am9O6NrPtLcASE4tYC04V8aaac1d9/cwXl7QpTaz2VjW+gGXmnCl2EV7aZRWUjb
NHGsE9sMFtyfNLTOmSrOrCjy1ci6RYwQJFsK4iHrqLcuseIAO2K0SIAQEXeqPf1f5R1awZba78Jx
3w8y/udfObfYN5BcIm0e+6c5st69yrA5Aglzr9/ldAZJufLrP9BrHTxfcUGN6Ydjz3Z8d+CNg2pp
8ZLXXYbnuI1XyRcJHlrbqaqEsYTrz4P+cceGxWL2YC5jya3qJwXmeaKVFBfN9fCErdMRATq3rY78
X9umnN7zkFPVhsguDCzxXJKNGeNKHLBpVEXg6nuDz4iswTXq63pOtmp7GZ10aSbKd/14eaTAYsgY
JkX+gjUJKNpBwVBuNPEf9R2nvZg+3VJ9p3SDDW4V5amWlf4ulG7X5OzI4P3UJlKbBIH4TVIYjsqy
2nr2pAnD8EziPUEqzAm7ejIDPj88fp7X1HfnZsKmIwTtKj5Ut/FH/Y9ud0lpe8dC4m0ZveUnW1on
l4Sm2YzadvBYudVb7mpQ6LcMvn+cMtWLyG+zOuqw/QWvcqRGmd0HlLQBxWoH/bm+lKrfipS/G7a0
Ew1uLfD/5RnN0yyCHQKZSxY43Cf9X2KLr+LX5ogDjE9quoFDJYZl13XGY6mvNPVwGPRBvF/Kv4Fx
i4rp0cqLKfDjCvENXaOTMb35KgLwzx0lTpt9CbhsxDcIQ8WY8uzTkZMYkENRgNyrGBKFIeP53lB/
+DTASUkS2o0cMC5Xf33MF7ehL2E0gYCuO5fJyJme+tJ2xY2NyQr2NT7gZ6pEjc5NBl5J1SqruRAf
PbNui6uG3EaaAN6toDVYmVNX7MRZNZfsGQ0Bca29SVuL6ZhS9efd4crxjMMKL7YxUwJzYVogg6KY
xRQMFz6hhgsG50DGsK7ltAVhq5P6ldyVIU/WIEEje9w286bg6wWEgfqdnub04Wil7pSTDwmgYOWd
WH51X49D3E1sp3dCYfsA3V55PpGcOYOg5muFdLLsp2CVsXIPZvmhBBvBF7bbizX07zk99XlB3KNK
05p3FkhBWzCiLjL5+VHdUN5Pb4iSple2anvKjEMRo/YnivWwJmc0XdqRPpqMCA6l0WIewXui11s8
jvEer1G1KTEGcZyNxSc46OQeUFMwbkMmvTqvnBQnJ+zcL0OEyh3/MLozAtg32uHnOWH+jxFbarrf
pJry5ME0hvhEZMrUKM4zeSRPppdj/wf8xVXr75u/ZTite/NUaDdTR4Ym8o4asZZw8IkgMQa3mCNW
UGOQ22MLZaWvyKOJ85fOYRQ+VUCIzBmN6i0r19mFAqVeUPWn3bpM7gnPXkTc2daZRTuOAKOPQM/J
6tBo4PPhYnCzOYjzaotaVAr48lWSp7JhR08uNHgGiMOnCf6RfRlgF1488xTh4AitZwZqPb9P7eTN
JMsNxuUWjle4i7ms96pF3b1RAeHhdasHP5Fg0TLFxfvGrfkLFOazA/ksgCDc8rdQ3dV7oZ5Rc46l
2P8zeiPovixajNVqQucR11ItKrXHapparCeAEAqJCVza77I39VjZWeDIViybvk4edUvhMPQVoPWl
S92HhDaoQAFf7szx6UQwda7Ba8Wf2hUKN1qXMNApFUBOGkFAyXuvojXJpHxi2wos/sxSCBYqZK4H
iOr/nnlm2Vogge3r1G9HR7UfkkTTlRRxlrCaqks/676bbq4BY696g5n8rmZ1MCDPTa8L5irgOQ3H
vBNf0w8INSJXEJ1ZNYrz0gOTGkkbQOdzH9FtldYRa/JYDZIf0ARLgMwapejH6I6CytluRvaAcclE
SrvjOQJun1c04as0tRBSl48hFou5g6QyP6sSTr+YbEFeWhpm+RCxhyAb07s4MDass0hdgLPCjVv6
bX+nSc30Aic78aePOdYAS7F8TJM1MiOE7gRSrXy0YZ3E2MnjUsOi5SbBNwaLtmhyyxZyGqcB/nTO
N66aMk0qkzFc5TJFHKww4eUpuF3f8d68DEaTnDEHXWvf3UNRU2XCRQ8Eh5bcoT69T1yLEUM/uqrm
adqnenbhHkxsZU+gghHpoYOBcFJgFxmDln/ThUXQWIErL/iSxLTCRcAsZYA3v1GGVfO4yOJy+5DC
eyAdh6m0xcD3+jf/erATDO1DxX97N5pe/MpkMZ4YTwl/DsOiMNiWcb4xLw9FybmLXBUn/fiUYluE
E8t48JJMIHKxGWUIKisdAaxNrUV5dYUS4SrVMxzuasV+RbZWNTg92Nn4GfjRgbj4Oyj0y/oKtZfe
6aQtydyg6kpm2GDSYElBfe26J79usDBvd40QmlM8ifa/jn4zAhr+u25p4eRx/O35pXlPkbzS1yLO
Y4m3CYLYMm9PsW/Ag7x3pfdQqr3F0SPT3Fq79m8i1CnR1kYYoNgk1ngy73LYEQOBFHpxqh3QURae
KQTt9tJ72bZZolXQd2P4H10+tkU96Pr0Fr7TIxYtpbMu+hWkLhhu/bjFr5kGSKpQYAkr5FcTekBI
YehJq2NSd8L5ksDXmOytrPhzFA30MCmArSXE0jDAyA11744lOHFHaa2QjnZMX4Xe2ugxNH0Q8H3V
W2ES4qlE29WARXMsqLLvxIfuGDUmLg8YJ/2HmRngfcTcYkuLu6e18woxu0qXzU///wUVCLIlkoFn
29XVHkZPHSvdYGlPSbiSx2I5WbR/lTeirH/ZvAJhOQ2Jbtc7foNkBFhPpOKFktCuCG9jvfGDVtxY
uV0rqWLOXOW64+8ZdcNRXwxgI5rnxBoj8UCviwM2nDdFEsS5Ta412xkhod7e9xPBK4Sh9ogYVPKZ
+M0sg4Jxnx03a5Y+ld8CI//o5P2gr5NnYdIdcvtoZSB4etBuu95gUQA0jlGCQNSIqUATUyNeM+Ld
1bxtKEv3h/mG7AvDS503KVv6FbhRCkaU/6CtJLOgJMQ98GCPA7xoICDAhsBZbfJYQkEgU0NkYhHM
3O0gAMCaKGj6GvGkY/jB+cMGHk93A4mcCFmZcOHw+5Ey5Wv3UuEOXG35rftMKGyKbdG2nWbJTQHQ
35Gdlm/RT0Y3Jdz5zFGhisOZwYLNj8HpkAbs7F2twXZJgF2TF0RPjoRZlx7+gP7RtXy5uRUZ6X+d
RNx7fmozzpKRvhrc0G5+FWDz9oFsqSeglZbs07BAlyVkqap8kqr2S9Ke19Fw+FeaEnNxFtE3xkw0
F12zOF9m64IbCT20nhQ+JJUwST221bNCtAx0G1wlhaSdVsTG3Xvud5xkvujjE0Yq18I0Da8UVBBz
a8uYUxbrj3XXAdI/U6YUKLgj+Riru5pvyYCIWuMHpEhmnTbM0yw3MAxiNfEV9gnee0p5HGtlztIn
RIjn+X8U6Wz8JhBbj92WBHUTpfegSpmqan5p1xsqeUyeoqmBlGn4Ln+Pu/6237hcKFWKfM6nOO7a
Rf5KzFdKT7R731wS+SSAWbaG+3kRHOxObVO0mlipRyE1Y2nH+JVN3Fmscled9IIhomr6RAWhsH6V
Zwu7TCZRDupJzBzHygAgMUXzCVlQDKMhqYYm+uUENadumd1Rz0yWyjjtNm1XunXqNoS1reH9/5w9
kn63tGd/fC9HpOvC9qX1Wdidpd7X0dcI7D/FEBQ2ae0WJj0G61FCQZJvSvsw5ydjKZw4qJ1a4Txy
/RXf2c+iqQ50QRk2JQ3CfFA/AztnjSwK7XvNEEdX+xBeK/Mvb0duqV7qI2SvNBVWQttABiuzblL9
sjCquovom3MI0bMNyMRefQfWeM7ADpyQBSn9HY4kVQP3OhUun5ycXF7jbQJvNhwxvjx2E0adcWD1
0JtbMw+CS78owzTX8k3E0MaX4P8rfA0OlYRKPhWYR57Ji4G4GRQmminh8lCdMnxs4FpGkY5e7XBr
umRgK+kUBxLgt9Y1CkQEVbRbGpHN0gDvVmUcfaXpmRrgHnVfkqE/gur7cg3U6YVrHeF+0u0oiXMc
tKr2IWg6VBueGvwJ/zIGO6ALaup6wQ2tgFW8pTfn+c9nZHYsMThIFuGxgXNN+2Ak5f2iJ6AoWLdw
LU1LmJJJ9J6symjJHWlMqwmxCRnM1zkE5Pwgh9jOgedtsePZdxRnLc9qSIKVs+QTTXf1gE5DEN29
Jhcivx0r03YBxGCg0BqYTuMdP7eS8Usx+fiyICR5FmdKjEUdhSUzReGaJ5kahuNH/kgejGmFaOCw
2n8tbQ76XLMWslLkwCyKQTLrQlvcM4RLhqPDKKauaya21vItUmlccKwR6kuVBSqolI/vVlTkkSvE
LNVkt2hgeY+LWfNzba8kyxgor9OqG0SP14G9F7JW3fVQylIgcXo1LNDxpPyyjbKKLkqd8hqGvjl6
ojb0f+UivVNrtYgsJpJL1eqhSiC+12FoJHdF/1pdATKZAKrTMNA+1Xfd8VO9favIqToKXI2JZWmE
ASll+9fwzoVtNhDA/SN18RINeLPTPfE2bS+rC6yE6zP1wD/ph1/PC1WB9XYFONaXgmuPVsC3n4Z+
jUtLjFEzrUos4BH6hO580HVgLPiRVRDwcgWlLeYCGuUbGVEG+mBqDcbVwz+QnOo7pJxVvZF1vhrJ
JxJknGeaD7G80d+KW4f3L7lzdLLfTUpDmd4hsIFs57f30YLbG0El7YiI/m+Ej05XVchSKAC0A2uF
Dnu+aNFm34gI0xl5MGsPbABecZDujYuZWS6l1OxXX40HfDOr/bi5nl7CU8M8p3l1nwrov0muHRQr
zobUpc6Q13NLoI1InfuHAGQK88cqEZPT6zmJuSZTexhMnZdNXBAX7ZVPsCErFWN9cfpESSmGBUBK
FM6ClFX4ch4dpsMCR+Nlw4XfY9D0VRBwjUhja3w556vTehfyV3HNlB4jSnIc667y8J0Zelq/CDEx
G099mZ+M9WyKYn/L0TTgYFh/0l01uR9yGEie6jbUOvRG8IEpTwdnAQJTrG9FcjdKJptAYujF82mD
8v1cmFQT54dt3ap8foNtPfelTS64Py0lmSaBfq3aIvM7bwif1Nk++ujuwzwVbiwIQzJZE1RWCNXb
CZqygpt0bFvwA8nlPF2rNgtSpGU+8GfWeaN9/m/rnAHDNO1rqyq5cppRxnPeW4IoEff7SWMNkvWA
DYRk3zzSeJmHrDQns+jYH1444A7t6wZM7ZIvUtqavIHer6PQ2dM1jJmyvMiMYyNw0eHaU4FCcAPf
F16HLxa1sLLaEITlDwOVT18/iwvL4BwzwFOpql2l2Enpl1Je08HYLvFBU5+uNIXRgWbKAPZCU2Gz
QOSp3mTyKyMoV5Fj8P6YzpSXuFb7kaD6n4lwPeCVwE+zwyC0EWe1v6m1UZcEGqfQIpXofdIIk8Qb
WtW7i6jLdaenRKZ+WodFWajIcptEY92XSPyGOjQFRklSoml5JnbfYFUnfh+VJsMezm7QHN9okxq/
SIS8aA9ycLVuzV9azo2q45qzW7vbwTtV+ey1i/R5RWaoyDuQwQS3/hcjeumFjrRz4DPgdFRyG88U
RtLR86ebxjejM2BMWFV12tcALYI7z9t6Sh98Kfwa4gVxXa4+R6Ev0HAeHl6UmGgP7b+k/UESev5T
LY79owl52loCfCSa85cf5VRrSVUDFm/Gj0s+iF1rVAVCOQ8F75bfIs7du/beukvX4wEGRsmmcCHr
6hJeqMMr9qG41xaX4DnMMDhxuGD1FThPXfPo0m1obB/EOjH/O2crW2YQrUSDwm6YhxE+UVwMkGoi
5CpRBarfTt4ocezIS091ODIRHM1QGv/AV9tlz46qDzsZkcWm7DClweNVhkM7Ta3Giob8JwlDElzi
il8+MaixnR1SKYfpkT2GcLEoCgl0CUmibk0lZyvolMMhtatKNudSNTmWVGR97DgDaJzjgc8gUYhq
Ge/1OpiWr0frPHvJPmegV2mF+9L/gHwMBZS0OwFKy7o4mukf9EBuwhFKhfhWgK7WfQdz52h6cGrg
orgS1tz5QfMPpcO2l++2xWocwf/2UeXnRm/DVZgtyPX/fN01QHnl60LpxGuoFFvrxzYTE6URxaPf
e5E0DY/IswsQKwmjnLVtln9mLkjUd+aa/BT8sRzHaLenKyEs4+CxzttNItOz3MHzIvEKoT5KmK5i
aKHxTibVgcnQweXu/X8MmL9JyQ+CsEfKaWnc3q+Br1ZVW0R4n5byal0HwqeaBGF1T5Q1qQ3frUZz
Ler/3KKCtkOCwZmdvl9G3Q0YxS6Tm+MM0Fcv6JUztU4Mk9+aoiQKqyDQK+miJLzcn+VkjWSyJ63k
G3pwjlCNpGSZ2tNGjmVd6j3Q6dsNj7w/OnPs6d6yZC4aARDM5qplms+fQ22hOwygVVtXvbiT107c
0E7pjF8LaO922K5p8hQcfvGKfI/KSeWDt17bU+8vfk3DCrBswzjZ3xTCVL9DyespK0t1md5earXn
+v5qACaRefbA0RDND3Q1FFlA6yi3ye1vxZbK8F1q8A9PJFN3GU5Vz/i/v9OoPNYD1GbJ/aLy4S1F
RTuk4+049TTUohiU/tKCFWWp7LSjHVLgimkXMhYxyOBfHEu6jr6zU4Zz0T/759LOw8ugpXr8elw/
J55QBR6IQeEJTqzMTNKSZGJxAj6wQGnZQiNDi4CRiR7cHTxBXfJsaBGvocayqQhVGtbF/AYCUVIK
c8vkFnr3jLIcSjdQd+9frX1OkYQV34U8iwXJpdEbmoTbYsWBTKFlvYnthVeMrDyXuoFE9BasKBuL
I4g5w3q+cT7NMp8go8qB+w94VMDvnvhmRYR4VLtn3YvEM+LXohRIKfsZQ91cnjsJibP1LXPvK+/t
1SF4raa34dFl/7Tq1dgXKSFKn7kGIR6Sg5qS6XEuRZf9/N1R/5zXLUlRCZuQqdUzokRU6M3qoLFn
G6hwwpP/hqtpBix9WSRge4Cgoz64V9XxWwfE0+IkrGerPfUcP/hFWAQVUNVL9SW2Tk8BaD3xKpgc
XwdFzMLpQNXekr4I0mef3yU/3v0M3Oxy8aTZ/qZGMU1EY0YwDhYCY6XyMlKR1+Jft1NN3expljuo
KqAk1D8EGnCo4Got1xKaT4iaccrhpcL6KqStS8RYhJ9KHStCppBydJDcRJBQ0u8hIpgh/z0xvk4P
yzW48TNRLqCqpuGdF1+RXROTez/SV4bkhdhacc8dgxk1aSvp0BvUUUjEroB7TuWa49BWYOBd5H+i
kcMKxEEwVQWH/f+lGutMejvbGROK9tqqVQWpIsXkJldhpungTziCN8vyAE+TjuaomCx5VHbDfqWJ
CjWdQ7Idg7+7F8vRD1ocL63GSE04lakFjboRnyr1eHD0eK/Qwa/3f1aa/vAEprpF0S17ku2zz4Xl
2XNGQBdKP7O5kSb7dSxEC3j1T00eXnZGbxt++Mp6t/QnpesJa39DW0OfnlT+xxSjhzSD/q+aV5gT
JgJuSW+IW8nU3lahtKEb3GtSfiTYwP+AoyDezIX3im5TQeigsIZCS4LujBRUaAaNk72f+GTi/y8M
wh6SNkPTALpKxQ5dQk2K/hJ5arE1/Ruge132BtX8+damiWcyGEPck3EHyBNKFDFYlsVBPH54xs8w
ZvV/D8yNTUWKxrcGSZehO3HD8jo0fm+ykvy8+Ddww37f8VUFS1m6B3bUUvKe7UqZylshY3QX9+yY
F/hycPzFNeCrmdbjG5EHpLTRsFlxRtdDD6vKINNCoQCeawTEB1HRGIUm6t5oJeW6EuUnm9qmmKUW
Ags9jEwzCLE8+JxVfzKKB74Uw2hZ38o0AiI0cP6FgUG9+5BJRDEsndN9ha6rFNYCK81E2XV9PDt7
pgMiJmwWz0ZJ20yq3ZpYBxlB/ZxuaJqsbvIpmeVdwo28WQviNbrE3hfI82eZqmN2Uh58oc1qWTI9
q9Zqv1PVE1PoIW4dZru08eZXfO7VwnqwAXAWELbsTesRva8uBvM3axiH0wHZTbx5UDo+8RpTA+13
LvUMXP2l6CI+E5RBSu5t5XKk6aPBvGUJrl6OkhA/5+zmWwVW1PMfABSSTpOJK0uXB/XRhQIpNE57
3GA8G49BH5HVa7Lj8c4JOMXj7J7fsfzbfGlmDp2XyCHkEerEKr5fVmw8V8E2WGjXOKvqee+NQYMF
FMknD6z4dX0q1U77mehD+du+1i4dgmiSQhwK/D1IBMKZHgTXCghKQOayA40sAonh2XnfID+k5YRB
dcT8BqeQ+cylxiBF/3NNGLTBdDg4/dF7PF1A5zooF2vu/DKVzVemNKfCnqPBof+ypDe6qMIX7EnL
uDKd1LZBgK3IRnnlJcprTs5078gW9mtjm3EWYtJEFbCxCW3BBI0IiLR6DIYmFmgGEKAfOwuQjlXQ
B8jn+zwRGZnJR1ymXrVomGMwvg0aECzMF2KMVsYh7wUyaRB5LReGLFwPWhE5zWvSlIwnDPdLcpKf
f8yl1ovyosoVkWpq/nizsehBiDNVTn2lECl9baIT1WpcPI27IEGmlB1DvKb9p8PqOYS6SaSuZ3hK
JaymNZWgKUn1s11NzvgFIGvLLFmX/PZwNYtRnAGb8s4p2VXAgWT5Trvz2AmDCLtCDvUvaFN2Sf6P
+chVJDBeA463qTlT7TnnbDJXP4UFjC4GqEq9Qc7UnjqwFZNipv8gEIHMP9J1fBhsGJqk1nEyuh49
woBaTerelubL//hPdfqiIbIUbVfTlLVBghon8fwYu4iCpqzEtHysAcKx9v4VZWVccRQUWHaNKE9C
gXZ8VfD3kKg5Upg/psWtck9R6Fr48XdeJrHczAj8noPtshFgIzJRLkQgHhLwEVp1uacUUNrqhf8c
ucJ6lKM4+tqc52LIxjAzRLaZXaTnHh3d6JYklqtKCBub/no+lrae4iLnF8d0f6X7zylabksM4i84
dhcRTYXfI+3Qz/ENK8mLg2yBPw1MP3AvYOMEO8KRC/n2xNClN4aEQTbSF7NKngldSD60yElma7st
ZngYEH4bINVwZwFk2gBW7uLHunWDjZktjHCTy5K2snGHLhm0MhqhZJcXMzehVoMitUfGBmB9av3q
niH+3kT9IGtRDBNfIN78nQDTdOv2ulyXCjGW5LyYBKlJhSifFU8SSEom6AKthhGN5IWb1NA1XCsn
YRw/iwAhRB6oAyQC0rQ+Rceh6Za/xOAz6YuF2t6XB6Ia53woVO85aBgRFEkyrgI9D53w8GB1Np5E
bjh3adP7Y7yH565oy27I90Pd/XfVU6SNVloYeyq5io6wXyvHbA3k79vbXmaZtginE9TZMtnX97BU
J5mGrY+HGlOTD9HXkjnA6sXICtFWUfW7WUkldIgVD+bgaKrPV+69XWUdQ8envXT2Oq8zqm06XQsG
Sshii3pWYXNhdCMLRpmxUA2mXKdbikUr2DcilIhvfqEDhJ0zM+ve0r14vWbcNytofuHeGs0lkJ3U
Ipx5R5Jt2rWSTq55RZi4G7W2LQmAZPVYYrEsGuarPwPmmiVRGUSFHbS5CGVvEbJ6nlTxSxY/yddF
KFVCSRpcF4ZhPzzP/X3utgQeNKlZq1dZ2614HCVGM08mc4d0E3TvakCmcb1YTKdGTCz/e7rr4TFJ
CN5QPMjsLmekkTrnwK2VyiTvNkJKs66s6lywFOpm2G9XerB2RLUklAn1UVFrJwh8+DOZKL9SxmRL
9msrJsAmHx0sgdWPUO+ycIUPnwcHYm/tWgfHXKYB6C9uhipFue1UvpNHJ/rBT1OrAFIRLKAvw+wy
pDSPKpCUzjVtsNpSFyXJWIUFmjMjGJkMXhV3yDHOUKVs57j6BqxOiu9pHRywZ9yZkMEJR4ZE27p4
EViYt/QAqLCKsV8c7JBMU8z4n4pZkESBu9UgIRQKHkHFHjsD2ey/abeNBAAbg03lLA4Iohdp4BEJ
Au8w0wUX9HBXHji2Id2gej+nWoCdQVyT9b6HtTXJu9rnvTMbwYVw3XeWcQ+yWbdz2HuOKme8BK5s
O1ysBKQpngYNaXLhO/MAVzfcerDCj85j8rMXL52k4SYb0j8MsL2IY/oEnhieu1gQwEbVAXceUi9R
cLs777bDwi/s5HuXjPMBetnKLy2YR7Z4xb8RMaGQ9qVWZWoMnnt4IILbD14C610HL9yBu/tMjpKz
7uMqTjvGVc1judgpDHkbmsNmmS5pDgjnJyhfD7z5pJQ/LsNj+p6feEUuz7/aNubsgdCpHNhwIE2e
NUDTmlbYUh1Y2OWWkjFyalMb4NuDTdtgZJTFlLypZV8bN4zcUIbUWZpiKgCsVsbheMTix4pVMF+r
sSfwrCqutIyW/IAIbtGwZVwszCTC9BYIVtxqyuYSycPwc78lv+GMRtYc8tKT66w/ZBlt0ob2vX8x
qk+K5iymKA85HxeGu7roBQyw4zCxDu8DLah/KS/+C5B97tgG/k3wnMD69rrcGr3wVCJaEKn0fQ6F
4mx77zRHL8NHY5vfLflFLPhmTNWJcjEtBi2u6NoeiS+WvADZGba8LObNPg0TLFbJRizyTN0suSMR
MftwN8KrAxpyoGZBZgHOu9Ir3+231GuKmHEuJXcowhtEaB/OcF3IoI/VBFt4TK1B1Wwrb7JeuYq1
TfXaamwKHBFK+PRNxx1cZJWKWJhnPUawejdnFQ0hdI5DTpqOihVkwMwyI+4IK8RiFoBhf5fP6kDO
7U0QHoQu246AjcnXGwJf2xhvAROCOKJP8jSqwf0uOYzyIXCC+ZpKG9TPhhVby35iNGeWPsH4ky9m
e1mIdVGe8xBclluDG8y+ghhZtAKUikUkw3BCwbxFsBFIeUAh2aQSsk2nhRsR25LuoBpUmEYLlAQC
uizGjFYYjTxSyPaqrjeYkhCN2iU5v1XKq5uDLVxwMi5opGG0Ae0Mqs6HLiX804Zpt0YDwrzAjA8A
B4D+5wLtTXSjMoLhqN0GTLDa4GHZEYs1CIwBa4kvgWhul5jLFToOOSPGVsjSpsfkWFOoCIiUij+Q
cemaj2dUwyXkXDJPUu6aNw7zBZZh9EELZhT5HCtUNVtGO3ewYhbIsucQ7NA0o8U2y6BNR4gIQa4Y
dZaC9aqLDcJVRD1kPvwohSMXabxJbxWXr4OTi0r1kG3Ioq+IbNdOiPtiQWMrcI4+wIzIs+Ka2res
d+rMla2/9biwmaZvPfOyL3VS4pn3noG6Fu7oDoYLpwRSxmMGMygNLRaFRtfbPd6T+NfzwJGcakg0
wBMiF+4vTluD6MiwPNOI9uqn3GcNwlKbdsJlLfalXKcvSmfAPcOYJSoP9yOKIiTNJOE7krJmaRl4
zRAz8Z9Z/UDsBYpoJ7XqE7QbI13esvh7W2R2FKJuX28moD60hxkMSevLP2oQm+qCQqmvM2WnhWtj
AhKWQqdcEyCQ8kAPs+FumA+uHkrVEPANZLtiW9OruDYrmC+8EjDmP1BC5iKGMotw58gqyFcuJDen
fpI3s560hLQJpWUIjFc4qoiWWnKRmnr2d1GkQaRDFH7K/Wzcv/T4yK/PMQkU71jeGIhdFr6X/bFQ
81qPaQ4+JRlZPbsuBdcPvUY7WmAAsi1KJEgQ/lXLMbReD+PKM8rz8Od3700Jj3LSSuzCV4DBhm+z
6/VG1ibftTMFWzqUOQ3uji2qzgm1gthoHkem2nLkYk1yr51xmMd9sWIUFuANxYWHGA0aIlUdE9gA
cfDYR+90yazPr2L9jbp3XCtQ0JuJXJOCGKxCMOAxU2F6yJXrpdsnvrEnVWFXhDvo9ZTlXVA8HfvJ
wNuqvbAE33T6DYO915KKRRJ/vHyjcQRdQ/7Y15BEGAMVLPySYWU3iKgcRdebKG3t0qvepUDL76J0
4rSYY0d5vZ/S5jzy1/9ldkjDAefXKsNc9mGdrjbDRKjS4wfKiViUD4kTj8kiNJworvFqR1NIMrwC
BRLO4cLAI1pyu+9Mimif5LIRTOhIYEgbJ0Rek5YGtXQuomwJ9OQWWmv6gEwJ+TUlepXFwNbBA3oU
7lz1mepnM8lOe1C68dUp22QTSf7RtwY4/yu9S6/yij/z/SnyTm+ZS5KfDbEl6LSizI0WhR5OH3c+
2ONsU5AnsDScxRVjN2ngH/fIS3oZVtsQ8pHJ2zU8KIafB6JNu8EkRSwwICwrifhadXgVCa+Nlk2J
aFISYKZyn80EkG21m4+qNYwA8t9Qog5KQvsu41SVoJIZ+qrgaBQzSINHrCIyClCMfu1sp3KquGpy
KBZEZUIEN4dFBMZQohjiefVfKk3JPU9/v2OC/306RbaguncWiVnRMkSgiWCc/BanNVA6MaEYKEv2
MZM1Fqdb4hZQoxJLf/6YuzcihcLa20GLL0A8oEcPFwzY5NAlIc8kS3hxkjDz1oTUEkXxlAd+UWPr
xFIIFQqhfWvAGj6Z9YwzXh/VpoheVOfH4AV264arGF7aRAvlNimOSbazRIYFTFXyTyoGpbGuPtNT
V8m5TVRFmAM40R9vItum5aVDfcje7PH/dXh2bfXxLuVIfuJPo7hHfAhzi0Q7GQO/qFPLupsbhPiv
ayFukbAC0EUW472tD+kwlw3Q773w+LZzxdoBP8XnW9vfg9AmGkVXvRHtPlreRf/MnmUa+WNq3P+L
fOhlOC02Uujlzng9OxfIVtkx8+eZdIb+xSQkVr5F3Z3CmMMsSX+iyfxEax1n8CJAzuwAX5FC0LkD
aIk+k4GV7+ybnUhxU/lMlwsAL0nInED/NVsRc0oU+LNUrhLh3FYW+xiwocKX5kdZbnOkRSR2tcyx
omwuq/Ja65z6xfohzA1q/TdYE34t3ejlm/1uyCMd+26F4BCrlOEKFNmlaFrXoB/gKjKsTsoNyaN6
n9eppwkt84zmtO4q4LOEzc6YoPubC/pfwhtM3/T6KVQDnZQE5R4rgm3gc8wzhYgND3Zg1GoYaAvb
syoYHtisc1XK+wdQKoSESO4RQfWS5uQWN/Hu2nQSRHdfhwnPnHwJXw54q2y5STbByf9XFVgd0oc4
qs8khILUXpI2NUTQeYBjnhgP96hUOb0vQtE1U097iwKb7tmJzch/4KSNHI6rlE3UeCnQHM+KEkTf
lVyBBBVEMfetGG3INk2iGr44Sd90iBFYPM0wAQH+yQ9An+BFzHW7k6fVxucDSUqOQnHTyQiFVFrI
/nwRIl/Gc9hjs1cI481UEFOAgrrNfV46F+V4QNMI3nDuF7BY2wxS5xdfxe7C08QpiNRzHj/YxKS5
16OUOwI/0EvxCO133qbhUYnHSiIcJpTnU/Uxe6xtyVEkjYs0bfHnwYZmU1/Z2gCAFOWc4W4AUMXS
ZO/ZTNkDKYu8kMVSk2pN9pJ6E9ld2myPxyS0BXa29yO9gVchKKvNLweUO5zTgFgeSKpQmKoPEFwu
3p8AXGLNNJiVoVx8QXSAUNYQ6YEvr0gKDth/Q8GKdkIVVAvIrX1I913J4dj0d/mA8kR/v28gB4TG
ZTdN9lo3iaz4bJBFiv+8vbJk9ENBHelAe0J4XPF6wdvszfI1LOBkIc5NmBQ2YM3NymJQRSZPqzYf
5CbUUO/bhKbOsIpqXafC9Fhv3/ChSWmBzfnWsOgz5/2SbV6ZNQSfE8j0SHP/fYrvjQ6b451XFgzg
2shT6EWj7PijtRX3/bL+q4N+0L2TD7z+6eaARfMQhwfIcZj7jUmbmjGSvEeJummQCqV0a3Rh7Zz1
qZ8KdsjPsCtYdifD9EKjyKq/Rgx9W43EmXmG3UXpuy8AcUanxQqp4c4LMXseBGRiwu358m4/qP85
LEDXeAGMJrGWEV0NECDKfGkOrDHL2Sy6BgC6xI3shZrVcFBVu8EY/jisuXq3/ey3k3pFI1Uzje7k
G3OYg4G4b/SZY5CJdNN7Jz5EQgMYjjx/1BBLLvvYTGxJxD9o/9XlJXq5r5o9d7f4GsD1paL1Pfui
2ne4CxVSybiXSzqChG5Oj8tw0S2JmEoY7UW+0wzR1GcDRZeb+8jI01BH+rsNpM38CsxO1NxwGODj
Ud8dHN62ZbmJ8NZ6U906zPjbXYn2ZGmyFd1/O8meH7THVhTHjaNeO1ETPYGNU6cGKwRDLSirkRHP
Hi6yBvWAgejWDtPd2LszG6/53k1dBcpr0EdoRI8FRde0Fh+Zhn9EV9To7azQ3+Eh9wLNFsSWGe8c
ME4KgRn6ISqSVDScmms6/FZIhdKpZND4tJyf/CwNCwKLbKB8Os05PNjPo4gIH2/o/pG+i5zGpWan
Aa5Sabht2SB1afzXnAmi/ZODe5tpDgvn8eztSe+Hmk2T/4bMNFmSfpZQPVdNe8R09ev2b3yDb2Ck
GAT7YF30FcmW1l2jejG7hyPSqaGZYe0s3Ayy8OEBeI6PmmKCSUkKmf9f7OdViJrJC+iRIB6whabY
dg5iRlrH7RFStzRqDfQgpy/UxZ1GD/ib66EGB3D1We2I/qgsvgem7FB6h/FAt6LbV1w8jHRifqic
CgH3iIe4k6VDG7DAW9TwEccfe2retd2qZKl0oCLs3OTxuVtt74w1ZUqGx0RJbWKtTDZVruqQQY/P
QmWUIFXTuvXwJhRgtn/y6K4LMAlUVeQefcy1+Eu8Nwmdlo81SEYPGnzkXbHjqWi26n0sjGPHc1gU
B5KjtYNPjOUJ5Lu86PZFrW8JDAZNxnuf9JqhZG/QNnAbgNsZZyEKccBU4veQddKdaKnuTuW4NIyR
Z3/5G+Qb5yaIpT2nAObrtk9cSm1rtAh3Wv99yjafblKYaR/9njIXRLyM8MNCVwpFRSUcuxCQnYGh
kyADx3yuD8ytkaN0yelDuwGt6Bgl38iR7hOxYfgjLETYp31+f1kLDSMeEeRW+JOz8TxmRP8iivG9
hBTyA7QMqTvYRpJ5seuLh682Cw3rKV5mkt0jxPt3FoZ2fK7zp16u7+HdEhbV9JP4RvqqPxT4XHmT
GT5Ev2NDaa+p2icov0GgCuxAv+XSJpR103Oa1WYljZ3eYaTY/zJWUmbneieJTFV5JCEIPOFIDMd+
GuI17avam1tsJI6HJNQagTV5HAbncR6/CGDs/q5V0P/2zuK3nZ7rEv86shz4+o3y+bRNYYGh2lxv
RAoIOJGK5+farLXdicLmLqfT7jWGL963S3bnQeLRcFt6Kf2LcCGEVJQm62hUbEMisYuSpFRsizMs
TmHf1mk9WR/lDWIXgC/zFGGQ2rQ29reQc9qm14zC2bfgMTj0BU/TY89rscW3n+3ppPd2RfOvft4T
+blF5MJfH1AmrMZka7JfoX2uBtgYy8+jBWv7srESVzJU3nRX+fyxldGjAfvYa+TAFfqKarh8ti63
1Q17U35MnuMac2VBss6IOE+RyOjLNcl4wTRSl7Z5s8A0X5JENZXshzZMUDksJLtaYblM2eWkzA+x
pdBn4EVlfsD9X0Np5yxhXD3v2mFGb9poYBEvesNxYl8v/AuWfGB11d0gexRHtDJsgXM8bJmrhxcv
B71CvomV/CGdMT3xh6vwaVbxmTT8QwpLIWF/RdIBWu/nsiMeROdeMFbMZGOm+N1srtf9sXt2NXiO
BgmeIhx1Ke6vFC2y1xdZwSZzAJoSxPV9J1BFuYkouXwwKWx3nuk32g9EGcmMtD5eW83FsrQRLIuD
Var1AcVhBqlipFoLxXfIYYx1M5c3PCml0dYdQTCwys7BWfP968Vj2dwvFTmoGVyk4H3700izHgrL
/80rJWsS6qC96QgfqJLfoBg05K2EuklEwyHeoYQ/ZYR5I6saDM2ShcuEQO7HysFyQG1qQ85stXFk
Pyep1vpQn2AO66m04S0tArGcVF8hyLapvHu1cOCfyJfktzqD9u3bLzPTsoq8HYT741/+zl4+Hrz0
CfTYb677baOBAWqbXuQ7XTKx4SPjaYd7vI9MEgK0kFcP0clQXaqrqqFmgXBvEtmZz4ecPsxriJcJ
bUaT0E3Abb3WL9lRlBt/yzeociRrrlvkp0C3Jal2GShE3GOs+1uxVS1Ji/cW5Oi9gZ7fzJhPrJ5d
WyDyR8I3wG8L4kC3E4WICUNtiqdXPycId0nzHQdgtgpSvC4luhmbQdHfiUEzs2XVUuaaami893qE
rO4LJz16+umj9bu7gf1dDRkQ6ENjXsCUUv3b9/lX5rHUadC4mRjYNaYxmcs54QnUNBYbrjXd/wCc
E6STefw+iO68ejaTTjMbf0ez+9occHe8CVtBNvQoETzxCIfw/hoMx//9mZi8wq/1kVtoRy752f91
4iny4kAMkaWPeNzWuXiQu7p0uwSzWh8UbBOT88zKmFPZVTIlgrpjlWSDcSUvhStIAk/KEZWXs3qL
cCFvAVWh7zqj7jZQCzoo39jIT1CxLQa8YQlh2QYMyrdMIhBaVzjExu6cVRnfwg19nrJx/GJjyyOb
QPPCNSNIYCKtsHVsgpyk4Dd46+BVeB4xPMDrH8Hma0JltUB3fXeEfKzcfCek0X+DOI/Xmx1qNU7b
pZ9yyEsu49GU0kBJmVSObiBnCYdfxBef3xy5kw89zHs9Uw8EvSuqap/clChQf6xRmVuyCfdqtsmW
TVmNEmJvLc0nPAkdQX09eO462PkCLDCUvAi333WqNgWgzNHOnZDeygGyUxkq8maT4bzk+6aazVF2
vMJeA36hFx8ZjiZGAE/bkYZ3EI3NFHPS5FauGmavXhvGHTTXhOjE+fglsgjHoVXkygfLCGkfntia
JnEUbquEE8lvayCaVAt1R/p7qBk+WG6XX5bh5e+0G0MlmbTzup6cYqRuWIkP6wzl+ASB5CQmFpTT
DXz+7kZpa1GZCcfAQFPXJ1dfzQhJZvKRWhnZw8f6XccrRY6AiuSVaZIcOPbuu5xjh1E2m7x8gy3B
m+HigU0HaXupnDjYSJr7MeBkXMdK5VBfW0PBvSrcOgnyjkt5wHGr1Gy7W1I9LLTy17v11sx0n7W9
gVWg7eEph2JuLWrydVnLDuQKeY4SWgnGnWhbdUKJ+A7uBX6Biz3ppclICMhV3EnoVhQwjWlBbgqh
rvdi7ZQMPQtx3dcpEkVyJsP9iK63LEasSbry4mxqZhuBuU/YeuaOb4jo//kCEO/kOEdAd4IWzIwI
nQ7yhM1Y3ITYU1OgrGPfwoc0svkZds80imS7TU4frITcgpLWyecfkiR75uOovSPWHCkYYkb9bgjC
rPcn4KbMgGRxU+aj186Vtno1HogmTnXm4Lsac/IN1mOyhwT3s9gv1Io0QVKkSROS2oJ2P9g5IkOh
xmf2lYUOzckju0lmnVENDnPb6eNdUoxtoLpNZMiaoHNvr0645LTnG0NTKOu7r09XEN75oiIZtS54
93h7WG3TwcQ2jhBAFQt7okrHu0iGCRfbwP0MewfSbOcqLJcLXGq7iYI/nO4WkU1JQ/R3nrhH9gSz
d1x9qsoiaaUXwJ4PsSd60VFODCeFDpbmG/p/iMfsFnFcKkNR5Rcw4ZQRRZwZTATIubknFZ5mbecP
06dYyYFl0sGvb37NAspsWgdjbueiDUD9HMYXTwOJ0ApqZo9vwAC6EOealAj1B9SJgnC34tDl5uSI
6O104nKzaXmBZGLSm7UAwJv6NUACP3/zQxsaJg/aP8PecgUMEFBKNfKfUFYeCNBWfCp64+mq/HVK
2dlzWgcd+rDWXg9+SFTIsl1Uc0EG4+65bvJmdKaVMv0MIPtqL4h8/tOfr0cHjT0uJFukTB2nETmx
rsUvEyYGWwFyt0MB3PnvKswe8g9K1cQIpjSJEvGvdVZlLG4sMkb7uMxRqcEXUhmxyfPo+PthTXFL
Gi7Aw3bgR+Vw/sY1FZOw8VtMfHNdmwhtI3+iQcW7Rfv0/M3enc3xpu4DEzTzjr5UwPvLTSnWGAu0
l6h/mKwuM0M0agiE+huggBMJ4/vdhSWFsFL1mwxx2vcNfFewKXOQxR4/9v6Z3mSB7ukfUIMcH78B
tb2lEoeELWoSBjVAnZkGw9v83+wjLGTl1dULBzr7Mp8XgN/e16A0zsR8BFf1OzzB0w79sDalqmC4
bVZwLCxq0pS7Y5cGgko1bcFXiv449juFUCMYmibFmOHCOrz4AwJ9VyKYGMnGMiplfqZY75jgaXfA
dj+rlGBkxQaJleCWWarnepfTqdytQsHNx+3lcEN6HA8ywvoBj4DIfO19AWyoj+cx0yCL00i+kaYr
XC2E3ISXfjhv+t2Dr1A9YuR4vKvJMGVKvmF2EpmjLDehCbY4wnBPp962nNZRKyLOqCOk4fCsHtQS
OAhZtuhk2lr4Y//Z5NVSoJyuWx8Z5rxUuWjOK7Mk16WNmFFzTqYmbgfWOSossMDjQheiLC43YBuQ
2eoVHgz/Yt5/GKrdzTlYoV76y51SnKjjkLcrNXstWDoe3kXdzz0JIWa6z/BaMkm7Z04ReNcwBZmh
3pb9V5wOFL1fcQKmD7GR18T786SyR/Olbd+zZ0XSoOoq9I6VEgCvAfrcSG2GY0ZzmBlcM+iZsZVJ
fEeo8dmpFSH11vsRvkbGDkZ0HHj3FavtOs0fs+TZzjcwOI+35POVgmfAdAKoZ5/as+ixagWeRO89
Su6AkPLDn4posjcNfibvjZ4IyahMltwaW+0gKoQL6Yc1pxABexe9oD5k4OCcZyjSw0UdYSuTDvid
j5Sd/hPxouB/j5OzXufjUc4R6Tgrp4OmGqiRwhJO4+lyL22JjGscdmvsIMuInEGFjhWgrB+5IUYO
w/cDZGvazeD0XlV4212wcpzMvF+7H9LwNHJ2fw1v+fdAnLFhYV3o1xuNEpu6vSMEYW/32x/UroQf
YBLyP50buvPUTLgjUHt2/TZY1OISHRwp/RPbxKruzzrqFduXgLnBGK0PbPmvTgrzwYgYfRb3eEmH
KjBwYuSxvzqqh2i9y9IysvhPJnMiu4cKv0udJTKEiemk0k2tElD0bZztJ9tnGP83IU6mYKQqP1/C
X4yAfB2QIaVwPUMiF7TauvUVIKQksJIJlQBkdJlA3AammpR6yl3tX07BRmevVChBQAVkdISJnJny
FSo31bMfZgSbuhlTHX7I7B3ylbODBjIB3coVyTJrG7fL9N9F172yaqpNtxJLs10MfpgA58o6rAlK
sWGUDWnv544cIeSlsjJRrMrAKQ8scDVXdsuqjVTnxfLVs1xbRVprLKCsRO/DUF50tRRu0VMbHK4t
HhrTUd4K2nwGCJn96jCA/1/1X/RP5aMsm9FTJb22avKctTHIMtSBGSg57mYoLGrmCtKvKkQ/7vRi
MAjvsNbwLGCqZwxA1wRIFPns2w1pgrM+7RNQRwptEPHhi37qMAzGYPOCBBCyz+8oBuIxh9fTxhmh
M83DAIlGehewgSpbRI5tTEbmpnSh06aPt3itkbSAE1n3hB22amn0pcye/wTocRYVsMnJEfVUX3pq
KEWuo/BwRRnOUTAFlb+wpNYop9+tMWYiB8IeN5jfwYTuP+xkyzdiFeCY2X7lMvo5mK73GHhE25kY
mAE+yUx1HuFqNijRVrFJgcdbgkuvAi8y77Lm+FEHO9CIkjM9X+pBh5RXkp6pyQVAiiKLznADZAoS
upLy94pxd1tFp805ayeZQeTLFhJbciwCWP8HbZFgLVnZc2Y0/zxTiGOgZ1bvEChXBMvQyxYWPuHm
p6IYvoi4pN7KMaJPhTtG5usmEscWIMsmeZNQdiScSVVyb82RG+MWVKBoRHQBd0t3aSwFAFbi5ymL
qfBEGcfTznI8sFOJVR99rJCt1GX3UjH0FcEL+erMTg9XzqAKLRQQooJ5nGzxiknZHsQ5eBUwW2Yl
BVXxSlDjI8HvMncc1MvT0E3sXJA7oMCTgaH5mPiCobyWWrMjTR00GprJYCJwST4NjFw0QIGHcaDe
eB6ixnbg0HicjxUsuC7binCOpgO9jX9ldrAtAd5TSuN1Pc3WshZbd2jwTR2RtpkQz7ST+f+t1//e
8VEFV2YrvKIXlIB6RWXZzMhitFkD0jiviTwxTLEbHXyF5l54G9ks+e7tDx+ySs6jpFlg0VbOw6b3
xIb6EKKWk11oSH8PzFeBvJYBVQjOrXEF5U7Sm02ZVjWqx/dvDq4UhERMEFoLqkxl3vw1UcC+/u5t
dtdFmjaiPkImRgAlr2FiaeqnLGZ/c2gIaUpvi8PTlOHClCrNiIRfQ2H6BoC8PT5i420weJp8iJFl
4QitLkVxgVBlZYMgk1tSijxqF0Bwie8ECHh/pt1gQ17gCX/yu7p/B16Ofg+bDfsFk8QJgm73etaU
hUr5qgmzfmepw5+Eaf04VNkb77USqCtfAIsxm5HNEukNX+EvBFk2c4asTlROOIC1mPs/bKstCc/e
VgA2OZYCx+5L8ibOxcClxKHsUUvM8l+j/CSipclARjZ9jV3aTk2Pt/TVuUmdcLGE1Ll7FeqFTfQ9
Zt2ZKp798eJ9CT3fs+JdajUR4j0b1X41cQs+7mtqniWPRVEIW2JCoWHMM3wYv38pQqXCkpC2/OFd
WR8jRFVaIHwWwUccWAsjVzwKB78jZfTEqvt5y1IXpLNNpK1CSRajJiCWXH0gVF2o/HZbPdGjGcNF
DuRwH19E/af0PkzmPQ4xMClfIfhE1LDYfRfZ2Dp23mNk8WzJYk3R+iiP7CefdmhXaGByh7TBc3ar
/HGgrVXrl7+fgvMk7gtoTdu8tNZM3R7TVxdEWwusZRC3RWROhpVhdEhnCmnyVdKv196DLI0JKhxg
PgBtDOJsXLbQkZ0Zsk7bqCA+A0JcAl1Q2nxJagm+4HWUpn8cZ3Um4+EFlmI3y/x0i62EkeaeeFBl
uPkaunAlG68Bs3VNj7I9rVQXhJAquXchGXUuUWR7Mz7ut10HsbZLzdlHF8UVSp/G/UvSLkW2xaWl
3NjNhDt/jKxYJmH0uUhA63V2olNtDyvkNrmFLUYatO9EY9JR7qpSJwxtZ1jSFR5udevQyabW38xA
Vup//q/EaDxgP+aQI1qDPoQ+L7+16aUr1tDBztDeuOAtJAkvuWOrXQpnUwwRln2insCznOC4nLHU
9xhJBJyRfvtt4XJ5O2/HmtXDEo/J8g5a6RZt8KBpcjaGtsBVuos2JIdy+Yg/Y3vnRBhpc3M/5oxY
qAqmxV8iHfT/APiG9Ko/XKHq2h21izk03twuyJFKdCnG4hTVvo/Vcto8MS/jcyA/U0j8wT0TBk7h
hurMnS/gBJzSXQbYuEyosq8c+Yh7D69s58vvbxyKU2Pr63BqwWOm5z+UlJZbUYa0XbX1FnLkKM1n
UjE6hmB2SVzvX6+U06hmmBUb5UnYT1vG5wfLVmau20giW+BScZ4pcVQoGHyb2ZFa4xvjKVr7mXWe
9wuQUZ3994Vt9xW2L/DtTfEWYK26cNIYMET5s4ktdNbHBLJVg/I/EAD74lho6BJAOA/D+fRbCnn4
3tHNIZH7uOrbIWGzTzNqSPXhjlbiMJ8N655gLdp3pr6BcmMH0luVQET+QoVvIY8a1xAP8GGFALNf
/nvMtzvAHgmHKv6ZaCC2bAaQUBZpjDeAqVnQiONWNXDB/TiHeH50Dt3GvGh+BWt9YrEeZYK0Kkq0
kWNOwjbGC5IVmXSdW7lPveqgubTjbYcwnBXszSOVomF82agDEepOpNaQlSUdJ08ezNJbDtTQ5tTJ
umyjhi8fmZamXW58P0X/VzZi3iAuZEq+YRDF5ReVz3iY7504TaUcckjgBZB7OadkIcOyMGM20SCG
6WDq+erpYOIkZDySPLdzhnB9kiSsNlS+qV9AcsuJosQHI9ga/EvrcDViUWT0avyuL5x4AODoXj53
Wqrw4ppDL0xaRD3of1ZhchBHq2bTdmXMp6NjFJn5aFGy5swM+SbkJgBtRMsYXYfzxyYjgmzSkNbR
P2lGTK7nM0Tf7t46NfLJQgimnRy2Reouc4doPCRr3tiGre2L7J25kk36uSF0iM/lLKyBBvMbr+W7
U2kDuJeof+ccG+xNL/JhA0uCfAgdVN4/TdFmPd/POqmgZQScDZpYuOWlxN1WS+F2Wi0iyqSm1gZA
q+7HJ2OahMIBZ2oVNZJmJADpi/XbZHCVa11eI9+7YEbc20t6Se8bg7jf9w9oVoCytN6MB9CjalXH
VtWywwz+PqpZwmxmG7o6ZSQhsbAMJ+PaZu0s+cySVWRxEEIpK3tgjPtGUpBENmCgXDoMXFeX1eXe
KKlnu+fFgTuw63We2/s0zA+KkNHIB8MIE6EHR+GbK/5kL1jYMJ73LYzajdQhbJzSMYsmDMWwL2YK
QEug+USznTsGTnVAq4TXgdpaYMFfMAl1fFsw1lT52JjW46q4cEy59m4kJSVAx2OeEGXnofjvqAKl
Txi1URpA2ey7niE+iWeuqx1K7jmAHOI6cJpeWm3zgjdRuuQp3Yfc5F0drtftlesF58SZmXjye5mD
f3mYpOqfpOmoBSfNOLhlmuFiVoLKMh7U2D1FI6A2s52Tw9pktHgvlg1tkSB9UInBMC/eNsc4JaYP
hFitEray/W9Se68Ocdrs9BI9C2WslkqGyizxVF4dbDDeFIR0E2+DlQL7AcXj3fGtyIJeYz32WWCC
pIN43HubkFz3PA6KFtbGSQTCqq/aY5b1deCTO6Yu06OhMPLFfawuWLRhUBUbU6kDq6FQ+jWRvboT
YfYy0cZsazmlK98nzDV5yi4T6MleuzNjoxXwJPWi6ruthw8BKsUfbdn/U74Ny6OZb53/Fn4lsnF4
9Yl5sG+mFNe3U+bpsQN1jff0IYPmZtZScSiZOCAoOvM0ExU6eMbIZXbdxZnm1uOQpD69XpFyBb+8
5fNa72X9LyOVsuDNjFHufB2R84TvSHi44C1D0PUt2NFnG0pHW5yHnj1sQu3F+zSo6JTl+j3Riqab
c/iy6J9I17U9fepW8Q8BC1SPUl2cFsx8qmTYZB7NW2BTDZhvAdoUq6tYqIjNIlWWCEM9sPreFU+L
DqJEqqCchbGaSADmnxWjiC4i5u+BWitqPYJ3Y3uVPUJyw4ofQ8a7jwL1ah7DhvcoIbnUlp026FGf
J/xmeynv8g1IZbjgKZTf/eyA9OkjdeZ7nTf6Wr3LxBUqNx+zkQ8J+7xAWQ1ElnOr5sKSM2alheJl
DSRXZqP8kLUWsL6gHnnHAxTqTVgjLRVyXunig8dAIyev1YtWXzwDfR/eKEPd+YkCN2L3BmB9T3X3
3XeVvMDeNiSE01OAUzrB1QsaAYPRF5tgKixO4IgyC+wgzkx0j2ilTaV30KThVkyNjyOYdrwvgX84
FXNyLdrp3ibJalg0dK8StfN4JLkwo1NXvR2AR7zWwlH4hdE+mdfBel7eAsaQN6ePay0hJrHguw5e
jv6MIPZhDzmoj7Hvx8bggC4AtWxtT4lDaw4LGRva1Ee/HgRWK4WyPtAYwI+qk3ElAjiCEKWbxTF7
SShDMR8NtR61jrHElvDorCYRwxr0xwltkIsQoDlmCOKp4dC/qlZ4bRsq0TbCWNsT9c9N9fKCDla7
l/gIM42fIBEpooSCi8JRw9vZ44YebxWBp72ITeFX617eko9K7u6TvAmAlrQ0d3twwXpEtZ2KVHpu
g+FL71pjRJsGLx9yysoOjgZhU+Rih1IPnF8crhEIY/QpUoHxunevWdKi8jipCxeT/lzZqsVPLCS8
t9Upmrxazq5DBEvGt0SHBUOVL9UDIe+MGSdaaJbJWMtN/YsHhkp8S7ngR4Nw6M6i8RAyW7ynfoHU
vCrlXmwhtoqwobxEhBzpWvuH9anZAs/ft7fhx0TMlOM/vRhu7SmIkPNKVqrFBntMY6edK+EBuu0G
1QAdoXsUQ9sA9Qk8vrL+ZNcSFrogen9skpApKyx36zDaUM+q/TG5RRXaB2YiYBFypMPWKYpgpiB4
n7vh65/ERAKagHOtADgeqBdNnoxgE4rtQqcAGmtLcpXc4uv2rd/bkU7KuzK0U2SsgIUDiBAjwkZs
hMwQ3qvaARr8KNR2HeZpLjiwy2UMBsGXlLdZgexGNw8oy+AhZd69d72a/kmpIurdOeNKXfC0mOM6
9srBCcxZC7MT/Q9GL9aQk3LCD2tscqMDWueL6x1nGyJMSrf6HJ8p+Kb+FbHGAcbHHpjVV2e938qE
9sBcTt0L6aa2i4cRCKTwFrPL9txdhjN2ATENzNsJVQ4xc6XmKwsqUwhfjSfyZVYL+Vz1MN7+49Kv
IQepLsBD+lC7EnUcW9YnJzzynl3XkwvpS3fLXxvXcUNomb/WFyIqw8dIbOE+pLiaPKaa9s++XQmt
cp53N8YTypjJkDTRP7y0OvgwxR3lQXiLJ34wLnKMhntc8v3mRq+VK+72MwBNz9RNVtR2MuLB8RV1
mN+7C37z+tSywbBuPkMVvVKwMrheYZry0LEsHNzW1kiN06/sTCeOwpAnaSA/suRjLINnhZ5QYPB1
nAqJ3X/u0IY/CChKGaNPXMlTYbakv4Usi6/udoD+HhzXFdokzdUnCEUjWtTMWWJovLBBscf3RTQJ
rFBu0tyAKYjUea8z6i3HxRG0LS1zo84DiSVzgTkOpOEzMw5h5cpsw4QEQ6o7jwln6dj+H2qx+I5/
t8CFr6h6cG2RidnCSp06TACalV8rODIXWGTqErce0cvtBiL93H8oz3AF1l7o9ZPwdadW1+cG7W/m
uM6PMI1VAhUPSd3yCNKOJAfrfzDPN56uj5x5ekNwiiyBOh0XFEJ70Xq4QHzhpRgDY4AEPB1i1fBm
8CWFXyzMNoLBa4XM7jmwAmAJJvQVEJlGvPyk0dOg2COvDrd3ZwcQhwWvVBOCVVeaQT55v2N+1BdW
2BfLSHq4tDF/qPyGAo1h4dNCiSYz8VRaF9PxBGP/6kdQO7YlNQqJtV2m2Vj3LIZ6UiUY2CYeb9dK
M1YR2vxvzyOSA82dYsJsWkdWqwEjhBz2RgZttd+PMBcr9Jo5bYl3WC/w3remXv3X6n69v/eFzlYa
542kWQA4KQ+hnNsKlGTsFmHI+v51kwhIUSSAtTnh1jC+NaERQBzcuDBdv9KBPbdaMby53dUlnKIQ
utI+CzXxTpnRzCDLURlY7+md90KBMdJaiecI4YnwS8APGQ3igLd9UPxTkstmnF0udrCrcsLKGytF
Yp+O633hEyM9/hPlbI6ptnjr1Dl0Sg0bV+8hdtgeXuI72Ep0YyZspP4SIhTptwZ0EeaTQhF0+c8C
mlpmRU1/9JN5h1FUhX9GmqfSxfX4Zkz0gKvqedkaUjaeXFysxHrHYtFvxn7ocTECLcm0cB42hKG7
BwsHkVyvxX6hWXBNijEAQLCQbgR17M6vjtP85F9BtVbnfDmebTqxFV77a8QlRFDHhO1i0DG+0chi
IoHwbAOGTmStjsq6oUQOUqZAV9Z/JU4Aeij1z48p5h0X4d/nY14E1ctk/mndmc/DPMGi122RtKsC
0zOX4jer/rsM+dBJ3m0iBtfDdXNjDGvlTNpX+VjDCKhcoMVyiK6dP0eZ3A8iTlteKRPh1pZQ9K+e
PPe0hEJwAnTDj0ZugPlvgzE05ePrfB6ATvHLUeo4q8beFok3kthyO9VoPpwZ2+lpaU/0Fbmh51ap
1zuDH81A7+Bsdti5B/ibjuiNoAhBFNinfMLU0ODsrFEUSIBs7P6KtWyXfQTIsmO3MQmXymK4U1hK
S8IxhS+T2a0F60HLj0yUUlVZ9OQcplKIJxLs7xYqOCwE+lztFOesFhWwO0ljtt2CJ8de9C1/LKsX
LqU7n+H0UVOEw5Kb7NlkEJOBjxNRurCe9a2Wid7MC75o77Yf3+sZ9S2mbaP2TJowLOa0aUiHp4Qm
rCTZZRPUJp3wZ5FUJS6G9xemp0Ty7RUrBQ1o7iCn08hfzC3vYdTcWimRZAKpueHLU2/mtlWoWIBg
Y/UUR+MjLjJPbE/x8LMXRT/IUgq8/F6hWUKS3OTxGBJei28eG76VlPKLRbl48lIc7xq5bmv3vtDj
rGbiZ45CRlP1ZnD6R8PWbAJY4nsNy5KCEy7u64MIHd3B3qcUG8JzH8SgoDuNNya4hZd7W7zeAOHJ
2ACktwsHjnnw5Ub9v9245lc6+ztdlGEjEpSF2WnVUip5HgutqygeQkc2ndtvtI7cK6DwQYLrfdSP
oE4mGk3qYTFL4mPY5qxnvYEOEPN4D3EvWTm9DH8yIMoqdu0TOiUPedr3CMSQDAtaob/j4nres3pW
OQyU8BYO9bCze1ZHRc1QLKLa9benZzhTn+pAjX/IJWF/jHZvcnJeQvsZ27DmZozBFouRSGHXe8oS
ULbpGVt/3UyTmdj7/bQnBSNFTNEuBPJvdttK0dFki0doY2gG3NtwD+99tfLPLmWEPa6A42dW6kG4
qV6O10TRv5K8s3roo/OnQcx2Nmkpi81EBZbnfZqODN1k+hm4QTqhHYvYEarqLfeL8SIo6bW0g+xS
KmYUNYoQ2GRAvsLX2+4FHOoDgXSmmYM+XNcna4rBzGupIhONqVxhnCXUk6qQ/3Uo2LAQ/TTH+xmt
PSmGhPa8iZdxInmNPvg11GyZ2OHs8F+/Cv408m59OtS2D9WniKNmgQIa1IeWKZcYgeuGJ8/ADU5W
nf/WXTcqaqHpMiLubTrgAlT9K1fT/UtkxOH1Aub9tD83DWzvZNa6e+gVMNR8275FMC+tNYlZrdNu
SGwzw2Exs7WduEulm3EM4djrzp/PryTo64jvynoOspV5GaekbpaYyb+lxGNu6L6w/LV9sHfFZmEc
lGQwbnviiriifkS1+3NaRvhhQgsZ42/oqbTADtoh8lf0xCNEJwyJZkQultFvLpj0Whr7wvHrbiK8
4U/tKbxXTF4BXWieGW4JAnR1a/wSF2RGDURkuB2Qg2qLyhfyhZqiyp8tVJ70F/J+F4xyznMKXiz5
XEMRg2WbN9XNmdloa7OWGaDJN23ilSA6YMsotp5WMq/FXyfKEq+aWgUrIn6T0g8OJkPNSwC/RopC
WAOQXgN4R/nwvf/wKmqJCFAOL0kZEW3k+LGRor3SD1KXyw5YbLFzlnwOYBn/j2NN69Byu6MQ8HGo
dq6OcAS0yMiP6/msXnhIVBV7NAaFM8D8gMSCQoZ+DIJ8/nidGVNS5SfRFRpBUhVGn4KeSSqdkhjA
/OLTRkpjtAEP6mIfP3jQ/s1cX/Fl+K2PWRtvVB4/Va+w0eIsTk3k7pj2mlQnVxpw9w51+ju8UgdF
15kb96cZGszWmtre1a0DDFO6t1Ey4rjyrK/KymdwdybQVX3feZbQx32WVnFnZfTCL9KYwfw3MolZ
WYmDn1vuCRcVGPm60872935uyatqT0hBnv8QMRV9lDu61WCcHmkPxKxaLAvimsInW4aZUnNGGU9M
u3b5blkZnJ1br/J7HQcTHlN3NyablNpkL0KvnN8Bt5Ih/oVJhzm68ZCFmk1udaYuMk6oI8jamP8R
QUxKgfbv7umg5uv1HTHGckg259Qx+XEL7s5Dqy5WDGqdsVnnYjS5ZrDN8NZTVkC4MEhmNW40F2uy
U//fMN4z6kn9YhJKgJWj/L/s6gi5U/kKsGGu6O/ZuN66aLZgdwQhpNIBAzdrejE32SWBXN9/2D57
KdIP3+SWNVIeon0OiIYuoBFJhLeXYW6ymuqolB1Zx91naoKEybNDMuEQu1LbHI2+LmIaJi6iElpx
6NjJ0ZxD3EX30wYhXp+mHgnx4Vqcnj2una3r5qsifMDvHQD0RDBlmPkwpY/Kmjo7dt+HzxEI31IH
IlAYOdITLy1y/g1iKl3UcB9sAVqbe1pS8ybNep7RWG5SprXSiRzRKWLtk+73vaaW/vKpg7RvBNcN
O929fqbe2GbNAAhctTaKr5cEPejER84OSn55OY1af1jp13g0ctiVKNh0xZHxUhSYFryH8y03v3En
nVSt65PdsAl6q2wjEn+tkBZJXeKypgQ0iSc0FyznigshzvMUHPJuDIsQw16ST6btQIcsc5rmzoNP
m48Tny2QBBJULxZlP5shpyHPIt0Zflg5ockrbl3hJkRHphdcbIBcOH5wcBpTiFvJ52SJNmO7D3N9
fQrTCqBxy5TXpd8MJaAXyaraWFOxUHA/nfyDe0ZdVr/VBxjjN5XHGoa4Ml634E4nXJnnQZKG4Gr3
/2sTpDVwT4/7pmMqqUZvhU15pPzy/y2DpLWwj80YnXMiWmbrpQ14p7MELv+y+8lJQhNrIslMyPRG
upFMhezIy7q1eBREHSKMEKwMUURbp9aQSkfVNj0ijcjMUQ8N6C5iDoee6DmOXA+5sRd1KNp7Babz
7pUKHdO1k0VjaPcbF45ufd8A8g+ZE0msZmAmdlymbN13IBnyCy127Oh3Z+Y0AFOwi7IhkUmCRPZh
eEjR03xAHqaY+W0/TDWkr+/aYOPmnDIb6+dNKfNSwZk+KqCxfiL2BJxpc/fWnWmJhu0W2HZ/p8o3
MEcVE4Nm6G2WfB/rBx57PjTDR9YoSDDR7CxcytX78Dxs2DW6jKgxcpLCsmgx2LcbDtbHYRyS1NVL
1dmEUhSVlJ8FbLyyA3OOL6CZkI2vrp8Y3OA9MfSuTTo+8YEy4oWoy/0lpUGYSqDzyldizhbg1y1A
LLFjQdptcjCoAT9MySDbOcVpS+J7UJy/u3s4ADE+Wjvtcw+j/sXnL1H867qXOULqXb+44osPpSXE
7bAdEkF1CC4xeAOHWYaxxjVohGB5y9bC7EYwFQDgid8y0iz87pkMa+aMnoVPF1gYHldMvQIO/DbR
7duaAwnKCQ3gDbfiPuWg4edwHZ1aIVuMyo/x9MDeCXFdZvdZXvwDdLkXBEURBLHmRXXO44IXZOiT
cZNwnvyNDUcbRVqFmX+YN7l6ee7iXlr4RpKNrLMrmYF8q8CxTjOk98GR4+lz1vnNda6J+2RmvXmU
F3S3w7z7cnyQcK1fPuV6m5EHdTNU3DJdVznNroJEgIzFyK3LEOfg8MHJG5NQs17OwUiCmPAVnkFC
R+PS3WuUy3FZHjljcp+NcyHeRUc/LOqQ821ULK8/AFZvARzRuDD7w6wu/V3GS/TzOTgtF54+SPi0
VtXbeZBOTKcxceHUnClMzpvP9OOML2UeXSWyfe+0oAoTiqr8zkcx/3JNUM5Pyeb+BOdBfvI6QAFd
3l18q0rQpgEtBm5P5h93gOokwwpj8YuIHbAvlxSlrzOE1k3WVxjsGwgIWGz6wjFGML5d44lq/5+0
MSx1VUEc8ZSyyt7sBWJ7XX/VyTrSAuH4GP6BTQ5Q8LPK9VgzByLmAqeg6M7Xqx9IPKuo+AzQioM1
0I6UEBX+0lnqOF4ZoXO58UeskTWCtZqhvoghQxDvn6k+XbzHP1AGBgNTO1dhM3pDfBAh2l/+UjWK
bsF69YdsoFF8+hyBAZbIKwKs4OXH5LX+2eQKceXt0bmYKp9PrgDoMKPrsxL+rZb+sDDyvY+WLqqX
yCF4JTP6mwPGmExTHdcM+6RvOD0iGSOmOWyc0sJBFbiXygHfXTIrEVXL3bLTN+xbyV9sYCLu4DBg
gVNdZP+YOjwMBQsfbFgzmUg/18bKk+i9+97dt8dRF0Yufx3iDoiK7xp7Jvsqy99JeiX5QcFNZihC
mL3W+qfolxiY0SxLEoUgYdb4MpsHwxxVRAGkwwd1deobZk481o9WkfrPkktMLEhnsvRvfKYeQWbS
dKoIf4zGSRPj8gNHjnj9bjum26qmi8Nop0JYXzqloNXJNUwSDCGFl6XyByKf18/vIUcRyI4fpToC
fSJCB1GraIAjy9HyoRl8e8gM9pMqyg8AsNWbiXUtIQ5xIlm/eZSzFZ26sW/7rOFiT3cRhZKPQgj2
9Arbd3XkN2mTkeZkqp1V0U1+M7ooVaql5L58/Vs7pi0DwOIkOd68eXGF5I1/d1E5mxUYePEcFWte
/wfhNzta2rqKpdeQpEzrQPMAJAJtx42M+UdP0tzEGUBjsYXY8B7ADWEt1R4zbC85g0awkkfdbqFU
TsRpyBoAOrp/fJrVmEloQPSjYT4gx3vMLpqkRxVzQglxbDYzoHgolN9UBPOY7xr0XgSgsK9883qz
lx6ispV2f5gLJne2ezR8KiN/M3z41i8O6jphuzlAe2s2J1nX2w6o7rQX/YRS3nNkt7Dk8UCsdVCo
XveD/8X3zupbrZPPrmZ8lqRAdBKWaXGAufTbXFRwWr24YXtXkV7EqqBd3KZGafsKfWs2nosVyciH
QSOlDcdrCYD9fQ+M70t1ekt5V13zrymX42RB8JqJWtrSyGyAn7BFTafYpPItzlv+iGS4oEW5ewXZ
mycue5GIoTxzz26AJEgKVJSLJ3Qrv7rFLeMJUpUTtWu7qf0xhvrDQciuvKY613zeTs9FUNIxLf2E
uraN2U9qcqnnN5IPRqbTiQWmg17DY3mwzzCYcgCIja4XQS5Sx6fCTqMGVuHgryDtpx6Yp7OivLuc
OafNRoYjdHtjidC3hkr3EsfgM87TGKo5Gxf9bMWHnWy67pwZ8tT3O2uugc/Vydlww5m/mLu+Q3aD
cs3IrZaikq3tT5wSPp/ytxJiXJ71wJJi/UsXHSu636DbZpUyBRhXvhhOANYVSdZvJLOwo68rIYB/
0072BFwkDJUJ/9pVn6jmGtYk2xBu9MRr2tB4toc1yEP+Y4GEA2uQOOYMtbtLFaQVc/nbByYtORC2
ntK3tnfRhGVCpx4dJn0VSG1wmB9VZLsGwzaLveY4JsxbMosVqf0IX7KkNi6jartce2s81HikVVvA
nxXqhw/6pO9B5640g9EA/aXiu48yEzqWGCiYQzXxvj9SDVdxEZWOEocwCEIrDQKFK9CtVwb7MWTb
vVppQA05SmS4lBNDyOYyE5IGCaFA7Q4arybEMABr+7flUmpadcRrI1n3IoGgownD+lABJU2FBkBY
12mLYHYEMVBW0BDuN8TMF34sKeRed/Hl0VcbL0LOXh9KMnu5FqViayduDY/JqbELxhDr6INsVILb
JxqOtDuEHzzFpHcGT0YC2ZTDr95t3/9Ui4Qb29xwiQAzjOErgJ9nFsi22ZptSV025oBD35W6By8w
65e5A/yw7HToIhrMfzXOsotnqlSEje95FjSeivzKjY0NiP1jv2bjKRDuEAD8SmnWdhRa8mkj1Pr6
V9nwBDxE9SxfkVZ2RkIx6XXJr+gUIHb5TJCDOZNlemnX8G1ebD0OELwFM+58fkKt1W3AnN/q28hR
8ChUnfBz1WxjqpjvZQ6CSuWrdyKFG3mO8FwzPXKrvwRpmV/35+O9b7J17nMt401wZublcod63E1y
Itxfkut9eVB7AJP4gymK0UYeBh3HCZywiTHit7wZjWTk4BNzZukl60/IbBP3YP/JYBFJrrK/5rNK
KXpEV+np70+xcr+hSW77E83NTrvv4ZNB3n4Vjp9DsqLG3jeUJhoi/+BjWdWD14KLOorV2Hcyygm5
qZSfixAGbbsf5Qlyd/VPxWE8orKTp94vDjqN75It5KIz8A0hVWzpHNdaS4TTOl/AYDbOII3jWsar
4Dg4pzyYMHenkMssUfXltshgDeqO0+KeLWF4nKwa6yc2Tw2w/oeWi4eU67rKIMNy6pO/fqhyQ2G0
X6OWg936dtRxI2fBclCKm0cQr7hI87RPmH5vgC6DXL30qipiyzIQZGoPjeM19FYMrjplv1PYY4yF
bsnT/7lj8G3YQ6W3+le25MNBybAoaNbOoXNQHc/e+T6h/O4M1zqio2DVfQrf0L5feMblJPqmeelY
OeiNGRUCyAJGKYwQy/g1pdnOoh2OkAbviWambc+U1kr9uS/pTka48Qa5VT5+dO/flU6U2xALOvns
679Q6jMNtA5GKzMQcpIdBXNmIzroV5+tlqK08Rk/YSuoG4L/AAmLm/2wjtOPCJG98VcqxV4iUDyo
3OixA3+GegBVHsQptNj5YyZUeYuqeCdFq+FooX79Mc4a+utMg64u0zxfvNMj+6ziOuJZMl7nmSRG
88XmfyLVptjt7YJ2GQvMf2gir7nR+U3xdzb+71R3A22g+39ZSJrpooo7Yl1n16i4utYZP01TvOH6
0vNn766LAGNH65sad2NeKb6Tq81MAYzs3wALeBbsoYItnHJ8PdrJxW3iYMKQxIYPDCBfQfezJ6Dv
dwD96ik2A7+1+nvfqEqpi1UlSBdNzvCOcwaR3L6IGGyA4/64PGzxFTAMgGyFu+Q6+ENM8Xf5EXvU
WbAsZHdIQy0dh5DsxfnKMBN6gckA7cV1H8MEjj0Tcq6PyQq0Z1ETMd2amqmlfQsuCpFYRiITQO7J
J2JKIHSthFrTly+N3E4tYfPgGs+F8Tj+L7o4efhhe6xlCzvacb3w9zpgMWCNp2BiNVfFKu/9JFw2
Gz791aHS+kjDQsdskRC1PNwVIAxCxhGpEt56nKe+X50v8jUjuj7oGBSXLbf26O+5TUQW3l1KZzr3
GG6/+w7uDwdj5cVYRsUby6zT06Z4H10xKFbZ9zZxherkgyFFUbZ/V0WDLs/Jv9ssyusOjUQt4Bok
HktitXrb8gsFbogDqgcOsYR8y04dloBz5zl/v24zmr1Ix2sPVnKgJTjQq8nLGe0w4kBt5L5Rmvnq
WKeRR1LRDmTQQ7FjihFz9RFM11HVAz7IUdRb1F0nC29bQaCe/8MdAQN5qzYwdK9DEE6IxhPEnu/O
FWVf8mNx/DpigZ+uGIEdNg6deQBkWGLns+GaTAiuVUNMoMZfgfHUsKyswfBAhRWCMIPr6elcuVey
ztRe2QER9v8CnDSM1GodCheCWCohdO+sgfCZKPsv9HehG0fProoaH5RwLWMJl/v2JgQ/ewOVwbVv
5YPtaf3L1+EBCSPsUGNyFH3SkWCmWlgHofS6Dmn4rFnPqvGRVQhAbZ2u1VxuYNw2rZ1OR+b8g538
MoMt4Td5qnk1CIMLNpdT1FEs8ezHkfR+KhiKLloL1PtVSy3rm2RCcWWJOsUGQ06t3CvKqeeSKz8N
Nc7L4RQ5i3hvUOrgzjbQS4Gzr+w6NutRsa2o1CAf3jSRDSyS/p6VgmnHtCs/hvDlLj1CVzS6HqVU
GhB+k5kKTGY8yq64VIOLtYqDo0FKtDHTE6nWnoTpP7L78TRJL+jd2nvcTZM8iZl6MRTU/S2EZyES
fEEONGnNlEGJXBVEV0OyccST2M+5f4WCRriC1u4hUuYeAYpqpnFmL6L82r4vIzntkGG51wLjS+tc
a+jl6z54HY/D3MO91o6Q4fmYgFg4imtjQIx6XUmY+eDkemoa4FCCMnsq+u1OP4ynq5yqCwQmi1g1
4QOo7a0Bfy+QPeylFt3WtFVV+gpQFXFcizJYW+jqGirbNesc7wBXheANTVKdW2ou0gaqWprFMGrd
ULfbSg7rAg4TP7WtKkxASmjs9QZE8sBBMwHstAaTkRnsSeIxumwdXO5WwBIvdFfonRYJ6ZWcW5Ck
ZbrX/7YPn9OKHv93V3agWmN7cY0jZhKaRth3NSUoQQMPyOcW1SYnkc5aI704EclwhRaSHXMcDaaa
Bnf51OmZRz8USfupp14U/42FlRBa1hBpy7xZDP/S8kp2MgZ6TeT44eWU/sovY/Zq6/+4E0qczgpT
6a0FI799WZt/F5ME0EkpgQoIq2EsaMyW+K6jKtKfUpcU0JSBK+MMKCOPbbxg0lkEsCgKuALoJWcw
ZlPNlL18lAVbZ2fDemVJgRo509q5/TOc+6SLoJvGDo8ToYl4caoflqMZEtaI31JR/ZS1qwbdxxWL
tzGS544cEUdU3XLlpZx0nhZjRIp9wIx/KKfl9DT//pJanA0ijKGcoUiSMWS8hDir9W8YZrPBoZ9B
GP07PNIOtzqmJwbhru2ZBcueClMC9i6YEm+elqj0tObcOhOhapOSdKZpDOkSjpPTCge2YutIhxqB
Zof3korbdZoseSrn3GVnhvIm3m8ocS5Xie/grEB4zXZighPwiwCRLp3xmbkpu55OLGKQAXCEVnsz
rQWcscfvb1K+HLUqgmKuCEsj73SUD7naiaZlbZlDvi32O/IKih87Kkibor1rYOIQ06eZK9JHEJSf
dI8IV0t4TBsPScjlecmVXF7brZ/yUmjwlqs2TPko4Liybb1L6XGWfpP/lizJnjJaQ39CE1UvyRp6
dpvDa85QJ/SibnJ2b2yY+7BE8NDUNnVk9WuBcRAsKq4QaAR5GEaCD8De6B42WvxjmfjDqGfc9jZp
Hva8XTBJ2I6T7jbUy2cnthKv3BICDffwSmhOZJ2vOY6hOKn+kTza6XwiHm4MN2ScIkm8L5iaHjee
TeeK2ydTvuwItmwDKChe++R3RaJ4ntx431843A16GEuy/ND183i+Iq1R2yoEc8we5ZWN/fHa3rqR
2tntzPEDfPTvoV1SyVtQi6FxISUtL/TvtuuZFm5BbvJAlEV/4wGPKmvjeiMOkpzDA2n7GHCDjJ0Y
CqrfREs+lt9mltqfq1VTFvsOi5xlbzyEVyP3gDHZYZ4HvHm8rpbVDH9Gxnzy0bAwTuq3NaY2SGMj
DNt2MOl6KYqUN9oltpNZqUkYYeikfE2aVguS9JVn5/HN8/OuhwYNYTUdxZpLci5p6sFu2u0qxa+N
n+dKthmUVpdGYtTHxfLvx2DR3MfB/5TUAhOftWVABZ53b5kkohvByijCwBpShBSs2FYcLHHn0u0l
raLf3SOPxI4uZIRvzu+0/DtYEjU7V/sqR0mfzkdI+LZRu8H5tmMZHhSaBQcClRK/WQ2tXBQoCGjQ
o5eMo62sZHFaycfLW3gXqqJ9moRsMh5vM5cM1gR+T+4+Xwp7ECxw6rKlCjJAhnSoZaFRWhDjRPes
inoTxNIauaHHmfh8Z+uDH4mGwfJ64XmD5vmSkkLsbB7WVG/QBy3WMGT6iWni900xWAJNeOCTlaIt
8yBo4UFJuN+VPYnSc0GuLpc+NrZ1LyLRdC64eAjxPfKqtNrtdoNnKKQVgXzmgE2ysGLMO55+ErcF
Zzpoos4eOQo9VnmbkStmmefDF+bkMEmjUHfqNnrdmsAtwcfSVl3JaDaGQjub/FhoLBZJe84ZwIeK
skunjlzusW5o53L7z5T4b10kWiMDmuMxb5yrxM45RsHUlTd8ejAkPwCePmZJlXk4859k4oukO6k6
0jvuG+mAW2ch/m4I4QhZ40J1iA/5jNV+P6vhZzQnafqSAjAS4jYsiKhIvmxThnC5ikSmbhHyPtTx
N58U4RSzciQwDX141d9QI5Y9Qk/s/ETtJzVUnPKPhRfYr+RYpfWO5DnCTCywXGC/LD+9mj4KCMr1
zD8RqKL0R1cq1h7MOdV2Sr4zN6Yx2twpT3EPU1ofohlum/rDVUoI/6cixcbIjfTzdqXqEB0DmWhO
M14X+Pb0vZinneggBEFlOkTbOFEOnaHc7l0JtQpqj4YSlmASSsB5D1zG+OZaZfYwxdPaIScXoLHO
DD7sQ0FcvUHOWns9qKbAgcHDdYYLaBnK6fHBGAph39vjmfVPkTBjf5uevs8GFgebE0v3hjBXcxas
yn+W/bD6ddLjn1IJTSfy49lDE//snR1+yJSKjZgjPQ0L6N9Dwo7gTN4o5QeYt3FZ6S3lDUkjogvc
6J+U2x0vpN6ZxvbPc+jdhKAK3kxdXSgee1He58KGqLVluXx1IYKISvxlEI7EepQrnUYDkvOoMh3K
/IIsomp/4C1o6s5xsxwjP1h1pJPcG8SGc69bbCBTS5w4Y3zTpWnU4T0fUbOzyTc76SrW8H160Vni
lvpA8vqBbdWz/NhPiaqBiXL95d5FDZIiWzLmoZrqtzFkwYIsOvNeqGcvUwMWxlMPsBDPZQ6Gxck6
iKjQkOwr3UNQewvRWTQuVzuFjDKpj2tnG3mEA+fU2BrEq7qtZhDYalO5IVd0MKha2emZry7AvI4K
bjhU2s/ghTyHR+JEslpQQHYBs95DQjXVo7db0IE8Nlprwc0uhutskCJznkZ6QhwNVvoA5Lwq6YWu
uhvViUNDrxxDVng3oRX8oiYgsPdf8Xxb/5E3QFdpL5veCLb1GMxG91HivYFi/TTpHDnmowTkKNO3
ORbVx7Gazl2cAqN5kqdkcmww66sxNbe5q5/tY/MqV8SR999P5Ks2BiS+H34XD2AW35i6nzkLgBqz
ymqGp0BOeDQ0SBmbfn7wN2FMuMf465rdCOneMJeNHvibF3vD9HxHMnvsWCMabOCslcarTwJ9gYrO
c32T0RQ8+ZRhpsOpDVfc9LCe5Oht3/hjF76hdLquxZC3r1oPqtGIJphHlq5zDl4uOqS1aRuH7vL6
FBOqryCBaMUFPoHiUyL1oReTFTtIj3KZD0YkOatDBikn6oyIw16cZ0NC98pRJgfGlR3s1s3edXRi
3KJ3DUniJyFET/NvR3pb3b4snUaR3olCCfW5tlFwNgHy7jCFj0XrlTprQcYb3b3NtGFff/jpR1Pg
q/SZHcZS0k0+9C7LQUhQdgFsPbazBgNAK23A8bY71+cq8H5+QA+46aHrrNR3qeYPD/K3j9GI8Bvk
vDVICtaLr+eTWPtAKA1HvMCHJf32gKKzCVZQz6vV49X44GsoLOXYtJiRZ0Xn0+TQf4uzZsxMrUXz
aJS20zFbbIHjaF9bezIsULylmaaBOjYV32/HtAKjYrzMUgInq0KfOyYxYXk6aufJn5aYKLX4KwAv
ZsH4K7aEW3lRMbGK/1X8mgh+vvhdhIH1jvu9s7wRK6mB4deyuwewp8rEgATST7a4R89pb0BKsMlL
b21+0/6CIHK/2XksmJpvbQvhdvC13wqNcgvVdOoixZcJKOnQ0hQYqEcwaT80awV63aLzLuwHBLEt
kOX6kHz42rz6ffJHe/du5vGh8e3cY4mXtM3EU9uq9EHbuUmGERc86acMCXRVxosJC2s/teENMVOG
ZhhtR3NoNu4T54jH1KyFyRHd2dhrXWnluq6KJGFeTq76WnbQQngnD7AvVRaXbaq5QJ1cFJM1pA9l
uiH8szWu4bj93D+0pp1AMciviBASjELwfNji1AxntAIFsVbUiWqCajI1UmIUwj2gPDbNR2eE0pAN
alJHOcl0J/3dzXV/VLfVJURfEhCKvhZNsu7TWAztWqQmcHJ5rKoI2yo1qVfSfDRi0GpBU8TNGvcN
aOXa04oEZG63R8Xa1RD03Zx5GiAnXAMnxrm3Mlixj0sF4UdMnk2YfLR15BBHYyNWJEQQuYPBz6XK
14n2hZXhB3ps9hbUwWjd655VnqqEQhEWsuRTdtUFZoPN3V7DIra3kIkVj0PsFAgoRbfoKYCWUzC9
W+8zWnlEHayEgcOT/54qQ4vWrcEZES3ew9P/gPo8uKEIwvblkUBzYAqRrxsT74UE1QH+xIW2RGfa
hgbgNsHqebwCl/m7jXBQzWSASwtqckfJYZ3a8Ud6V7E+V82a0xG7GcIlT4yc2G3CjIuMPEESrrUM
qYmZnmvxUc/XjZlJwy+eDsOUZ3HIQV9/gG7FzkAl1oO8Obz3iOoqo/4LxFUVM2VhCMNNDeeCjtkT
TFkm4B7CA9tngMOWpH7Fox2/qg7AcZz5HB8Xxu//K3JidsuhjVMSeCA0P7/sum7+Y9I6YNnMF6CN
rtsIVs2zKn+1+2pGm1PG52d5lEJ7VxHs5h7hAjoQp3nVQ/kAWUCvy4nVx/MTiHdHAIoVBLBubjn/
U0i4v5CxQLgxJCPtBC2O3sZKdyS+tYY17tEL09YZpaYxNvjrWX98Hr/KEU7e4rMDK+h/a3Ukm9mc
BsgY0pfoatsYk+sJCyky1EqgYyw7TwXV6DfzDDlfYmOw4mBEVj9/rCHfHTN//DcqD9A+A28hjOeq
2xsmAtS0+4Vu4oIbayrPgjIHWQ2ky2lF/sU4mBiPJVf6XvbnddCtSd13Ts5Byh7EkVgAgYBPkh5H
h/Jwr3SmVJFmGPCHHqavxOOMTJkMB0HRQqZKNGGZtffugC68F24pBsJ8aNnkeYzD11Atzsy3y6BF
fA12q7l1Lo9lTZnc29bmTK3Vq82vZD7UuFm7ZqrB72pWRsBHESlIbcLABw6vuMBvYJzDTSDyIw/0
eihsbgiSc3WJs5JC7UGV7Cz5Q8VQNQp2GgiFB/sMrW3MMvgcN9AEoEFtI2+CIqso9ZfoYZuZORFA
g4U664YGUoA6AJz3h8yyNGNfSzQT+YiIcClvhNoM0PCGYu4QHhopvqd8yF1EafsYu8TO4qc6ZUP+
botgDiJ/7TTif8MVJqJDl40Mp0TNr5Qx5996GevZajdyP41GER5ffKg1PRVz8kEVkUAp/PEP9Rnt
1zOT6L0+2jYs6oPmbPnhAUMtLI5PBObU0YU0fg5aD3vfVG9UG78diSK9g1RG/Uw1F0hO/NTjxh1U
pvUDEqWmtRrzczLkLkmiLlQcEVFpHkQHb8I7QgXAVmFEB68BgKfVZWgboji/XKBgPNoONCLWjdZ/
CfzsSsY9xwdPDwFL6MhdwhIJu8qdzCAe4Ae1STEcFAc1uCs+4JLmCYYLaBVl7r11JIDzi0iWhiVk
pFc9ftS+3WPqkBcQryDPSWJ0jnewkB9n8mAf0BpUk16L165X6U125XI9PWha3OTniIli+mXGF5D9
UZUPiyd4n8kJ3SgqfA51v1yXcuVKhFoxz2ek7LyHVXpKEcNV2Vyj7lD4u0LLCv0mbDblE/lvXw+Q
Uxn6cmSkDJe95V3BhARtedS0pzUaUbBh/tbofhLQsl7odGgummVLdddjpeNDlGIcGHD9irBvjsH2
SLBIVphhMF0Vhn0mgl1hwnSy9KLo7HU8XZ4jRfaEWYxWAmnN4TrpeK/DnSf60Vyd1IRgpTm5ap2S
IB14+s6DumjRbR6i9IJ38Zj/cP9urf9yaBwSZDm9KwF0bz0CmN+j2xJQw/2vucsWbuZkrXvDHOQ4
M2R8J/q5ygC6EgTinQyBXyDg1AC1zCVIGi8GDdlujEhu01CslCZnC848YC2tuh14bWrKEZFNIXJt
mHbkiCPjdNjPxUJq2Ba32yeC84C+LADIS//fQd1+Ahht2m6VzvsO9N8z7xCEkev2rIA4HfuCsbSU
JRzGISjO5z1S0PHTp3gxRl3ycYBY9FXuF0+KiReSEqUNXYByw6JGnAwYbyyv2DTFGOaOJPiJZp3g
owmTwI5aMGcwMs144j9qDaxZZXAYKqZ8R+szFCkd3ygDjHYbxBI3jz5X77l82Y8nZ+GqfLwCy4GQ
z/lvUGsv1v7GHofJB4U/oCytQaTl6P0rKKUCgXjcHGAp2M3ky5eG3CEfxkegr8nD3vZSbeVgrYD3
E1GIISObuozFbr/Kiar4RL6NcArUQJSWTgUHHbTpkYjfQmhVS4rddmDWchuUfld47eQG4ZXbYtAV
otHqtLxdE0BpzhK5mi2o9l8depVB/EKYOEGdTcofzzzl3iVViuTbKzJy/RA1C9oOtIuHvvJ2oR1Y
3D5LkrkvP0BnGD0W+WjFNAq47pS8ollmSnLF4XS+2JU1BvhF0KWVCYt9oJutixIE/sz7/oAY7Fcs
a92A1pcK+K8cGdvHggOqupPTvyv6lelik0RNo3p9knk8A4tc2aLmeHmOfCUqODQ0Tq2GhQywvV6P
G/6oQQeZaF7UXz+BmWDJPF8+VQGK2anq/YYmJIFYlkFEIaw8bUgAd+F0w6NPtYlCijmwTjdtBwQ6
ceoNbAnUtYpsCJ1EM12dAepjqA3p+PHNvIyxLyH2BL5tULdRb+hw5AADuk+zVLWWWJuFv7EalbBF
uEke1oP4xozlAdHDZ2y5th27BvXSu50mlCPSiwO23lA/jGgb83DWoOE7btv1SCcLuypEIlHfuzZf
q4bSXXodRsu/Tt2BzPlQal//e1/M0Fqx7/Tta4TyzvYdr8gSvbMssddxJ5M/P4oJHTRFLW4ZPrey
zjXkrj+ORxQQSZwjSX2IIPr1ZiJF3xWCZLMfSlcKlgn7TApU4rbX4qRrISCgJROfvLYa4zJxzHKF
Cvcj0ihrM0Cwe7wZWcyOGpayiaWvQTZm0y+NDSqbqWuGcbpLV7Qmo/d9CgXLTSuO8eIvSnmrfCIa
c3F/UfTQxwMrxRkB9+5SscFAT/PNkUi9YaLlHHmBXoOv0e7Y+5IgV39inWMhqmlw82RJpj/hsOlD
Slxca2tmibVe1tH+15vh+Q1N+932leJL6wDNr7g1o7EWccLCXvrchNOmkpT+U1wM8xhR722Slidr
Qx+j4N8LwHxWV3hgf/O+BqjQrf2dvteP2/p9nPcyhH+02Z+zW10ryfH1r+nHZRU1JEwXTYANKgS1
ArWnUQ0h9aJbAX/N4gPn4sOGbO2qk5MKtIqqfRYFdCF69LRhwj7hv4zFZ2h8+e4xxw2w+O8qMKWg
JYA3tOYWu7JgK3fIcUADGGywgJDoqOqeHNuGWh5m8CSuOS2IhjjWqwfyOK6Lzz7Sok34cZUMCeCe
We60WKZN/tO25SScWgCu8asZPbNSsIXCfv0cXAE4odP45x0Eb35Jl8sPjs14b3IgnL3OuHhOLnrP
gmPLiu0HcxWZZQMczH4jjBbQbTNHrvd/8Ugu29sSbIJmU/oFn4wEA1TsGPUA3UrrDovKQkcUIk6g
MhuA/X03sKqw7nI9aKadSbz8KIvuOvUyVEqawDFryf5PjNjNzmS32oHseVThcJ3oO2m3lRcNGPm4
ehSrWxBDv0wGjc3hhy5JMbktkFvxrdQnUc13OAWrYSWm2R9j0nuwztQJ2Ob1WgIDrpcxT+TyI5K/
D9th7ObHiBwh2huVUgHxJbamb/wOB4D0IxJZXC0jMBXhV92pL761M+QAUlXlEqv4t+9dZ67zQd9/
qks/VdGynWwW2XOdgIIBoykcXifYhfsRQxjvzZ/vI/yJj5GqLuSUEKm2zm5Sv1sBKFG2c6Ny7OSV
ErGcM6hlfHL5Pk1QMDcoyu+gYpUQMtqWa9FlG6YnUnW0CFYB6Y2P/YiTxrHVRCDq1gE34kIo8v8H
+Sgtf3Y1pq8WXt1eB7ioGEY2auztwni8VbDEMi0JCWU1O7LVznycLbev2d2QscUjL4r4oYajPYKm
WmMe21+0bXZQT1X0Zf8fzQVcaAuPziX7xz4tsORIMe+Eq/oreveHgtLMUaBYWAzQqxuFJaAmaFJ+
zQPHXEttOBXE/kZaDIY2qDKU1FFoU4+AebO/Su71ANj5qAgbXwNaoXwwDg9c+aEJ20Kfum14Zfzi
iYeAMkL8QVzXdBdX5AnbDOCi67If2zTlYQOiUkUlrSGSX4X0FEfjFxEgoTsd98UhZJav+iYReiSZ
teSBzrCGG+dVo1E/cEhTHqMvSsRZyOQShxB5f7ly3SuaToWEHGu65LfntKGdhD44m5YxDRI4Gv0I
4Z+V1N+2krUcZWQa0zIwrFDFPFUVaev2gVLGqi8T4UtrUXUuZnLxHubDMsY3fOkCXpBSl4RLSzdv
YsL/rM1/mbvb8XC00kLU1FuqYY2xq4cqWNMicg5lIjjMHsRsbA47/m7JiHXKsqP3GHlCS8uGha3v
a3TENsmgML0vUd8Gaw29rA+Cu24KFD3Wce1zoyX+Uze/za4SC0Akr6FO5+T8RWUU1S4BOT4mEoJy
+gKHh1meEt+fz6HLmSUJliB4u+pQKeYpI/8H0LxXDtZQdUs9tX6t8ggYoKF+XcRPozvj7mJA3rlP
ZE2xSjtx5FG0hVpqzfB7+ZmJ7nx6mliVROLDKcZ6PR987JJ9nVc4C0/BXU5xQWiJ7b8jmjHSPTA3
+h+Wy1XZmwaWciHxJ/L7rGxSDt8NHz2MrgfE64Qlv4eKHb8fO1HeCcv1f04z88kZbIZ8lQ5RIBDc
hmCHm90CAitadGW+sjJkQItz2B0HUpQCh1Am7TqJ4/wiyMNBYak6VU17IIHC1jeXVIJa4p23vmPU
fgP5d+nGL6ehClDhImelyeBOisJuotJLS4L9r9N9UOKq6jtjVSLPPaHFnxZVh2a56H0uDj+2mkcR
xSycOAuPkvkTytr9lac+rF6hq+jTdEztT+Pq/ZZdFxFHO6QimsAVw+YBVFDUYFnh2k5sbApvI9+g
Kc7JUqrfHh37gRY8xEjhtUnQ2ywstYQRhdLjxJ3GuAmktOLZwetSecHd7ti/R6w31kUplmgVEF4g
LP9mFxTQ5eSU6TGSC3ut5w3AQnTnTmbV5QAcTPb0YYAWw1rrX0zKWCMTUrbDT/97BfzKs1b8NMiT
fXM6pzQt8oJthnCULHkojXSa+mV5FbBBRFFXI6q9Vm0OkcJ/EmRH8RpprEy4rcXmCnOJ/4k53+lQ
SkXzctkTHCqT4+A3uXxIaGsSt3CHDdyptdRdXXwO/iet6q2LHG6iAAZXL4PXQAFoHscghwxtCB/z
cWkFuzC5HwonxLOKEcwYdSfH7li7wJ2FZYxDA0g5djvaPajWxVIV4wtNKDB7vLJXnHXXdgNEem9q
wnI8N6txnOUDYPChMaBH6yl2F8YxBMR2tKrVm6QQxYGu08Y5xAjiGDlYPqcin81SLmmxo6yJIhj8
n5IkjWz7erhvdJCcD78VG+tVbTzyP+r+jOqt4VilZ6RTUNmUmavLb6GX000xK9lY1hmwdNelIxPr
mzSCVA0qrf8niYtgtXdFatiC5LYj4hg5etDnf5QmFkw9eOpa6roDedKkSlilLSO60urGkW7KpX7A
59eIjttxWMfeiEissNFIaOxlr/aF10gBdHuJmnsuDY38rFibBqYhhcIBSq/vR0AglANvDBR3yhSF
SDr7mciN50Q71BHcSnT73fYbwdj2WMRE//2C9/sqFwycYmkFTYtTHzrROUDgZFOvpLeoAssRG7nK
njbauzYZ7voHikhb5x5PTQL47G2wgMyUinFK6ZiQToz6LfJg/30rOUgIMd6Ig0pVMZB1KaUuvMj5
EjkS7RumTEnGkeqTyKMIGbsofTsErp1DEuJD6eYvUHfWxXaKafW0WjaU9uGRAQXsmdVcnW9CQO+u
6qApz7r7KBU9lJJ33p+1ipcf6oswt1M/rQqbPTJ/bFELLYbVF4NEeKTVab6XEYSCjMZDpMC1McrB
e096/3ZO4a3GLokZTS06PaRd7fPTInQa4kqJkMMNTy2qciSS3LNGAZS+N1fyfWkb40jwHZwYwH+7
u1ffBi30Z8VbzX2XqDAeukKCgTEMANf6aqP1lcXuESNCE/V2DYhWwKkBBAgMe8Nrycraugc8Byx8
6Jg7ZVXFNbELi3PiqCo/pz7xmIqkY12tgAHJdj06gawR52GqS1axDKrowDNR3yQOGUc4zEJanMRv
AK3jR1M9bfRVDkGs0vrj2x6+x+EnGxH0DwMYTsVW6uAXFtYudJptyq2EgV084cmYo3Y4xEUMnntW
N+RdS9JXjpQUVZFPiVRkG+TTcSMFug6c6XhhT8fgKD3Fyocr76eJ/VQgC5aX4kgjKQVK4qaVvXj+
g8Zp0YHSiUk23Yto3s6fYOsgoMI7+dHqXZO5KUPxjbu96pyjwTHWRY99bHSAsxQbljQiuXqmuUxk
TztfldObLKKjLOfuWT3DCrEqWyBzz/lgcWUaX95QBa6VfwycgkHCks5qY0URb9iujbABvU8ZzcU/
K+LfvdSLnFQ8xcg7eZiC637lLSesmpqGywolR6/AEjHi3rIoKOcDfOkqV233RiGy90aob8jWsQW5
a7f4h9HTp5JaJpfKWf6Yxa5j7G6yD7Bj1GXDNkCAuMpwns2ZEsgml7TZlIIQEVtJk0oRoptroEXd
pseuQG6AsKY4QVWI7MkYPoQwwa6zOlcG/4FFkhhymNG/fgcPyXqI90rw0THjc4C4rArfy7L8vSY3
kFi54J7FpPCnXoG18vPXWpnI0T1hmLyXqiFifhrlhf18yZd/iz/1q+7WBcwh3DwvLUQqNP00ElgV
e9pMhyPTGaxvvtCGpp/s8vbNEtehCCW8So5Aw6VtCm75bZ95UZwMiQt9towf7aNK29dQ42IIZZL7
lHlaOFRKyve6+nj4swsKD2vPaEW9SNjIhjBENbzUftIbT1e0DB10ilUme0Puz53RhgZ0QV/QNbf/
YhEIQiD+1GDtbq44TfIgjVrF/0HrxNcCCvdaogoCiyxW0hEyeKNk/oespGs3uIB1FQtQ36go6o30
3atQUxe43ZhGzmVYM4g1GAElLD/TYjK9gP8S/AW7OeYRgq6Y/X59JDu3utq579SPdzl5z97Ue7mR
6UmvH7pfbIzSpIzPFnsoZTa/QltoTE0O7FA2wgmDVUJ7ex3yXyD5sBjI1nPYFU/O/stgGPCsVcCm
5IQ7vNOUFjnsGvMR48OCTblb+54lq/XCqOONIWhkyl2+0NBHIHElD5rHk1r1rWYYFn1SMYedYeK0
BOwAmTXWeY5Uzum25tYV70/55Nvu1TcDfjS+mtKu6igxuycxXRXHf5+BDRt58DIF9M76NSJKz4Ze
fSPEPxRpGj/LRvF1SPZgHJEb5HUex6xpNh6JKzByM1/EmBSMcQWZ7isNkSlcmkD5qoqDRcpISbLX
X0fwsTMmmVw9N80Nx0wfwUp9oocL3t0UK0HmRsl1gFerfti4RCMSZj6WZj3rybJpMUobr7ds7667
Xwt5Fzmpk9UMW87xitnXI7DUkGheKHJplzppVEAgXAUrqRvXeWwAVUjIRVYMVD6UrvqEx8DruKOQ
nfCYrlSFMww//PQ5YvrlsBgBW3WYzTgXHcglnapXM0QDauaemCO89+u4JkG+kMnTmZgAnMYzcjIa
A3Ugh0y3xz2ZU03Dt2v+VmioKxbsMBo7o5NNdciOOMLYirDqWQCRbpwv/+aHm1N4wJtTrLmHrQ0q
GQMOvjpUyUCNvH8xbFNk/ONgCj8ALqAv6CVM/EiGNlte3u18Av9FGn7Spc0l3bNkzmCNSrkYGh6E
56OAsfuoqcuAvYVEmqbAyJ7MlmQsOsvnPuLODnaKIZWNMQHW4ZRFGGNvknWuKEYoLH3sZBT8omow
ehFqtI8g8Iotg2ps8bzZYihx0RCjG1+d0leOuwSWXNROyRyF2iUuKDlVB9kS+lSLmwkWtG0Y5oiT
Oj2iFi1phjNJPLwdRj7q2NemXk51LEmfBJJLmxY4VE1bct10L7zgOWpb5kEzf5CAoyMSvyB5ccXy
ugZGTDngQYrXsv8eBVIUa2gzmh73pgOYyN+NrGwmVTQuFHpo3Xkiw9Kzfnmphnp6iV8unB+lYBSD
0q2k1G6CZVN0qhLq7KSfsNmz1keDRKSfJsd7Ju2dGnshPx4Mnqnzi3a2qvUerSHY55GrNkLGRU8e
aGQ/vOqPOIyRMadQg5zn4/4zW+9iduIRO6jwApTHPIJc78fZ1hyOIXM9fVTsZqVw6gD9BCcq3D9L
zt0yQ/J3+j+IItzvS5AgfAG+Xb6K/fQDzyG6ppSNbDFlHo2VS7k3O1J73xQZTlpO2K+EP1SUqqpZ
XBA++RSQEn6uDl/uiwtB9PZBubBKj5DHFnvN/y0C3pnwlkharCekNlkloYcgevkv6fBAIThQY7t7
VG1uGRFgALxGaAq1KyOQ6XAh2RVEQtpy+JhL87dGPYJXsZY1S8vq3btgD/UfaRy+X3nTZ7aO/7lO
vDnrRIGmonV5x6Vklloy36K8AWZI4X0jEvWOiq3t68ejdqBovyKir9GHuQOulrL2HScLWZX30Gkc
+JN//wFMF/AndkiircTwQw0L71pfWcwCVLxxo+mwEgtH322fnF18mUlNwQckBIlQS8agh2LRQ/H/
k4sjMlZ0AyrQFPQpjHXSDvLBFR10wA3rQ8+QBZtNDvzyWbTubvI1MGPnkCq+3bzK/Q7QBGlxcwGh
dbqJFQwqTeqdLQrbipuaa8WU4opmRrk2Cz3KQUlpx4zF7cBHih73j87iu5Oobv0xe6ABGgcN4Plt
WB+95I3sL80SRO4pW2iFekxfMOqpNoq9aQMBtApNXY3HWC1U6W1V4YKu8OzWXORYThgFNF3tmvYp
VOwVg47Kq8PGohJ8FEGVceuiHZ89fJMXi99uIgOaKmN367yeA9fJcbElnu90lrx2i8sPZmwUJm6p
2jnASOHsvJbM60Am1Q1qqgIzqd6T0iWzn206fddNo1b2wLWmBemXy4BbSM27MJ4yUofdBReIhUAQ
8ef8XphRdEwBN1EEq6lGrOby3FglJln0e2+Uej3f6FbpHjHYkOhMPnWEg2oD7IARZvw80Gc8boyW
38bQ36gVIn5WjWdfaq1rIOtrvRZsAUrm4oOK2dlH/NB34zuDgR7uXrq3VtZvV63gM+fm7/TrEye0
xpYAxokAFJyzzntpf4dAkYhJ0rzZxQAq3sM8lYSorvIxAc2aZBGnCEdhMMflcqJdzgRQVZFkLOuL
u9NYUZKCuab91WLl+d5Q/x7a/6q+FW6Yva/GQUfZZqfZfCYEg3XjSjxxhNPetKmM70PSbtGOsaDb
p6hrt5Uf6gwmPhdbjBo2MIAMV3dTsSWaxfRvcFJvU88kgWbOGWSlUSqpW1+cx6vFffIB+Ij23s9i
gYy2AeqsoUHGfUQEldjU9M+N83Qx1EiLhGqIyfejAv6Rqs0XcvCYeIZkHF+U6FyS/QrTgAxUZRkk
e3p9e7oJCf9NPWnXUW1y45/yjS/s8xvLS+b+BRCmGODck0uBksXkElkYXRbv0zO9IuZ/yr+ZFPkh
Fevai28KLjc2yaTMtthSKl/V1jG5XQLzhiUZ77VbYhmuvCDau5zgc40WY67KXzl0QxMJ4QIoRPZf
zy/brdCvYXR35I3XzCSLQMfgQNQFG+c6ha3useb1QnzUuJzyoxT1ehoxmDnaJNtd/Hi23npLaHQM
aN54BCNcH9+vJO/frpWXIJa3nGHw6B8sKlA7AH2gJR8QkeZ8JjkcaIfehqV1Yob6HwOJCwtBpqBX
0Ei3X9qkvNde9wO7yPApB09BmlTFudrpuP7RDRdsug37IaJGJUXH5furdfOB0gwkf81M43dd8tVB
QxRfqyNb2iL4reTQNI2estQgU/5ZL/MI48X8EHyjIpYtDPF+KOkJdSO+LA794UDy4dRcbfWVw8px
te1iLr5WbpG0xaBKWNE/UiEnSKzgWSiLq3sw+sic7zZBvkZxoDwBI8OtV/iZJNwKjK1ZpgSQ09JJ
3uFgnQuBCFef2KsfXkDt6ysZofhehhShFnrUc4v6vM5l6zTOe/CSgyKJDkl9ctm2T7NO/b4va6Ab
4Vb2hoA7WvjsbnlhwDwtWXmXx3avawpdPtiFAtXYBW+RvYnQgHlHJpzYsRjyLcv/kRT46bwuZ5mL
6ENTaxAK32u40ALEKFy0aRuDkKe6/XurWEaicwvJLDM4eZc/JCIGSN5B7o7mlS/Y2Qf4gse1m0RM
lQLciGWF701MfweE+i8iZJ3te0M/gTqIkY7Rocok598xwLacKM73J+/kzeMuhyFqFrxvU1Zdp7Qi
r11TITBDoTuB23pB/LvK1y+uwlqy0Dy1MS3OmjGog7FHxdQzlvOhLiojkRFi8pTnz7RaONObcXov
/z4MJRfR21RVOd1tH16H5XNWBXOGzeYRUUucosDvtj2b8rF9Hhbdl+UgYQw/X+cG2aIp1zafsCcV
1MiH996HFmi4Al1u9Ix4WL+E6lO1dj8ck6JbISrkjzDA9lLnk0ELvLO+3P8y+ZGB2++5J8NnQCYb
fvD9nnlWqoFCZEMK8uUajmi4b2uFHii4Sibsc87TaHlj/5YrHB+G1v4nZZNkMmfji4oXXRV8nSi9
aaO02apdFr9x39JBtFxQArgxtVjMLmmQtMgMxGhxGhb0PdYyRBH98dlakSTyavshd+XWa9ykT9V8
jgVgAmQhYMbUmm7B5MbWWwLleR+LvHzLvyDY2jgIh13Yjn2B2F2l19OswczD0oqD4i8C49eJE7e+
2BF5gWdnwDVVjXDPVJLoTl7lFiz3EZwk01vFOcfquOTr8/Ze8UjMsBTV3GOFlrF/oBvs3n6563CO
gg75ylwmZ1T+Z07vMZ27Ieu8c2M/KUYTVVY4WlBeLICOHbWvs1szJCt7/RCgs+oZlAzbhnYsHmMf
WrFpyGpEOd2+VEr5XfFNvYH+ySk51ZVeI+DsTR4lU2Mg4YSX78q2vGWkVuHJocxyDPuAxhFeexIm
RwaPAoGkIFNkWEGlHihp8yFGYql8b3YhKRBT4pYF45bc+rGCqM1WcE4BYHPoatSHvwayIZ/zoM9E
S4C5RY16vi98wNQ18Ys4AJZSUXFgIo5AvdqTZmvhIVo4husRRHfaXXjxqfJ4VPohVgxN5Uv6Oj0r
uOFdkzcHDEqvvChE5Iyjaf9ovlJPJT+IanMMRzhMBJjQTmAqIx6oQuNlY8kLKkk2/5aKNrbKpCcK
Bx2ooAAYeO8HTxQH+x6fbY5fvZdnxfKY+4OxX/bduHVc4blzRHg1zWRFFa/wt1UM5lF3mSTzu1Nk
dsdNdqI/kWaYCgoJV4P9Cqth79q6L0kMhPQjK0aox+XuMdQO9bLpc5goS34FJ++DurT/IY4c+qlZ
CErT8EhFDCpANUcjnJAFRcAkNtFUFdXrKIYFjIUtTq1dR8zF5b8FeC+KjJB9ZDmzz1S0RvwJqP/W
2sZJ1uwwJwWL41CJNlvib/rIflKFZ9gcUhs2Q33LDyf418WwJQ3lqI8W+oWlIgljoh1IVNY+rrcK
RBFHHB0GcFLl4wf6EwNnwEwfdlRSFzA6yDt4ZV6TgreNZJRMA6TrInn2Z0t/35SVeWnVrOSGCjH/
B9tHtS8/nEUsh0Y44SpgahhXJkiIdOjTXdGH9yxWxUkeD7thvCtRAU/r7Dfd9kC7SXbst4gfQVKv
HECXMkLIaOrii6xbPbMD0E8CNZNEzUZETGa/NVv7qIDYPI471uSOf622ZdwJZPqa21c+lqbWST32
vloZ3pKcpl/GW2q3REH/QJ4DSBzPYCxR6R8+t+i/4Nv8GUjQ6DGsEPavcsoLY1MwS4tPw7yy7bAs
pFlHnKh442HH2xzFIwljHaZs180ZaTDc4O+fYG7FNutMPOATwb6xSPHH7/2EOKWF4n47xPMHV3TW
BG2TW/mBuWzOM3wNnz9cqFFcs9osuZdLAqB1GrlZt+yB1PMc6AIIhyeSqm/gqlWOrGHFUy82F7K0
/DNBruTjsIS8bbhduMOUP+1nxgtgCy4JFi7TqaIA4fR986+/dlLOfMmIhx4xUGfXN1iw2k+/8SLI
vLLG8NNmfCROkM02vuoVOpzEvbiC3jbB9GrDMxfSQ1TwRE9+mZEEKNZd42oEemYUZgX5wZLCphtP
bW0l2FzwVgOS5oO7gteIvl2CLVm+zAWhga6zRhyAhJDfZ1yFSapj1tN4RFJ04+cFaKKFQufIxfB+
wHXE5QXB35UmgSgO1R0r/i/X7/uCT8gxDUrws1daT9LssCxlLSucomcbFBb+41fsGUQh3O/HqQAB
w+hIktafKUFfEsJ6ZaQXQxe9gom+qXMrfoPFyU6tDT09kLkllR3uoHQEFlZ+6yxVNJtl2dNn0XUN
Hqh9n01PcPUe0TqTkfGMX6qVAmOxL6gYB1izP50SyY77kJJRzHTMLaO2L63HLy1OvPE8GtZpF325
bEZkQQ6DszSNuhSRYvDAcvixcVHm/jPDcOf3JqN920N7InbiW4vJyqfPQbqahNm1VFbO4VT22uB6
evySXRU+mej7M/V98HKto+mFm3wYuNo1fSSy+xta29/bIuCuaiCfcVbCFQkX/V+GmMJh80nyncMJ
g6IIT5W9U8dVK8VUFn3eYnZTHqs9Awp6zCp9HuJ+2MIkZZ5sIgAvcqK9wszwAnHnMknJmmIKJyA6
rPxyIlxG0ziDglaqrSt9ICI25BCDbcHTDHV3qVKgLYFfZYsMAA3EaRWSXZeOfEmB12aWaJ3K1ZA1
WurqI64JjdFtqODmDoZc/GcrNiz/EwAfKSDpZ6xzdQaXEMqcn4239A7aiikBBIu/Y1KNnacTuw+u
t4D5blglloY4onBnG2VDxXLwB7FQC2SONIRk3QSx4wwcVXSb4ZCHTYrcgyfJN5GSwGigRDJLErtJ
vova0JzoECUabhqrNxyBN1o+yoFFyxplWv76nQp5T1U2jBsdvXfVDT/jGeCWtckmD7gItFtnn1OO
xfhKA1nwH2BDg6wQ6uCHUpL4E5fQMCt6mJnZhLew7Y8TocMYll+99yZpyBY1B2f2GUMtwQJhhc9C
6FouDsOnmIfeeyFhywilhiJJPz9BmRjIQ8qEa2ldPLvbNeqpEKf7onpTCs68BWDomHQr1i/lSoTC
HiyRsR1zKdrZQw2VWoS6jHhpwzzcqSuCbxBJz07lz8v7+wwWhEkaJlC1FqgvqtD4P2j1Hqz+wfrt
cW0geuT1QyA22FodYd+iou7rw6n9nEuHlclaF1y86lJA/nbCnO7RMfWO45+hqnEVLWeikfupLvsq
M2KzJEIReOgTJTVCmIJ5bttpskl8tHCvBMlCOFUfIhmB7vCJCUoBcrHEe4Q+LBBvjeR4AUnva0rO
jWzc9bGbICQJB2bPGbQStrw+R0m2un4Td2ZDSatezLalSsgrbSJUcqoOTMYPjB9nleKHrahxzCgj
D3h/kl/B7ThIjz790L0lsRLgIU4b5UO6X/aU6HOhdUA/rVfvZtCLOl1ldR2mO0wga0Rz3QkiTdF3
3cGKA7wApSfvCatNExdwniU+HMPl7uVFuJSypIuNGrLrw1F3UUfQrxEO/2YqdENeXPsvMuUN/QiD
ZBF7nk0JU+hp5RN+AoWhKXI+h3v8G7/Vi0c6gujgTc8Dr9N8De3v+MyXdzs+crEAIEHtFT9Ze/tY
4GHHKoYbNQMmiQMXyjseXsLoN2tlBDqNwL+YSD4ome5CTo1Z6xVZ7mydycRmqJCWe9LbGREbMckR
VYpsSLyLMjR31enAK2xcvM8t/XtE9RdEYAQuS+ftFjhwgfmFEHmnmYzkvcxbFMI3LP7x006+cIVl
+rODV4RF0VMY7ibfrjudr3T2f1UH2i+uG7ku5NQPTfoqijL3mLVZzDhUjYvR/6JhJxAgsGl/6tK0
LWYjBMY6xYggKs6AyXpx5WIsHi1eRV6RHZxEzjwEtU5C29Z9SBkqT/6eW5hgmq/PP90ASUcYRPj2
wNN2a/M7oGZwQrKrq8d9rrzpy71n6i2+wiI24YdX68ycu166udTHgUXNdWm9bekOyWRf7RP2l1gq
ZabzVfe/TC4qpSORP9f9Q0ILcO5rysH48g66NMvT/aeifWz2x9xn1AN3cSvhb8nUrTJIlTSoCVS+
TkEfu3vyKmWb78TcUrTGdifVY5CUe0a2BZ9yTpBwk3s0YWx7NifgRfTsb+1XNqsm/Fctpgb/yYKE
hrbsezFdOAdwB2vRs+BzADGzhzOLExwD9UgiZFjvZ3IaSu8MYda9z2MUxhT+YbbMfm7iwnGVxpaD
857WQEj/QwExIduYL6URDG+QwaYqiflEim11r14RIFLTlt/qfPTgKGSLcEVRAYhTlWFE4+x1CdmQ
5crIz1aIEQD25IxF2wTGN9DtT6gRTx43I0W0kFeNWvDLs9mzWcp3P5va60I8gLEN/0ylHaFvAfxj
8U9gK1a1N85+gjLIsqDpLEntouig76TJ3G2jxiIv1fAL94BKcifUohOAUF05zVooi4q84rDPrnkM
kbbXXkPsE8wEt9pqRmNp/N06Az4BqLLj/6v4bGe2lwTpFiKFNkmtqt/2t8wlSt6o4JBPGcmGu8YH
xDkbqCK35o6rQu8NRCb/vDE6jaPrKO4sPur2N7XuXIANLdYNW3oe5vtPhTFctmwPI6ByMHXts7vY
BtAUNleMzZg6lKhGyZUJAO9ejJqz+LxSfH8N6duZt6G/VjFIpi6u13AjF1NR0PWpIxPRyfuMfdne
EWkvuRzY37h/kz55l9ZdUk77qjDs3CIWZQkWiPhggs+V3smY8vcwGBmGezVHEQxqnQ2k/ALfaO8f
wE84soW5sVTxOuukbUzYOILEP5NN5H/CyI7wtx6/eANAmAzeBGqrbuAOlov4ezzITn5V245Z6T+s
t23x9SWGbx/Qqd/4u7avlf+hQFxWICTGlTILH53A2Iu+pVJMgNbvdjMEMB6aN9aAZWMAWwNjzHpQ
UdwzsnNBeW3JzjcYwRN/+HrVXI3nhWgu6M87WM+SwTzOREFieWcQavDPaWFaXcNxn+hc7KYi3esw
rQPISxVsFl7L/6Q7shmOhebj+KUUOLdOemm8YZ+KN/W+tHIsAnJGPihutCkjdac8ua/ci2pC5xnp
jUjhGCh8exfeHhw6KkbFdjD6j6vrx6gjqKvKNZH/PMZyRPq27fA8jFEF027cZnMQ4NJMGB0KJohX
kZBi5sXI/QPSryQ4GfEhCJZeiOFQh1r75Rtb9aYoN4tVt0dBfeA+KvTiJH5EeNkCwW0aA8+9GDRZ
APfbtAoYjNmqBpKIOx0zxNh1hRU7yIdI9C+pGk2ZmYdaRStijut4WZGjp5LlCZB3BlREJMdEGaa6
5cdfYVV+hRhynuaoyrVckZphCJyBQSbE7siGa6phpY49MrgKOXtrpkMP5biCpAbDW07c6T7DahvH
iW0GJTZWdDZkKcBJeCmTBF6Tm+9HCw2jhWGAxUHqaydDn4kkKmgXzOb9pm1xpe6uWUauNXwn1a/5
lnKZ1rOzyTTEFtETs5UzG50C5cn+uhF708gIHNIVLwaqjcLD6uVK4fYolvl5Zkstx5C7QLOoLe2d
SQe1gQ0vmN/qeHbLmG3n4lyAMg0Tp6lKXfxJXAQfY6hlNlK1rwPIxO+d+NVVHrck9uTz2wBG5X0W
zOvHiY2uDBK3ZZdhgHWpaygyXyMW8L71W0m+BiHyBu1x05stMVl6uuk5TdqqdXtn4xAuCyUIvV/r
GT60Q7jRrvvMbAw2ritnGFxLyNXx04ciw/nI8e7e/V04qznY6N03l18SQS2R8DNdHeRH0hRcgoSG
y0KHkakq7mRyowmtlHP+5yEqv/cRyXNPv38FMUM98IjQb1tmytPkbL+mHzHH2QkHEBK62Klyo7qS
Ea49GM3dSS03VIZ9o6KBXY0PNf/QmB/PTvfJpqTRXovYQpbaWkwkqbLctY6oua1yYO6bK5CIpkqx
H/t3ERD3nuV8okn76184NlxRAEYqBN6wxFtZ5UljfUPoGLiI8yeAf9l0Y0q9Hfu21jws/yCF1iwI
TQv6jSe0Rq1qxK5f/FAFLxO1qVwctbZSwhTFIrbPW7PObxsROXpnfFg5K/jnxur6AMUwike0TFOn
waFaHgc2ZyT+SPDQh3AjggobvcU9S89wLtpX9f7ycTYZDV6u36e0zxGYk6eIhltaJ3UXvkWRmXtM
IWNKZeW3g/z9Rvzji2ODBrTaWyduRtgFy2gNVST65JGY6PDkD+W5Gri/H9jLDWjmAizpUOA0v68J
hehbYaX4uL9Ab4v+GVJeBsYN6mPsdVVcnIedqQCjc2VBXplHVR+cbj8odSNVGbTa9p7Su45u/3hG
2M3GOqelPElk/owZ8/IyqpVz09yFqzYH2v/YMJKrANjt9x9exZhCaIL3otwAtuHGex/4Wx7yg0iq
b1HtHAATFzM9veOlcUz/i3mvxT7OmaoRM9IBgoYt+8hw4LjlCzWiwLSkVlgMGZAqZAQb4/15qZbZ
hyIjzYEcZ+bAbmmXiPahb/IUdV8RIqT1DB2tnr9nS0VVJn2K1nec9NN+pF5Exc58M8FNsJJSCdR9
0wCGoBXuup+2hht/0PS1h4SX65Dx6x1+fbeoKGJOjJcL/HsepdcC0+l7jIRgvKumpVQtVE10ogK0
lpKAlRzZVBJ1dadY3CnEhAtgtZNnZ2X0biAT7zHsShlwRy6bVWXTJcWWl3ITB2Y+mjUw/IuaLR7O
HM3HD3OK793pm4ui0hCTRAUdBf476h2HT84kdzsUgFp7D4tfZ1TuHmWaVXr9P1ZRRlPpmUPF/dg7
YJqgdnE5v0+UZuRB9qLUPmRByztuLY2PiYCa/bbkFKcBQZS7NWFXnCsyXMbBIMasqpb+6gtDZo+6
co1PARXvFr1ODRpGESPip399qdU3k8XyODOb0sB+7/1AJogP4wTlGjEYg8i6ySjWpInTmrHtxZGy
c0D/Z9lvPenoiU/NUozxE5TovIl/QUgVUXhR/qfvKy34IkKPz96UnmJ/slYwXSeN2mc5UXGpKhJB
R+WQKyiAVkYNlzjKDHBDkd0sEAdsdeY3LCmaS2Gy3pVVkhSvXNY01GVvv4xKlBzni/bgonjeUnFt
DTIku+16OXOHJBrGCdVFRzm5GOzohaSHv2WUfX+TAkWCs+MexLsxX/hCeDbmJVTpbTrxlmrv5M3I
TAuz24vrPLUNBXx3qI4cseqDv7sd6pL5zgmjw6pdd9zMRGeZb/O0L4g04moGteb6rC4QW1fEffFQ
GuocwZDTnaKwWJtbvslZjdvNyA4wbRXYlaXsDYBuXdih3chLKy5NLcbhENT6GQvoiCwcY7R13/zm
dmMUtrCCKVIOkkFECeyRm/V/4z7ZqiZXtA8hddpSNc9D0UBim4msnUmgjovU3R4uLTD6vosnjucW
92dfjRFLNnn2pB/U41JL6ccWcNyyMYmWPseJT8Bq76X0nx1MaGlcEesHjEQRaHtb3Ha9gG57ylXE
+JKiTrGnU53PXD/YYohKTLf9TXQaiIQgqKbvhNUKy4/cXe6bIRvttTdA3K7S8jL+zzDq55vI0KDp
lf5qtbgM7/1i0ZLCb/ay14PnlrFvL54EzLdGqko7kh5D8EgTMD21sVpjHltlSskNysae53aEllg0
15M12c7MY7XWfY1AqoFuhWBEst347xyiBu39hpxulUY0TjDdBnBZAgkC2W3Z1z9Yfjm//qhxXxnH
iprE7WOjaEJgSKMTMzq+SZqf4IXRYEscynwanrb7LZwpbTLI3b9yp2rFjb07UmY8W5rrR08G1UjG
yh9RDsK19KjZVrejFLjGuP2yT2E6uXBWoiPCpuCMuQsg9JjbVxSVFuISoFrpd6SeeTbM8gFCDLXJ
ne17oFeVTkBy8TgrKfzoWtPdG3FViRnn35oGsA8yd6C5pxCcr+VGvXaH+0TGOMR8LrQSJz+Zo1qt
BqyPeC+FE5hmAnxmUWPyV9G/OXdOMqmT7bfbpevGZU7d0eBuRelqHckqEw/qwIeAs8yrI9sHbHOq
EBWzjELqeOBVeBn0dAz0dGKqpw4Z1ptvf2UFekiUwv1Qe9JfstHmlONqVdbukhs+zYsbdRBwt1OC
Q71s0PrBvFnutUSatEfkw1tAn+7+UO5cOFFYKP/nNpRjzlmb3cCQfw5REgZiW6TfPHqKj6b4NWgy
VKkChnK5cajAHTaHGqKl6IO+jfXJbmqjUR0ypVFJxNgwDMLycMTEcTVVSzfLpx4X/G5jaqzIqrLK
UtSZM+p8ILX4ByVFBHFwJ74KWJKWAi5jDhDJKuYhduXTFCvBSogKHZUk49nJoqC17J62sPwkRga9
8bS6rYNaBVRRS7CoV5bx10U2RT93k3v4B/1pIY/z0dyzZ0wsCpnBeDtMad8tw1gTb0I7fdT1/5vN
BV/fjj5yZ+jMg7s45RfWjySeNN90OSeKvuiHm43u4CM7q/9CIsI68wU8eWgGXBrkOVox+Y7Pra13
epLrHfj8ThlT9Kg3Scq9/dv08IxwI/XtCIU0Tf+eubgsrgmSdLJXKujHFU4lz3TmtxhAv/aID2H1
EpbwDkLesKO/xa04VNdZK1blR338DsHFirUzyC8JTAVfEKEDuEa1p3ULfqKbDmj/OfgSfG7V9DSC
Oa2XFS/md+i5mSQZRJDjMzMMKND/fG3rjmHK9ZJ+A63PbMcDoMT2n+Tfrt1mVw6m5NR06etdnhuW
skve1M8gvYV4oHEjhyGQcnms6fLi/06/Dyj37nQQ8TsFAO4N5bQgckj9BXAdSiXFFAc5J25vvm3e
uYDFevXcvjhsV97Y1y7ljEvIOvGOn+H/6WYwyjLaBWNAorKqzRwxCjO6/55csUPXHtUg7XFhQXbA
73E3BJQgYjoe0UZkUPJDiyBP6hckvtH1sK8Qdoop4XwEMoLfgVMw+WoglQIq9yfydrBW3+Y04GpN
0VAFCiLadYExhqamwcQEwXV6d0g116mfCrccMII94vEIqQx2GkcgsbkgL3ndGMLR17RmXbhZzzzk
5yxv4wDFS9UR3lq7LEAHu7WytJgW08WARuZb9sHrXtPLvTq6Zpp94tImp2SNCG4lycISmH4H4iKv
rPgEYdxuKuW5Dkf7OINoMR2BBg6+CU1AlD1pluklOoiOuvXo0NuBoChnrRTcd/8wjqAJKGL1J5A6
yA3rK3T0mZQNmU9/Qc/ZNHn9gho6705PPb0dtrE2Dtvc0JFBFr3VgZlOrFXEDC5oI7dZL1EJoOK7
rRK62o8jUWfQF+N5np3RU95Khnif6CgGPM5L0DRZQRld+0G2rE1aETqFClrRH2TpG7B1HnYdOyiE
1tJAQqVntNwqrZgvzRPsLsF7WRZAsxiqbccgpiP4TxwzloXgaxY5hBTZkbXszzI8Vc8TSDCLkHDf
m1J5JXbdFvpbBPCYqwMWhw7R5U3fZdbTNyT63KCN9QT6aOxo9gAgSKW9lO22/jJVD7Rcwxu70b5u
MrYkIw3FjhJxYYvJztzkK6W5j3p077uAOiDmEgHp90G38lzMzbGt8EX+aTd9imnStLAXJbFGSpEy
jicoRX/REZ3JN8iNALfsJ7OAvDV98365EfklCo/85ORQQiYKYHKXsJceHMiavk+9LEVrWYmB6uQQ
YbR8uCgq62YpeJENal7tr5SxI2s8rysyK+QzD1YosJA/tt4VrYr3gDMQSnUNnSxyinW+HlpM2XYJ
V+Ynu9zy1e/ieNElXCeR4razuCWk/DhejMk4EKhlq3+kFplSTgArJJ8h5nRzHQ+7C5iSQ4rkzhZy
qCIRlzCyye6LZC4yv5DapHR/4TfFOq7hlWYST6zG1funHOHj5Z1Bo9cO1qpewnNLLq6waIimZwyA
NJxA84HTOF8/UkCIM6CSvZ9ayU2smQ5IbUwHqxBvtkoijajJEtlUG1ZSGWKzAR4WxDxAmlpJKP1A
35SW0IYe9RijYRaAiNhafiVXkKQ0ISlv5UDubfD1K/t08Ujz2GaHTUyL5zyCtdFc6u6y5u8ao4WH
+7tAOeEbyffSCjto456vXE6Ky8w0BIjsQVd5TP1FYofU7EXBKOqb9Lyb3gIt1PwAmoCoHP97W3ut
1rJ1qTb+LgOS/OmyvyEJ3YvAyQfCXtnBR/Hn6eacPipOZifXBWYoca3LyRX17zepHv/StYR+JBLV
j7LiY2cqkMrgngaBl/yCGX5sQFApndHWYxLh+le9ro6fSRiP2l//xqxponl4JPmx7PUVCvyT+ltX
aJXLBDZb/Jg7Yao3u8dCCE0syL5EsqkT/Dv3Gp5K4UY08aYJocyPE5jQ3w0Tl1LWwC8N7kkdn1dn
+RCVLVC3KSE636s6yXKyFenpOl0Dw2UzCnMEaxX6aQHO9SG4OeFGywoefnWR/VTiMzfXVC6TM/3g
EECc/vh7jL5psnvBGm7a3MamKr2kvc7NMsaeWEJ4/Gd4sNNBKxduOKz1CplOFMIsw++3t0xCZBZ9
Pqw6JnHmNoS1La3kyXTZgExD79vrb3YzrDQ8TJHeWa0RXTLM2QwU1EdBLIfVj9Ji5wGsQOm77l0H
5z1Wig/ZCNQKEfEOfNI9F+goZyVf3ST0R5+uEqokkbCX/0N00UZiMprtUiAPCosCSDwYGVypnmmx
GIWdg/8h6AXadmeineMsok0XMYBEeZ7ZC3nNrjbjsTw8VvGbx5pKAPnT2Ec3n0epF3KB7jIlwZoA
ea4m1Pd+lxR61bqTvYLFoL8wNV1xWkCPb9iQpwHnaQBAYrqTUdnpzK6HCntu44aFx579us1FV+S4
qH2MIC7IpHDZJDHfBAnS7jYJ99Z92ByvkjHar8xbuWRv9X5trVoSknR8ogc/869/lVYmJhENpXGO
+B9X89+Af1vReedHxM5aPt29kqq9j98ueq7KIFauN+x2Xw6TTWn1Ey3avNbNoCZsZxwuNO4STd8r
IsE4XsR53h/wAk/JvJV5jzk2ayjPMjAFNiOT51yUzziEUyeq9kg4ZeLfIstC1UwDSJNQ+a1qvERg
oMjJ63G00ll9aWCe7NYJlcgQ2nUXY59dBWq4yr6sSjv2MwmbwaNV+biyiJLl2poOlWwIVRSSJajg
/JDyCdZ2JUUbWIFu4fQqRTxXooxxYQZIfHH9pUuT9vWOs6SHX2eWBKda/OsWaFWW/LcFyFffjbEs
irXDpjFP9yDsWLBlOoVbRVcT090mZ2xQ8LFnvElMlbK9z7qULMD4DMmyUgnkJbaDKnRWBObe3pZX
0SkYhXgYYM/y9rTydeQFKtsgEj56ct+jJiM3NIxr7zh0On5Wn+esGzXkFjTMWLCh+foIRZZl15qP
Muk5i9NuXfRtAkqgD9ah7d633CMhdd7mgHyu0V5jxv3lNRGaA9BV98BOvcc1+F9BqLBgwh1vcYMH
2qXWzghM9JnEtPLPH5+4g/9PZB6iYT+JX8lzSyaJNtH0AxL6d6iFG5vVqMjcPiMVwrlVYhO/yMyM
4PqeWRsAV1Y8cMqDrpUvSnH4lSNV5Y2ELGNjRpUj4mwa4wj/9KURJj6MESc8IFqcxSZ83gXt3nVV
+1yBjKKv9RbNIyKNUf9ZTmOVUJjRhBH++Qg8K6LTZWiDdJjpRnaH5wnF5jXdPD7n/6LjQW+mZZqV
PVklSJFE2PEhmMeFxymvnILq5vasJH9mdG8Kipu79A4YhcBAH/kB3xJmOGik/sTYEfcfTeMXAY9H
e+ArzyGoai7aGIlTw/uQr7sEfLiIt6ubve5LkJgzySgq9uet0s9Gur96Nz82rXS5jCVutcWLqiTZ
kbMbtKDG92YrBrQ/hR+7+B9wNzrQ9wl0LmznIzFt99WF62GqMbZEFLGNid2lEvchDfP2ZnTASCOT
/RMi9Nc0DkXEGpGZpQrAai0jE6PAvlhiz85qXlLq2q0gvdZ0wSaMY9+AgLA+mIRZSCvqhXAWlNlj
4Hae1AjbzI3txXnxhMXWqn41+39heilI+se0fZxr16eTmuLYJdksO4Dht/4yiWdHGQxzkfUDr6HD
mlTJf2b+ikbqSiSR+YvWSesle0RJ85MieTjQ0Va3DusbfUrl5qxfiFDpQ8I9LlYOOpAQQnpzyjF+
Sw9ca1dR2wxoi+S8Vyy7TNYB/RVqJfZzUxbXZrEZciWnkeBllRRx09lRFC4YGQF6M4GYlGEnZBW1
V2/znKvDzJuyAQExYAiamBFlPQbZtrt789K206HSPtRe6kPUmfZ3fm1/uKX6Vefpg/akb4+Lmw4z
UJFze6sQkIptY0iKmDOiZVccMOjfkZ7SvAAOf/2eFCrMzAj1mgdXwmXmvAMNbJEi5ZNUI6asG1jF
llu4mOqPrdvkZwgG+lff+9Pbu13HrjznJD70hXMfhNbA9s9iQ4UClw9i/3fnwj5AE6OHxkxjx0oX
FCcjEWME469sysVQkbfyORi+etgwvYjC6Paarbb5ccgVDquc3wjrb9Wgf27PXdC1/C60+ClGxez5
jnKhy0v/cKQkRdAz4olX8oeC3BP2EVw1re2D+MOMDKKLd2SaQBtMm27LKT5Ue3Y4iiFjDOT5dT0i
vJQfhxPpvvwexAvQQAnCxGq4EU372R+GHk+pUdQIJdQ9rqXPKnIMVGYTfI2OsZWVnRKVJir2GQ6O
i53DZRUdQj4F1z3Rp4aPVDkHbFzI3kqgT3CawSWqIuXwyo8jlnfsBYVeSRGSA8HRcnloVHBvGEZM
9WafkRHImtggVPGp5Q65ktoX5Tm64PSEViq2cC34vVzfWrjAmajztxfmJxuvdIn4d7XPfUZSl2Sg
HAMT7eOfdGUids1+32DDFoC6POAZ+67kiZTlIUZB2ggakX5SHM0HKb4VdmSirg+Icv0LN6Ij0qi1
rq/eEaf2vi5hQngFD41/OkPtGQl4fASsbQSDYB4yo9OibUNtJ+JYTqVX9gkZktvihlDH9gIHYxhR
NZ+/2Scku+ByB0XhaUpn63xh5GNf2u4wF+DTaa+A54VHe9eWwbA610LsqtJEnHVQaPYM2Wv+t1bD
AHitcZ0ZnDsZOGgoPclKpWxsjcgItjAFs5Yw7ZgvS5dzJ6HIj5Qn1BDQt0BMKyfLce9qiT7RYZis
MAo1P1EH1qCXZ5BsifDqnW1X2nxAEqBoKbKG4KDex2DZs+6CbJLaY1iIoONyvlpZeC4kQbtf2Jpg
0qZhCATxGd7bz7/2hj29b+Ng0m4/ryOIDWtlH8V1rl4g/SL6zJuLuKG9uACjKfW4NONuHozyc28e
HsdIO1VfJZcuVLQGDZoyncAK/JiaUJbo4e0RI83mEFPa8LtaG6chU22hUStDpZxNKiXc0yhhplqc
vmfnttT2/Eeuagz972KRZCfDJvz+NOeOITj1lgMabPX6x2oxFIQ6XDa8Tavpa4pol47yemt0+zje
tlJ8YyVmuzZDp/qoAGWVVJrzT24lkdgi7BklipINFcAOPeFqxIyv9X3bE0jsGnbOF+suR55148lj
8GOrI5A90d8tnIN3n5hHn0be93F9ft/MAAL6ZRt7Qr2P9t4r5OH4YYghAr6yrS3JPb3XBAUUsjle
nSYyPKSRtdwxl4tCpOuQwc30gZuutCmtKBVhy1WmnjXm1bvfBsD6LzwYkEDwF2Z2PPiEc6bKV+26
KNVlLDOFEEFsksoWWeRyqlHl8W29oYxj8BPa4RBJVYVL8IvkyfHj8Np9PadlTdsI4+d7Sl36e1BM
50F3VImDn1wbHNtLJgHPHyzNL6+9hOPIbWNDjn0QZ3ggEPnvqsO7qgnHhpMr0IyWUtME3y6EACkf
dDKXWR6ccgGAldQoPSK3S7jIlpHGoUJNYgykdEXntO3MmSwF6x2IADVNr3cD37pc8MD+VY25AYma
nxI4pvhJkv7QMSy9jBRMrB/FhyiFqm3TxFVXG4az/2YWZvSaGHqLOOd1QkgeFlzn463NIO3FFFiQ
JtNJcdeGe4RB4qHemgul4OA9nwWyFPaNJaf1+F85jJKYH7HMdQZbx95fBq1Bi5725+cx1wKVcU6y
Lwo935hjQFIiT0mmrGsBqvE2y2L90r1T7dlWAQa8LF381c93R7qHqeAvd5ZnowPnnuBx0Q/rZEYT
3u4WVwbVilh6IuNTSN4mnVwevKTPrjOM5m6eiUziLaUGdCVYXFS/HxMUs17pM4yD4SZuzXSMEz4F
Np9WW5wdJGwnRGb79HKoqOmFrOvmYHO9vukXvP7NtBStU0VrBDMp+xECGY7KSq2YQnrZtKtvVQyS
VxrBQG30cAWFMonlRt4bomOTAjNwmYg0PiOMG4NPOKqnLTf67dkb2p0BrPMH0FyPiYmmbF2LBuO+
X6bXppQ0dqFIOf7tSfNe83q4P7vClKjtSWtRX9YSZx8VeU8bKC8S/kemX4Tvnar6q4mPg/UIviTU
AkikPfX8Vt0/yCrE/o9SkP3kw/7G3PqQhlYZ/HRB6xi86Q4BrM65qFGnDSLTL3dwBzOC1hxaQs7L
c26ioDClrlSL/UlJI+RIPx5h2ZKvqXZz8If4eSS56/gXihkEnQDJeh2TSOEsCcgULj2MDACSsDsc
wb0yz9L9P+2pZMevCbgjGWUptL3S7n3aqgucc2O8Ltw7d6IrxTv+MTm0/z81IXuPEpYmwou7O/Pf
cKM1C3vNwCV1pGAiTHsTZ541EKOehHEXhO3Q4ajQW2xjVdX6Tnsq45oCr/HrtYLRFGmxBTm2XZKB
yJvdAgexzgFOoCY9yeY/x7r9L5VkfAuLPzl52viywPnsRcArAIWOMLJ6rFgJa8FL+7mp87v12kWg
fgwImAVzGgFJg3hOxo2tSS/iuI715BtZgMdGQnpJxNqa5RHBc420svaTGb39pK+B/haiPc5//Z/N
MubDMn8B2At0VbfJbCyVWjqEmfveyof/iVxtDT/8N2KTkG/ZBwbjPRYKIdSyf1wv1D29wGzVsHep
yFsGQjexVBNCo1ub/PnrzOq+H+4W4/oChO3TjVZgzy/19cekeAnuykp2JoC3Dr+0ZtPRuMDTRPDu
3gaxiRCBOK+WPl7qY5Fn2xW9y9J+BMSpJ7pwqXTShK3+wEIW6ufaXprdSOCDWW3LTM3alaH7QSie
jGKfa5KByDckdh9rdel8vdv/qceM18RfWzD6Ox4GyczIY+q+/TBn5zqaX++vLCEh4+HcBLPwGKQr
tvmciZJad5QudGYd0n2msnnxtf6WWaY+hCWHaseLXAgf5oN9PCOfpdzWJdsbfX19VSlt0RvqU0Cq
EAxbuubGJbDjkjoSE+/YWvy49YwAm0ukEnM9ZF8JBBT1v+tJMXMLCUj+FtBOOtSsboXv07B7Wgmn
w7KKmfMhGLX/KFGB9K6S0SAcffe/+4U+k38s05buPRHzUD2hLr4U+c+z6NYcR36w7Laxh6dTI6JO
r5FW2wk2LEkdPKMEVXiELjgF5Ivh8Il6+LaVeu3tqg6DiEd2fpkfDKFG5RU4bc/Fm0lpco/GD7j5
CXAFHDF3bC9aQVa5qHIHmA1ztEaz9Gj+vpN3CgtFkYP3ltaN1oUF3gp1pEjloX0iJTysZXEbQHaG
UZCXqirHebgxqcM93mE5eKC0s6Mhpeo/+8J9EvHXI2UlnO/LDl9iW8l4SrVkUfw5prO7BMF38eTp
Jm7BqadgTycvLEkEGbmXGq6E30qUl13aU5jdZygn6/zzMPlLE/WOmKjSoyW5HTe/GxkjoTP0T3VB
kk6D4Xu5p9G8kVjzmGNKF++gtKkksGlzLMZbbU/AFfuUsP/eiFxNNWlqrA+x6x102DzhrNiOhe5g
jrp77Nl9zwuYWE1F+hmsmYM/seXjYXiRMzbEprPFmyoQ02gSAGUvirWWOH+Myx9pqzc4za3WH+M2
isfX9AY5pSFmXN2czdIfuQXz9nH7mxir4qOQwqALfLeqIoTYCvNpS9YLnyAliSGixRIX1/8OUrCJ
nGUFMVxWkoopy8VJxMGmY/UGDxV4RbkYDBifYlsqRmGosj/bbPDZ61xUiO8pKOsgT5UxsjgPA040
wgTC59hL0PggD9l/052l50w+cYmApssCPOhvNh6+QuKc7Xt6LO23+ysb8w2WGBzFjcEpUeyVtny5
EmVMEMDO9yyS0hxpmFdiuCw5g5lwJyrk0SPzGVRLk/SYDwA+RcqcKaPIpTHY0S5kaxKcamoAq0gg
oD8znwABffoASr0BAgApd1K0HVFJhBf0CUcn5MfrhnlvsMQJyampcF3fbRgY85v1yrCnWoaFqun5
WI1c0yIOXey2mTEP7KyautY4ZUWkVF3xXJW7sBi+wIeRvVbbD0wk2mBT2FV2lZ4kvpLAQfn2xqCi
UWp/oWJ2WEiujI/Nd3Tg/SCv4RRwMck7uAj4OQ8W6/OW6r3CHqcRQINMTiozDDQuUIMvbiHf4kg9
sux4M3J0+FudOLOF10TEjGpAsqNT4Gc08Xp9GU4VAysaMEj2QHX9Uw4jiSkAvnO9RUw8u33jubdU
N/gl9yUJxc7BzqcGNL3amGv1QK3PotkSmfAcKsaL2D5qerPe0xdCKQ+O8+vDkreJh/DUwxmN5mg6
97EdHhYExzIwo9U94oMG3Ju29xSC8l37dasxhT+2D8mGMomhQS9EJX77Tszv1ZbIGqmdfXBzayZZ
uY6pQ8iT2a1Dzgc399ChuLNS4zELEw05yuIOCpCSI8gcMvmvYqzfe3kb00+xAgeCU5NmEgl3tcQb
T+pFuUWObQQ6C7UZ73bGXji4YbkNWZEyjGSHIJVRwtPeFoqhjNEEEKF7QltHGPFniDT7755qSiRo
qBjNZ4Sup86V1iBdaU1W5m/1mm5FwsBbHEvjxXVCrXlGq4gudkZaJQ5uYuOF0WbrfLBRW2RvQehd
LiQA4a4k0kyoVbRWHY8YYv62qmf75SWNsEw11P1AIaNbl94VGDfNrChPARnUnUKs5sK3ZgVQPA29
tyuAmib3BJuU/8/y1h3poEPtdr1P4S9kQHoyaGbr4EeC/FlAJHZnKNvLHZNZFlnv87s4yNNT9GI7
y9xfLBIsBu6zTKoEplxfsoF3T3QQwO88mu40m1VjWrCh0g/a6ylkqCWpRKK0vA2WhvDxzupeyVef
nFGPP8xhLlSSScnGQBXIj2bfJdBPs69bMH9bpF8c7f3fe2PpuWfqbQ4Dwg32ir5iCE59gqGtEsJB
X8ty8gPs3tMTLuA55yau8fQZMFrWNpmXjdiZpeH8nNIjc40lKVgBu+DWo7APxN9kBADSBB+jORQ7
KrwdvVHfWuSwQ7I+VNcuOnenowXJaIXxFE91D+YV2mg1VP54kv4BInWk0+97mzKfE2RdHcSkMCQ5
4j5AMGfbietH4CLssOiLvaQaxqLBH5bTeO6AZGPL/rAQIarzBVT+jNDY1bmY6cQLUSPK8167agXK
jCnfvzOzQUnP3iASFkSFZQXl3GsaqhrSPVu1+D4l58ooGmfkZSbAjFPlyhAPGH4NIHqysdZPXE0c
ZP5zkpjyMsXxaOoIpB8lwcxOdwnacg1SQ862VP0QrB8VR2KtnrQ9gnc1Gh00J6J0gO51cK2SzeVE
GE2soGDb0ge3DnQqxUr1O5PRPrO1uSZJhGNUUdAbbPCY6oR5c1xcEW1j0Sp3w6nOiYwnT7CVn99a
jKINl3mKQZI/GDszcXP+rhkR5hZQPhOj2QO7AXXXeP3o/gGe3cN5Dj6Q6s+rxFIjci7zfdweTJIg
wQjbOp+M40rcmgkJCJ0+2IvfFpc4TSXI7hbuETekc5WXjVcbCwK89Gaa7nJKANXJ0geCbHxqZrqy
myXEo19ajwNGMLSguaq9PFeCxJ0WLqxted22kJIwQE8ZnvZ7buDje9quaFEO315bfIh2gWtwqbE9
4C9NBaqalIOG/UjQpdO7dsIhXs4uRMur0G5JkAuAJqNXU1GhYrpULO4LAXQk5+OJxXK6mnpJI2nl
D8Rx7clgIo970uJGkeWTbSvw6ecl69sSw/X0s5xjLuwzFxUkoen+xcr5FyJigE+lI4blfaoYb0TL
oRNXVfTfZymsQ/uv+CXlheFyaCjoiWd/R+uEczssrltEzPZv/SM4/jei24Id9zuBCEIGaSSUL+Ai
1uXteyR0eRrGP3tcE64DYHJ7j7/1riA73LkRLB/+VmshRUUru0VHCU+AqgVIoBYaivJ2qLtClc2v
/6dwsvtCYb/RDuZV5fo/gnDg6topKPblVTQFleUK5YejZ1UaKZ1a0lgcqfBqOV1YM0W7XK4bS6Bi
b8osgzHE6oEg50EtN6m7l2rMcyF6Y1wnLS6fl6RTcA8mRX6m84rfzJwTdkjLqV70xDsv75ViSyE9
fF1MnFwQtzXogCtWSdAUDMue16DJHW/Rjoy3tnTtZo6YLyjov4H+MovrUGMZwJpTE+aQpGE2/JTf
/UclxnsJUkZ6Utf+vuvi3CWpTM26RSqeuNWuGog3zfBUA2dYYzy/csSXs0+o70zA6dWA1g7Ui8Er
G+CqcfIQFVWaXy5sbHcXvtr7NkCWsSi3OjiHAF1k6B3AoSo3ylNrRbbFgcssDA1/vwpeU34pTfRv
Bjjq8PTbv+GRS1ym8s0UvuyVotzSC72q+L+UZfaXvzgPuBI0hdekE1WXayT3MVwT8UVc//zvgnRs
Nfw7A06V5i3qeTNY+USjPo7E+9ydL8nZPocEQ/l6r6L1ZUyqaNLV7G4wahiaDVXR9xZH2djgYYXE
slO41SKA5xhX08L5mZ+uQEH7fmlCJ0zHk9HBr4ZaClUTz5ixuAKipkLSG2CG3z4Tf7piPCkTxWOe
96voxqI+FtGmVG+2nxiOk3iU9hq7BdDECk1hXLG8ToJXGQ543HzebdxCnhzKPRKlT0MiqO5FyU7h
iyXZwxlFoYy8Soj0LZSx6aOagLX70ArIouKXjWeGcwL9jdTOwHFVfxuiWd50AyxdZuba+e1N5Y0i
y2zbpDH++f5mkAf5QemTqtSXeHlUtqVtUcYitaSejHDD4cT1BwmT1kYxMzl+9nitWFkcw5eSTuiy
uD0pu3iBFSqhA+If/bqfU67WOi3vMn4OnhSSN5hseKSApeUVJ1bnI1rjvi1/EB98RsiSayN3aw3i
7pqGypTRSXEY6e0yAadOkjsBaE1G2Vv5XuvV0mlXxPKu4eGR44ZzFAm/4xv9CxBDRmyCsv+kARMQ
/e4Ce8e++1IiqiAiiBVmcxIB9/diGEMXQrD2/2NUMNXb+EuETBBHSeJxMFpqpYOZD5jpi68yqn38
jxJSUXADu2w8gHehSiHy9bQcc1WxiL4uRw8WxzEB9jgxwS7u4NE+WJHSldzhCgJ5VCILa+2pgveF
JjjJo49/IresS9Xfr0sDIt3kHOKxl+shhopxlzpoOz6p3r8YzimycnLw9pPNe4atEaQV6js0lw0+
w76lLc1e6UYF/R+XHbJbytC8fDCCTiUg2cx3EWB+3s3ii9zKXJ6XDxJQmmj5wCeKN9M4Yu6PHbgU
SLDKcEiJktzfelCmp5Rdm0BSfOSZVETM4YSR1jL/POp09n+tKBWmd0NpdglGvONfPe3QIPK/4m37
OjRJe3ZOqiKQQYBS3gon3wk93NaQaCoR7pmRoh3SjzH1+lNKt9K22OSTvUZiyjbP5l4/JZxHjv6D
bxGNvgqicwoZxOvfKudDO0Nhj9mUyF8SIGWiYsJVi5/iiKLb3oq+z59kdRcNQ8T+onZK2Q7bcs4S
JSaUM4z1dBSlW6JkySSIv9XH3Kth8lVLLMXnbEhyAeDvegbbhKbDKfLJCcXYz3q0ZOBQQAS+vRd2
NFbRAgcXblU11sm0f2qOyKBZGb2Sao5J+X6NiYIWQW8FONw2mzb8bH6F65jNiZP3piGxBBtcYzeA
o7oWmoc3Ib+n6akT6jwmyxzj/gSWfMLZRgEgQTl8kAOpA87ZYWGsuCJ74I7q6/PzsDD9B8Wq4Rtv
cppbxDwnfFe+yJy1mZbESvo94SEnwjtIqHw+RtKLFy5MeBIbyw6GFlfVS2iRzeSXTyLs4HMPHJRI
z7d8uBpp2JljbeTEWsSiSd0Pt+cHnpTgb3jeJ994jFV8OT0nHu8AOTJ/1QdA2RZY0yg5PFneL5NT
iIRc6y1yg1L6uzJwt0TrniC6F0oLnkzCnU+EC3d8oG4YpK7HNqa8HXOyhSaiRunkRiYDf1EUpPww
wKki8fB5FZKaC3a4g6fYrcffD3C/+MweoRi2TIVysLVpnow2c6wzWW1/8ISUbP8u2TvLtVPJjyiw
68U3Ev3H2CsvOH5piKSjSRXcxXz4iFZdZGMzFM/xDkqDwgoS2QDbe17MRn4zRd0p/YWcSEuyeLqY
9Ljd5Lr7iOP6M4VofcKD8z9l4zq9LreRnbqROEweJsn4Ke3CWu1vTyzmNYovRoyNsf8JX5+ZO5ak
ggP4crxm11Lq5RUm+RdfpHxCVTylucqM+4NKOMLRHqKgsdcIfW5KyugH2q9v2eOCLnJYr4fGi8ov
AN8BiRKmX6M0oJW/DOEBvqgnx2+tqcyVqOiwgIqEbSQ8EVoZ4gOg2xwplfMo3l9zzvS8pChXtCVA
8AYJ/5wbAQ+x0NGGxalaUa1AvNoaMK7+n5iJ0HQJ9jrrMUHDwF15JHU7VlPOP4JY+5K58c3dM1zW
z+lhGUXTzWth+i/+g6rfgBl+eqGeMVSv8++LSsmpjuWVQSU/XRnrrL8Aw7Y3pnLNeN/VEGScF+bl
ZxzNMfs2nS7Es1ZeSAHtAHAsiiM1jaIGlWL42CkVo0Ywr8IArO2NQQtfFbOamwSoxCutJxtiHRf6
7BJPAUiBLZS1e3e3ESgvocpqd/a2LxFDkefPqr4M0U+JEZdmN1lDDmPJn2L3axe47Y3dsKJ4MRS+
HKkJmRYkwJtoXtOjtkzq04WQu/+5fmTBPGs/TTFq86p3w4ZlYUVAp13Djlo5frOYlI/WOElS+91v
GXQvyE8HqhpjSaq0mLIZjKm35X6RnwKWfil2pIADewUzU5NBMx3LD/hd3zLQaCAbpQk8jSjjAqwY
/0c4pdCJnnU8VS3I71ElKCRTOnYWckxGLyuv+ll+iNS7BJQUmqNlK4o48sg/hgd39eb+WLvmjJEi
3FxNTsdRyhwwJv+Kbk8zq0X16stjOST5jwJ9CZGSgfuHPtwPwkBhBu+4GnZv2O24putYan01BJDt
QXKtBrQUYtQ8RM6nIYZI+AcTAW/718wGDOVipdr22L1cTGsgUzyFcW/NuQnOjq0H/krR2G3+p+0I
oGo3V9WmQr19k4oh6JDVWyXlINVfVvja2UfltQlxxSSmEU28VQIL1rDPJvWPMTQUsqnogzkFIXt+
ZG4y8tp2HTpb59Od+Ph2EnX1YWXe1ltjfSSi7ALncOJWTjAxXKLdYAndCRLBcLrNjEOjV88v6bfH
4eOWmN2R7tFmR6DQXhiH1auVL/DWF7nqw2M4IPt5wm23M/de1rPOangNbQzlScS5kpL9JUbVUopQ
SGIvJBypZ4rnAFZUbNKOpkCmJnB+a1zZopYq0lfGnMvYERg4F8ovyQpjjTlF6V7b4PF0sSgzmDPX
8taHtcLLLhEkQKt3hnBMjDNMGNFfzabbAdAVsFIUUVK9OrtshkRmfyGe5IRKnR6ZtD/wC2WVgyt/
4+xK/4h2PGpEAl5Geyqi9KMVBy/loIGqHv6KPfvK8wkRJ1bgt82xiY5LyKCmclDx3f+zCxLu4GUU
VGz28b5D4MwJ+zEPJe9j1r6CbfVaRPR5nFsCncRiegu9OcHYaSo0E7eIJE0u1zsVPSGYpVnynPTl
W/pVS/9IVWJzYklY86vg3JOpEWvRQaI16FonJkDlriKC+Bdkc6WhUXdYc2nRuvJhVlIX2Ubv6dmu
s40WaWFSpJwo4rVuHxoB6Sy0w8ZHRROpTf6UF8J/qJpRlhuujHamOisa4+BkiApP91SfFcljkfAC
SupBD0mJQNv0hHMv0x2WTuFfNscr210mb/r972KAzKgE9/zHoRzL4t86y6tEHbr3R1h5VUbKLVX+
fa+M6gUH1W8/JkuiBu001Hqm6kAVAj/6HfalV82YIdB72d7NTjmBlqCSdUHr544vW/JvXnHaS64U
J3J2t1F7pRBgMhKYbp/d3IiYF9ALIJTGlEu1iBAK2VNLJsS0UjmPZx629thS5k9dRcKGYCIGd8mq
Zw9Bx4K3ojezeXJaFWqTuEc/nMwzcevcmr9dXUj1BfA1iDbHwbqPi3bTi5/vohA8gTk6NJAjIfGJ
n63B+TbiuLCWpFPEoCe3WnSWehxXPNWNxJaujxjIFnui2fHJx1U9ODws7UMl7xg50jMt88uQ67hO
Xa4NKUWt8HGFclLdDeWxjX8nuwuWyjWg/GhQVR8mhhiY0qA+Bm68LLpBgew+L1tW4DwGXJ41uS2C
oeeklW4IK/+On9svpS33YdOqaBD205FtuVIDQEfqEirUzYIUUwDmif+hxJT765XsYNMK7El73b9U
o2ppJwngcACJ0r+RVzXZrgvksfpckBr/UwgWyBcqQ2cHJMEB4QTmSmCOVMGoh2w92mcBZT7trPZs
TH1Lo7alDr/+y2ljfbwfXUnd6b67Ed7tZikX/xeMNSi2QAcWWlNYWBlNSSPD+ObivBKNGlL+Kq2d
+QEiAA8hx29Lq35ttMumLvtmUds2tVvNZ7ae2gK2Zp9QDL1T5Y6i2I6H9pmBg17qe3DjvCRnV2C1
8uhltwemDJJiYXEQh7Bd9fSrSDl9R3ETX+vyBb5U/UZ0YQqPUoJaGw0sfV4+dLnBa2iieGd7PZH2
j13WByYs/PVZOjZvRA5aKyykg4YmT1eUlJBTCik659WFrfgWRfr0TuZSwhv1ug+EB5UNZJnHF+6X
u7lnAOeD2bXrItxoQzzcN4iBBWfiGVhO+sE4qYWNHQs68VWQ8yuc/j/HqRKihsWjGi97CJ//Ttyl
b0wMnMB1jCCJJRSk1f+SGmu3VM0DYFRqPo+teygOJoP03+ElyWGD/fUBbKB1kaisWyUp4PN7oEDT
I8aAlD1Azzh/qWBsE+eytXAOs97k8GHAhDqMhxFMa7V64U3RMUI2LkL8Pr03gXPNwnKL8H05Bh0f
dOK+GEdZ57LPXqR9ElHcpXTQhMoKiQSPl3csU5HcodQ6458494LtkNWxFWG8TgP4Wwv/iWHYIwti
Rls6qNKAu6jeL/8R5f9r/ccwdJQbe+7RVeMcYfqwYongAWLzF+ABmCqZqzsAKIVu6y1Vv6S0vfNR
Xtk02DHbZgL+wGu4ovj8/gEsb4efiC89AkQN9S/Z2YA5jka46ghD4LAN5UvPLQPzWXxVGC7FFoyy
xQZNUWBcpVPnMsPWf7lrcXMkTHZilAnSfH5ECOAp8pt70Od4ETg18m/Fp7hI3SDZzY/W/ZLQaQbj
1S13f1eCTbkY5qqTXVOJWUNWnsdZx3tE+s5LutdfmvqwExMgHylCfZMDD1EKBzIGEGpRUGvfrBHF
2IFugRW3sqjRNg5Mx0v7UivgzG1YlDS0grUpYWuJ50BzT0TqPT+G9PEk7yNmIqusEFvCSWOp8bSK
syB2QWlBrvuh4QymoTFt3hMruWGJpN4ACbw5KTqVTUdvl9QNIIAXomdYqbjOdcBAHzEvDY3fJUP2
aAapgTeb5b0AmHfl9FjZ5+m+3u8g0hXM+Ygx65WIqH7o74+IU4fo92TPsQbDAdcMfNmIezk41EHI
4PuE+WSPAQjHJAu3+9Pz9hK3lIT+26rvQSx0cpUg0lo+QhWT9IDiFr47OjOqasor7K0IQa9nf1bS
46CEiGeaV/jl8QLTb6t8Th5Afx2svMCtyzThNnbvmr6Qm6oJTlXsim04w+glE4Wz9x7x8DwrE/Wj
DzW4jwTAjyHiNIQQTQE7/vLf4R1pKAhM8om/Cy0JRn1qyjnZSPVykbDxq3zpJOK2ri1pIb6Xpiif
8J89D81TORN8FT4IsNaAFUaGyKwPhWOb7SlVrbOrc/ZMoTRaXqgPzF1aqlD9LfAumAHZTtQn/xVO
XRoHT/fOn3wChGHHou6a1PUvJfisCi8syigHFvQTUJyQacjncGrDrMEAvPRtgUoKvTAS3RxhtQXW
pRrmpXj+DE63n86cfb7pvbRqTK50uTsc0B2vcVArj4TglFf8eZZYUOVbzDiFkbvAQAF8qEeWEViQ
92UZvH4j901XkS49Y/MTtoKHSiBzjpbDphR8LUHDe4ReM5F05lYsuw7FH80f2JBTMXpr6NPkc+US
wOY1VVlKWAytKHKaT6RLZlbuSbcwXisNBZSsq/0yfmtubgGvwLtNjjjYD747ie+prZnja4wIpK/z
MnaEk3KLDZoRhF1uO7SpVEm+JhoS8sSoemYQn7oswkNYVMk/D7S+LREMkuiD5vDOS+OYLM4gWgne
of1PaWfW5GzmqLRtWAiaITQZ/Xm8GsKwrs/ZuNMNiQmnAh7mRCN4RacUC1OI9cZ9jEZV7+oY3Cfo
U1J0k5d3zp+WygX+qQ9Azfz6WV1QPQWLiVY4WRemclxfDxtvtPWbC/BpJtNqbzTU+83O3Mi8CYKR
VpdUQybNmkgQ9Ou08PRJrK+68ZagPnh+Zfy1DggVIK2YGt5DtiJt0ytIyr94G5Cz6+2ggFw/v4sn
BFcytCxxCFOAp8hnzgFiZsk+W3sY522ybjFZ6bHfZuQOmyb6v1aWM+7z2OVainIvmYTtkTVgwOtD
lEJ4XI1tYn00PIEVep9l3FDivo2J1Udf7PqcMXm+VDtEPDxh1pdig4s7sH6cttj+WJxJVxk7edb5
lo/oizKxCUrAewyxkmJStUyVHwoept7dYJX9DbaNbNf/Pj92+ts5fjeN4857PplxnLC08Tmz7kkC
apfcbahPlmHkCHyEznwLjdefzZLs+oJS7pNLJL+AqOwk06NP2DxIIgTmxXLSR0GGAzgCUwVUB9Vm
qyOoL6B6UMnHcxuTjQVyeRF/E9ykPCIiOQSCZCcbNLwSs9+qy8V8iUUlENl8DYCf3fqbodH9jf8J
mPrg2PwYgf2cE73pF611X7q/yiNGGP2kKkt+TMEBvGasp8zcxSJbVIj8CuvMtaj5/x5MhCeMHgsA
0lyts4vNsmYpXK4Cy75KAr8hZcFsZhHhUAQj6I2tyWWSETbTE2SfmfQ1Aa6Jj82MAYLpkXh9SFYM
Kfb8fagxB4HafAkshRdL4m5/het4FQ+TS+EkM1WYZB2iaOWe9PGi3JjGSqLXE8mk78bz/FQF+1vZ
oUA+0/zB5FRubmc/6SZkAdISM4Tqm1da16kNsjwlYt58fUihdDo4DhfKu8wpAMlGXGD2m3b0Ppg+
rnJScf1w+E93UzaVLmiw5Ir7+x1drqpzJuwOFXrZYsT91Ai0eVaz6+lzGdU+Hw3ZOHEXC+Au/ky0
OW389gVdJFXCBdBN4J/Q9CrDRIVMpdMLFP6Fv3Tst1ktYK2wO4ozmUfZBt3AcHfOcFd4P6a/kb6i
dJvBowNGoBNGKlrxlQPPK2+uDbV1H9wZZ/Nj75X6UxwlybosPaYZfYC+VFq1A7C9omHB9rtqAWpg
vUZ7xY3W3HPCVriVtThd6BKr+3keLyBCaD1l2ujhvHqv9Qlau1EvCFN6yyPjjIUq2VewkrbyE+1J
wCXHGOhjEiqCKmzGFc/9JFOQTgghFkMD6eu3CWMDyI0rVVSGKt/wNFxMhiRpQlp71itUga6pIndz
PTMrIdQYeLe2d36UdeITDgcAHKyUpaIhB5unqHxjHcclDQk3ScTwjVz/gsE5nz6duH9ExZdQ+xsk
WrMpmjCFC36uHDXbqEPlKWFGZQ+F9T+RGdf+KN5ULRQJ6y3TX3xEbqzf6Em6OUdbX0JIdSqXEIPu
8ki+Yfo9ZnpDiCPIgN6QQLXTmIuzyYPERtDAS/E58yNV/bVaJ/xxS2PLXJ4ZAfhK3nehrbJP+XFR
ghFUhJR18cQNqtYCiLGcY2LPNp/gVXEpNJ7unC1i9YoAZ6XNUnnQCADfao2+q51vdS9lZul4zEqW
ObNyjDgxaafDWnK/jQlT3rPePAOIEfbN19pUDdn8vsz3LnPwr/fvXVsD5AWxvkfsbgZFmCO6gwb8
QyKuz4dME/sXiwbwiP8P8bRUwS3DGTZWOuMGMCuP7cyefZJS6bT4L+4YuZfCViNkGdbX2DA9XqqF
QD9Gx5Q3+l/ETr3mdJcmEW1PY0ooQEOXOy8sy4S7hgTkwVsCmVYOewq84iBwhb9375YUc0hdjwEc
kdrLltbUiGMvLUBeDtp8cMpDiwxlfQpnSSYYwDS886RKtYvoOfffXp/J680yrDBEZydo2ROuPBz+
FJTkqf8Hj0gHubONd9JrECAj1kX203WRwDTWpyF0R7W/6ukxgiMn1W/gJwtUq0ksYvdmcBOE/MEz
xa5j96LEbQdEwz2FWTO+ju42TBKg5V5h6RPMEqhJGl77Iy/aOUizsJ0iGZu06yse3KN+G6LTAHUP
gdMUfrIi7XKHkX9jTJW7e190PV3+HkwOlcIJ5iZynWNgYzzZ3jSZhCMlZ5kevG8FskgN6OwKSWQ3
oakNFSFXdnNyKAJvO+7qymlV/jWhRRVDZsz2ar4IKTQgChoCNTOxU+Q0gMY+MzwFKOV3L24+mM2w
4LEFyTWlajgA91ZXDE3gBMtmxh3jq4Z+joW8ARM3T7l4Ro+M2cphrmMt6AieZ4eoiaSCE7sI+kVz
Ade7HmkPk2s53HhR6UnJAVnMVf8pt3NDe2FhdI1RKhCguZZvw+XbrdKWkn9wMKOADHC+A08YMwdH
3PhAKRAQYcZfyvWGurQBaifjD7L9c7sJyFEjk8SZSisFifOVwsPBZibJE3HqrTz0WEhvKwqqGixg
dQKiV74tuirwx1EE0EAI/D9DWaGqp+bpOsPcXb2DWEOabwLJjtZQ5dAi6Od+uWEuMkGMG1vTBtnt
wY0IFdN8+C4qcZC1nbj/mrsAtc6bfC9cq94A37GUoVfudoanc5VTbLp7iymnRawRVwxcSgAa5nhD
ZylCx5YUrh2r0fPfPQzFQVeePiY7dlXs/8+MYIWLE+i+ju/Ah/48kDbPuBtv7fxu7MWU+bHexqr9
VVQMT8hB5NnkacOW2OCc9yqG1lJobBg/85ziwXLneH7HUsXb6bDcLVYheN7L/WogV7arFGVUciA+
Q7Z0efh8cFvXR5VxsRuRzXvaD39/rr55jkd4QlVHX/fImqm6NcJNhwyzvAVYtDyK6dB3RvMwZkY0
1QGVeESTMRPJkivgI9CY50XmI8+nDsmwkpzvD5StQnCkTNLjv6NTHiF9v4nqTSH9PULcusHmdLST
lRIbr1qSKKcBtcD/3cpcKKyB7HFeOPgdTNfA2jWLtaq35ImAHEMHJcNycm8op6ZAYO/5eyz79lNQ
xECzDY8in0lxGmNNKXCd24dgN1YdUmsYkn8CvHeYpP2uO/z5oQugAM3w+Aea0aelKft+Uw0pt6Gb
0Wnp4HT7TF75OOxnsoos1exgvRPCrQw2W9e8ZnAZ2UkKBt0ll3TWgmw2Zsef1zl7QPugjGak246I
LEgU+/FhsMqlbEFd/abbe2TWfem7tjAASDZYb/IQWPOFWQzDynyxUl/ih8zCcySvfx1jZl117ea3
eHp4N+IJYwCfMRx+q/a8gBd97Ixa/9RKLUqT/klWCqPFJiqpI9QsHs6JIWFdzg5wEtSs2CHOw7JA
ci+IRuvea/fFMYnRTMf1Xd4TgqxMBFTcNR7g+UXYKLoU8gSL3Y7NANt46rLnk9h/bE36Z9vERuz0
OkDsONZWZBEIoHhlOfdmfRxeId3MJPUIJ4k+XLz17IZMthf2BM71qtYSc3mkImf7tuM28oUSlD87
WdJKpuV8DsikOPfVEFaoRl6C4esfsRXzrEeR+cpP4ntQg1Wmb7yVjLUL3k5qAYJMuQV3Wt0vh+rh
PpnRnscpRcU/3Ca9P2VHAlaDDaLEBcYN2NICzgB2BhAW23M5OahhbmeMw+G2IVT1W1A1L4iIXpEO
GYNgyUJF0xi0n1woC0o5ifWh57asskog+p5NPJ2V6yZB3r1u8QAACyI+0TnBaIrL/82D5CtSQpHy
vfhAnVg/BDWyZJksSOnJEEL4L0ZuoyfqNvAk+cIR4JxiPq6Ue6VFLop0me5g1fytt5avgn2Os6u9
/1W0dUiOrpwsomm6kxWevBQi39rhBl+8EmAg5z7c7G02D8vzUogAyGLqwAX6DJLMmk89A6auzoe2
bGUeXJSlriqV0s1i999l+hP7UAxgftxkdnMdPFUe4RkgEpUrU3j4KdvS4O4FAWOEJ3fVV7YkIvnD
hSeneIeT8Ms+ZXugkBZwhhhMRLWG9ShqAXcidH6qenbunCuA+AXVF+aLH3zBxV7+RJtiQASsLWHe
gX+M3KzlswbNoQkV7+qk4PVeQeInO6NC6507JaMBkvE5+J3jdJbe0L/dADEiCFsCJcvruK4D6D06
1/J2Ez8QwZPTP88IrtvlRcIAmOYX9L0D2fNyksrQpzgr0go3d5hVbBTjONa13EnweF16O06zdG48
k/umEFcaFxOq46HVHbkpMmGVhuqJynHcjm6LiO94nXGW6nCDp19cw4W0rvo7ggIhSdtHc7zjoT00
FBFka+daG1SKfVpeQvuQsW5evlpdBlaPoddAb5vIsjCHwIhxLoALX1xOH18uSMBr+KUayEO82E9v
sg05gDSE22/FTK8j4nSyZz55YP8SyG4V+n7vMnZ+8dDP7Q4KBnqLYmY45SYfREcAPmSG6Jyo19TO
CIQ5Oq6X2eKZ49CjC4xtiXpU2Dm4X159qUuZvRf95lqPWKx09MAUS9sXh3ELCchbAtanUGZ/zNg3
8kXr6Lera1p7lC45Klx4X7Hht84dLHmBNKbXkzm6gIoy9FVRTfgfuRhZafjInziTusEJ8+44J09X
Kjeqe29+akphoGM6vTxDdnAUlKc6GAhIGoil8ZktZYry6PxL0gTZ2DAoaQrFNMQCy+EGgNhiqqQF
37qInBGicRDY1x12YePoVUdcExpgM3RM7MIEl77ib/RNUrxU9LZ+BP807Mm3fx1NTTJkfXHVt5vP
sNduhRnQ3zsvdVumNJG7A4aBWMgX5LL54YK9gpLZZ9LHFRR+XL0d11L0cBYoRhW92EPxmScagukE
6AxDPBy15pxl3Atoebu32oqm/IFoikNaZb51yrIlXga3dheUMuutRg/ctYsRwFCZPkVZE9sD7saB
qAw0WWrlJ3eo1ufFlMxU4Bfylap8tSJuLmL1LynbTCpgQOmtBRJYiNoMtPq+7CqLL449rVIGROV+
W/xy/I05WlGeFrqW7f8+N38LiyVjgiBgN3ASaJfMrCeE0yl1uFoqlHaaFFtBlCrw5qxhkLOUzW1H
vtYTR0GUDHVKr9/uJNAb6jdoq4slU9BDjOU3s9JFtjUUsO9Eluosz18tOAkj6EJU9x1iTV8n6DMA
5/mTkk0raz0oNSfSPgS3kVQ74uKCTI5fWMsn9haTWj0yGmCLSdb+MhKZxstJgxfBEevlHP5lENKD
aLk6EWFOkLo0oDCRUUJW68VsTpMzLvxETyFJS8RMNFTSxb0Vil+Qc2s+R9D73qTxHabWMWU5OFXC
T52yy1EucKcMeQW/6eY5zklP6Ole2Gkk/5zNu3qEkPy8yLD4ys9g2qg3Wz7PCqh/vFBWKRsujGqq
LgUtCXZM68IIVTBsEUy9cHgPqtRCYR08UbhmLBAut/mfBL5fKFAmL2oDc4qc6/DFnyQuHXrLnT9B
RY5psL3h0k+tHBwaIrSjG4IEZc2ExsvCS0m1uNGgb76mPcJrN9J+Cv4ypTf5mP8VOaf4Lqjh77V3
dXoYukvwpsKM1uN83giJK//oiTd+xtosvKkPz5eqAblbTj6UbiafoA8Gqp6u/k/Qm4+pIWZ2QTzn
Hzs9bFKdCT9uzAU8/nogiz8DiBGRTZCOlUKCZhTrnu+5DFGi4XsD7tAykxtfjkf8+mIsbgJYoAQJ
r09/+CNy6/452g47xHhVH4/JbC7p8yJuHWc73MyQPpHGpm/99h5RNOSUlEy1RdmrWJS/L4LwgyWH
rI89MXLNhNFzvkpxoSRD/qQr8TIjO00EmuR0Kq/Dhn/QK6YJEktg2CtgwFLRH8RwBrBpn6oWK4pM
W1zq1mB3jGPrGNAKOu/f3m0yM/I71P6lhqDATTKYl65KJu2fmFmAiKzmWxud4WGVOR9i1OxRag2N
oQRGps0eo8m1Zkm5ZmpQefEYQfnwUqn3zJDXjBUDLRNFZ4HteCt0RyHgcGf4KO4iaqMaY8VMy6MY
/suj05T2Z1QAwuLMbDijvLQRGVEN8gnpBOCAZ1U0sZB7N2IvElP6IXBPcYAhC3/xE8PMK7i/Vm6I
yfxgK1BbkEWv7fm4p8QoTsDfcCjitIeqbf58juHf52hx9IBSddSF1GLcWT7wnFVNZ5Auc9Nise7C
cMqgOwA37o6U7tkYmfD+77v1/wpOMHFFzz8tdzX1HlXECG5JLoNkNiU7zJbyKi5d7FcTRVuabM4L
9oCp8NegfHrQlA5mcWLIBngIlMk25aeblj3nUWfozssHtB5PgfgEnERYht/DWwf6Y0LIMUUbSrYc
Bpm0SwvgaCsDNtIdf2FKLkQbnT38qA77nT7o7Z0Ixt3atnpe6FaqV4OhsMi+dfESN/Hdtr9nwtVq
AGqo4XHAj2C+IuyEqamsIvRHxQ7aPxN5zTGbMhxFW2ZDRaS0uYylWXQ+JPVf3X3z8ET/tLMiRNeK
84skfyQl5BTdGRpw+kS4burSMwMqEpzT3/VEu07LjEPnzWftzPj9rtVtp7xKDUFC3RjZ2XJ1BDfI
qyXM2Lh+7s6BldcTKKEa5F93bJDin75vpr6j+ZqD5ZFyXBLnJ7E70a35HLhUFrKP9fvIPorNYq1o
UyB3iCoVwQU/1bH892DRqLCIkV/kyC8dfeXGrqWmmal16rzacW0JDd6Zaz4jp7FJzw31hd4WBeQH
1TAM+3ytu765Aa6Wsn23Qa5UxIsjYoihT/OGDBcpHwvRVoivQ1pckeOxffaqW1o+8+XJQeI9ZSy5
+k2ARKr3KV1cdo5IxMsI97hpKoAjx+SpFGkRF5bWPvl21XV0w28Yce7/Mlsu4dF/N8KWn6sTy9Cq
OK/xgiE3LkhEJaCiif19np9wvGwlkviJ+4JEBqnUZ+XdD9hbfCiQTemRiV/Z6W8OiNVU2mEImi7+
gPCmee50AlpsJo2rUAPCAnz/3s9AOw02FFhp94PDewh1BbRJ1hFckY7AGTmh4EHsiQTcVMueVTyb
cIvZ57Ykt0dIhXwVNJLtdFd98jm3ga83Cd0tRK2QEFIY38vY8n7po7tXAr/zLsVnbye8BgvqDW1z
ucZ2i08IJhZJvlY4NEE7BcYgLOokeInbtn39NUou42UyuYoM0tZsDGSxvMY4c/0ay66ndcijRlyN
QiRfWGsFCi8/E5y47l1bsFD6GvB3P2awaDemDp79OdA3X8SZNzM6ecd3FyelqJKY6nB7mDT8G9Mn
j82UANS1ax13nXI9v8lh9NDUwtCW2/Zl9H/N+Zl4ZnQP9jMfSDMTGQ2cOddPbPTfcSqyuBHTqVw3
7HYNyxCnHJVKzi5WC84bjz4w6lUdC/uR+CdPRS1slIeDnTSGjGhezkvzFlMuKF3p4jjAzPpjeb2U
Eos3zvMRf9FKjUFNzcEQohm6nVEfHCYeiT9HpKIWiTwYR7FehETfChqh5kRojGBjTcOqW2Bx+aYf
nGjpd2ZnrZSMCYgn5Sk6fgw1CDZdAEDzmRD8RHcpc6Ukx8KTo+cRjw4nvaVlAlki9Jg0VVIQbvuQ
bYfjFaJ3op/ZYlhFi2ZdwrL9Vk6Vyt+jtIksrlSCIgcyvdnCpRNHZOkuaPLa0oqpsuCAKx+niEAx
XUpc8WzXJvV0Rrtw/aXTtsotmytGPcvXkfhmibpzavMNzTkiVCJd7anFVfZ3jI09YFbVJqaqvehl
sEgTHNhjfeyKPSYUERyBrWEdexfD8jxV0QHdurFYVA7R4zPlaKIHB3jDP96qN//pX0VpQRPamzVk
tHZyknwfjH0hOCvBR3wumeMBMyziCdZPpgTYtbg9DbWncqewvpQjP+x7wCTePem5P47h5MkUt8Be
zJzQwI5vhVf8Z/rKtqY6j6oVkAs3Ckr+OKQdqZ+ASVcoJBGwzwcLsT3POhZ/09eBKm8LGqBq2YV6
QSTypMJiLvxc752VkwJ0WGgBwj5WqX70pt96juzEq8bxurtCMPgmUGCQ72JAp1/CraAkJJuq9ziN
ea+Y01RN5UCxaMCcOAoyMCYLoZfEPmyHs12Rh7af2bNZGl8Xl7hcPHlA9esg5tAUeAdfZTm9NJQQ
F7QLdW9hjyynOl8D6gXVWF6C2vlRemacAx1L2UC/yCDHEODEj3K7M5U97w3ZaFs6VLzs4y04UU9G
rTr0ckj8Nro0WORFlZxG3qTefLVB5jyTU5edye0pb9VJ5octD24w6o/V7PkBdeB/gOVydqDC/cRW
epfO1+pfeAMKk8kuogPGE46zpKCRF6Ml8nTf5fgnDnxWJjo42Qj5WpsgByxJg0N118+yndD03BR/
UvA0oFGNq6sU5jU0+dhN98Ld3esui1zCrr1MCXZ0BB9B8iEI1Dq4AUXzMX3QvQWIWwKgNL/LBDsD
/tuNnCFgri1hCZDpnEHtrqkSTc53FGYG4w0IcHWN1qY67jDxVCq8skd7HmPgqxygSmA2/STYac+D
XEqgIU7gqJs+aboOeaC/2IF+4eywb7vVYuuylmc36sjD28r2zqJUZjVsKT9/MXoQVRzd0fRO52Fg
kfnQFA++T1srCE5P5YRnGfp+5nMsCH4dXQIa/IblWH5sIG8SWklm8Hx/flRYBVntm9SpICi+x2gM
y+tPcVKXM2OXGvlUSVJnrt8kTf/J7svWR4a0qqDJsV3rh5sodn7zBB66Ob2u8K9v/6l5YS4b2GxU
e/+SPRbHu0Hy/oZYxDOu1GxzMRKP3uKH+e91EELGyZjQk579A4TW+ZzYbkjTAAKK/R88d8IQCvJF
YqQuwUET2CKGqiKo7ufkWUR5L+NCja0OJgE/15I7KkAsiZW+NO9xVffdT3e51bIQrldEumnzRsOF
GuZbh7JZXPQxI6biJoeFC3pMpT9t2qMdOu/gJ9avzWmq4AKKKuSrUXZYp2CjyXQfxfoTat7Jrshb
qQYsPPH57DgcvNEQLu2skadmLoxUr1pvR1rzYfTWhmo+FDtoCb0dM+FvRO6p3ddbsX/IvgzKk7F9
pcrbXn1m0rWvH2NZeuR/pQxSGS2rEH5b5qlkVbe3cUTxTSzE5dae+lYrDy38GmVaoiq2RzXqc3Us
40iMm//MGBaCvayRaQVN3svtR8/himiHb86/QKAtmGA23f7/Ua66eQG8xjHV5o+NrTxDrcYyELed
i29DbLbetJ4/FR6lUPikBk793scGSCVxWr8Aedlzuc2HPVg4N244DDbG6qWKGFEz9cYK13Pp1nn3
QVtbG+VxLh9MSQQMMor/BUh1ZqVb6aDlktlRT73l8Gd6J9J3B6D++9DzWhivKkr75tqR8bhtrNjy
0fy03EYY88A1aItQT7KB8AtTVz1XU7YlBmcjciAVblCgPidHsBkUe8IhmdT+i4Zp2SSqDU80NY0G
Szb9HIpQ0jruhQ+ss+NoLZg+tmX84HFoLLhXVuoTZIg+xV+6hkSer4CSKsI1PDDuYxxwn+OfQ2hg
Hz3F1gygCmk7SZ30o5WeLchpKqBuZ9Rvl1QRucmptkl/Rm5wRZeIwjWfs06HVfF4CbUbFjI3zPWA
J6qN6TNRie7CDI/jAETX+K1FreM6vnL9/oVhnIc/ImNlhJZYKXpL+oCnFQyI5mqRIELzAcMTSTTB
rkfslzq4+CW8aZbIMZ9ljdRMHTz0vMOgaBqeVaj/cjMBGgJ//cBlnyOAZlhonK9Rosa9SufVy5fp
Q1DUWkQLX8F/qDpCPKPBc0nK9B3fKiCj/GSveRQN0pbyZWfYd7bLYFXVeLszWTrLUkn3KguVpi8C
YqsoVg832z7nPjDnjYP8L/Fn2zIGhAAOR4kGkgdmYEFoxy+6EwQ/AA2Brnx0PE/lyyvzthK+qEsw
r92moXNA9kymTetlkqJNmgioIt3OQvfx5tvor2TSEalwmhFO7Yfzpr8/97TQJMYORubAAEZ5XM1F
2fCM6mIbd2j9IFKVIKeVOeuI9lh7ae1iAzNKtmjddaV3916Wp5evaVN+/8EROrlzcgITJ4FOWYBc
WN/KwmAR3R+MkBBlOdaJGY2hgLea379YXd1Bi66njWp7+QbnzC9s4L50+cQI+pSlsTvpnZ+xy2Qx
x+SdLvFxgzOqKLgzNuqjc814WNOOjQsuJcO3Z/hFsshE8KCym5gXy+ezVHK3eBcbbwL+4USBUmd8
/QttLRdpT3XFHZZk1ptv+Es+loBVdI39CpCWuK7Kkl0JgDs209chYY5Ve6+jUp5lWgPLuU7dBeLJ
OS42IZHEWtJeeu2o3QLDjHUiZbfUtGa6FizxJv+VGEnR5tyJNRqiXM8llj+uZgMdKHgmmr36bFom
FYuG91UwtbfULpbVJzumuEo1h09im5kb3H8uf4rjj6aeGDfpX/7/CJJrUECwPKM+ILJQoPu5Pptn
V41tiyX0IRL8i3Q9FP2OHq5lhAUI50i0h/dFs7OKt9DFo/UG48DvaKjKm6iygJVyfcfUp+qOHOpF
cKUKmrTo8QVmFFEwzq3AGfQN7/q1Ng55xHCDabm4qkHKCuHl0VJUHi74Pwo0oB4HGXlp8VfmCgz+
X8c0VEvvBYF+7NvYMFwn5UbtjCMfO1haeEocn2hsh/0yThNa6oaz7KQDhBUHv5qHxXkyS/d2oEmO
J2P0/OTbpodAz+WerpTi4KPCW1WKTw8+3Hjfc0C1nwzwGMsHn9UAvjFSHif72rlaylWDImUsr9NV
Dd950BF1aHbPH+TXG/VolzrD8g+qjw7ON5wO/tl7WqiJ0UTfCWIMU0wNzvyZX7gHUhrXVmNZg/Sq
8NZtbB6ZtZAOZMSbrlfJsE+l12WFA/h5bnIBIw/1q0bEUMsjuMp16bRgIT9kw7DMq8By4aoDX9FT
ZzvUe5IvCVcw4lCyONi/N9n3tGd4mBIrakXXkY6+8ym2Giachk7g1muY7ZMkIPeC0tXyJmrSZ0Se
7c+2Ha+1RtBwAthN70AHeEyPTJcnyHXfVS5zKlan70XKmiDKPGfs+zFR/bpQUZpVUvVPv9d6tjL2
uqlf9E6/+JOajIMbA4jMcwBxyf5XV64klHixxMn2jHvl92cdT58cCi4dhu50oVmZUSjXgwajPiW4
RfJyAT9KxKOLrsFKANE3+m+d2HETvfddCexG7B0xAaWLBK4XlCny5qrl3/bbUwGUdEtFJKDCasju
9VJX6c0p+egskTYp1DsNQo6Wj17UXH5AiP/16syjuRfXq3SbIEv6uanzcS80cMWucw3Ie4UkTgLX
b5pyqBNR4urRYzVLRWRYTWHOO7ZiyDPNJ2I+gGe1zPiTZCEOcd+1o9PdX8UZRk0uqnPaaK+2TzBq
qmW60JQczl5sL/88dMdVoFqKjRRznOJH+jaLLpFj9SCijgwA/QggaCoDpSWdu+Ma8b+QrD85c5RW
8EWDLVivhBfRUCyCKNCmP0OgyrqBt+xcbprBo3B9Gelr1eNaZkk8+rsxNYdOpl8g9iIIOxOF8M0L
PloJcjid8L2QgveMV7Iq9fe2iA9qIznYbfmxId/95M78PjnqnugsbI1mSNGwcFDFT3kfb/O68Vvf
1PgLfeWkxiS/kwe2+ReobEnwRjsTs/AB7scMUCDONzn6FmP2JJVC9KwD19n7Ui2M8vZhArQbQ7u3
37U7VbXsQOq4+O+yeZ3Y6EwgPgbqBgi2lOU+Frrh+/AXRYWyCba5jX1z30XYP8U6Au6mvSHL22rW
PFWbT/doAU3CTtzcAXPa+/PDaVbVmZvUbSgLbYEkm2qhevTaHjRvuwC8UegnGaXbo2Ng9c525yRH
87LU2PdhqzKTthIPLRucWZRlDAqe5nZB04I4xdZRO9sMyLB8KMh7mXOsBxQgHtmX0dxQr4zbgmh9
ju7ZyPRm+n/QijBVCgy36YzIO3WjWyx+XWLe9zU8gcyQJxbKPO16bLqNgu4dPayy9sm9JxEiXi9e
+FiLOO02V4QijmqPycHfLzxn+MTU8qfzISDKQFATkFp0fDk5skUU//IqRg6VF8VewjZTvTdlro0t
Oz29Ja33axS0GxoqYUotNuoVHpqvs4Vgm11thWjlViZOCqHbyVC1iJKLXJjHJhgNgBWB7+61HbcM
3+eHC4odBv0ISytncwyKibO+0rTDO79m2eZe4635xl2V6daivtW7EI3vqJTeHs3cudeBKLwPBcUS
ve37OO4tJ0Ost6lzcdOVxWhl4q05MQ2mGyZwd2a4KtIka7mGTAX7F2c6JXh6crQHt+Mh32/EiHQk
Xmb/oj48SvFHc5RpG72CtC1uSGrSMN1gv66ltjyf7xY/oJDOxQV0ljZ9vUH+FAR1ZRVdIk8bzrri
pcd4grHOwQ00azzKAxYaOxfIaNZkqzHdhHQtx4fYu5rFukGx+dWdlV2a9Lm//+KAw2pVmZIHjPkt
ALW5/9/t7R3/DdwWPuD9CjCWygiGcgn5b+ozrcwJ2E5O4ZePGlXvufjn4pTTm2bQziYHH1RuhGgK
uaIbxBSIERh+JzBVRDhicMBbpvVrZcP/u48Y1umgiZgY0gc0U7zCZtxFygXgBchV0lMTMn3fS1+R
/YPPRVYWDg6aSuJyu6CEUacUQdy490O30mjPOoTFpomxMZMQSrAw7iXiKL1UKLtsC6xI7Yzc9djO
5AIfR9kI8BX1b4CfijTMd6nvN7BOjSRzeDuokRJVMb+5mPSWm70X5QvCCLlqownVJ/OuPuQOKOPF
0fkIGqAuXjz9WV2XDQlTsCldhAykm1xElCHYVQNb9lgeQu8dU/jB8EpBlUfuyljKslw4Qx+NVIzc
L1vH39OCqn/Ub/JBnG4o4C5bDlD5dfq95Zi18FUT5qh2HbVct3lMAqOIBJsXENmh4+ejhniGaerq
uYdSYMmDfXDDbuVs8JOOX3E+tdgF+/GD8vaolv+aq91+EPhIGSIIeIvd6IWr20g3zcvppmUmbQMv
1lP10inK7n1MEB6qyWcOgdhe8v8EymN1LonUJIZJBCBBzPndT9fL4LyVKjgaNGaH8hTU/SkWf7ce
YBSFJUG1Ohe2AS0y4KsOhgnAXU6840hcl2U3jmnMyY1SOznfsVdKrP3i1o79sIVxc91VAXjcWu57
QnKtNGHYpUeDcqDJhdF6ObW/aIwO2EWKbKP7Hxn+rWFBPahrW1WNa+U8trl3+O2fca1ieJAChtlc
KMhznncc3Mp6O9ARXC2P0n3PNAiXzmR8qH2+UA5iW+LTuAzfpOotqC2jlKgP/YbJH91C+v71Njyu
S88ijgNC6rydIJYg5Ypv9Nw62IYMROBJwNfxFmtQlDoXWZXzzc02MnOHHR6f4JyvoCCAvYQydSG8
2feOtp3nAyl/UqLFJuXbUqBhgF6hXdniXe0aRmNnKXmGmgJ970p7JytDIQM/vntiriV0hGGg9wYK
ZYSTzAp29g228L+zEfY/L2YvgohSP0MUl9/RQDD4lURSSgDEQtWyBrZvmtN18O2HRHf4dyUtVCcG
Hqak3lgj3rJzojFq/HoGPF8c2a+vaNg8m+agtWVDLX6mr1VIuwIbjRVBwnncMyEgZSfNa4GLJMbQ
np23CPGB6ypKmXKsl7vQBplX+Rx2iYbnmdxQ4/QnF83XX3VfXKFLwDt0YWx8mIRqamwdLg/hgynY
B0PBJL89SDWzb1NBQcboTGl7GidOOzkD3XUshRrZpTgic7+pA47qbQFw6vH1eRO8Zn5KS0gJegIM
lEaPu2hRKQqJvZ5lajl/pMl0BP+VUBQ2ieynG5by4jLTGzrIfATaiCvw54q78O6WE/N4X0PKUY1p
3strN20kMn6181P41o1G4uLO1ZzMWpyaQGh87hiluBcZIZ/C+I4subTgpbhqDWIAZHX9n17XvcPx
kOC0KBxm8GY7j/IFowTgm1ODhsbwSrrIYxbOBWcTy7gRib9pYw7gqwQW2JhHzhi69X9J73Fn2mcI
QFVtKfKLb1KmLRiaqO8ZbqPkOWZ14h1FqeKHOcpjFh+AbCH0nxag70inYezgKNIhM+KrAZzsSb0Y
AyjmchZwUszlJcybyVgw9zaLFt8BtyJoXz/wm9T2iuhvpkmGPKkIzMFYNgS9EOXNgrn3xDisTGBc
1dceZKQ3XDAWb9PP7eylUzuDqmQH5JHilp0fnH1MwbAR2B4bueOBJKUOtZ24OvmN2YH5NPvq/SUQ
fg4JYoprmJ/XLltd+hEq4W9bS4ZzX8s3TMEejQyvtzi/tx/9vQRKAcWvHFqqOLtZyUJ81PO97tIH
yiPiO4pmzT/z5zsOqYdAfNkwf88Owvr5S+odOqAyPLg7zaLxX/GHR+fq6269MKK8qbKKq89LqS6O
0OXDrCCbJTKvjDyv5uo+qINmDjYzEtELhMIPfibrNvDJre1USqZwGmAY/4Szr1d2/EQ8pmtJbkG1
z1xeWgVqlJpG5u3ewMTMlt5fzQNQpGWlTRshGDmch8ilHQPUIBbfaKN9vbU0vqiKWwohk8NSgdrR
16fg6RX8viZT+OOv6YkIOB5EXreO+PPb8WHere75u9gKwsiS5m/ZZgTW9o3pCF/0iqKo8O6VAIlT
WcES3Z2cYxSGVAiwZW437lsoWljeIbFDPk47GsCMuGS+k0hH4QtKHWXHyE9grkl9m20kS7KISoxx
kONx8Qi89l2dX7iOlNLHIEneeqCdPGPEeijfDAr6JlqRJsXh7rBce70L2KOSk6VVjBlz/e0CVOk/
aKKaz06HOhTEMt6nUxQqOyffLMR3n0dK+WxOxfPJJT91i1qKTOz8zjMYOyHxvL9T7DNKiK32QBYX
k7cmakQ2hl0CXAbm5z/hTUv7/DQM7nEWs/UbseFgJLxGU7FoDkYoLwrNUqzvHIbO7Kwsdw7eDVgu
iSyIsrK53X3gaPNfU6OFG02Z9Lw87kOJxagB/2iY+jH68qP6o53jWk5bV+nHI2UT4xUt2/Ew6HXh
dqifXW1P5HTS85TQ84/sj0wi4/MbDQrFCFS+XllXh5QncOJXbkoV+N2VLpw7bOA3NM7vfETeD2aa
ZqjH8dMgqaZVWhzjna8jJiNHUPypWJdcx2hbm4k95XVZ1JH9QB2mA5Gyxe993v9R+WTY7UxKP3Gr
Cr4rQdFbPConiaPNPueiV+IWb462WgC+yj3e52gP7g9dzO+0738pxJeC6O7tv6BQ3bHk/kweX7fg
xiFmT0oXAbrSg3FtdzYlgYFjDCg4BWKnmJCuy02yhjmuyrAYgC5fxNiKbKLH88OSHvuMEpbPLxkm
UWsWpMK38KdZV7ZEEvwYmqoIsVvY2eW/4AZDA35P85e0shjknN/iYaWsxPmwGkAU235zvTYkZ2Kt
I80KW3uK7SJlZZeb7+MoJEFrR3RGgfwdkYn9rR7+r5YGkTUeYfwb7iQ2woULd+6xHM3UJB7nfKF0
B52BpMPJfjtNGSLMqOZiAjiEpeucLOYup/5XTZZ62Il28X9DJTfyY5pR/UxFAboVbX8MzFC5ur3c
XJq5LsKbBzZBCUQ0aJJ+zOiCmpyeUVsj+wB0dSQEA+6blPGo0ndV61LestdHrW/+BU0IIqG9n63g
UMOl/2nYgrgFTy6hdfcD9sEotsQvH+5qObNB/UEh/FhJkfw+OSO5w8v9nwjMrlvCVoflzCJGSF1m
QrdrJqSDaGnoud6kLSDHvuEIQIqu724cvQHbD92R2ugDT3Z5Pmt2pKVubBZOhGR/9ZIHJUjnJnky
C2wqdGhHSY+X47aEHO4A63CAA9JVQ/N9C04JR1y8WqsWohp3kc7kBnGQtbYMI99h2HR4CLiupJYY
TyPs5EO729awEcB9ui1STYzSEkOLTgEdCdd71adF6k0dU4WVS6XyrUbdWGFRsQs/RmK4405ELoai
MeSr72FRJ5mTwwGks+a/ra8bVC/R+DKEvmbl68J0rQe8Urya0bYpdDXZGtsXJpNZ/QOh24shUbjz
XPfB8YC9VUFhQhPBTCiTrM4UCqWzJGC3Kq72pPHDc9CIpH03JrQUkTiUfcCeGwe/MKzkmRyjJspE
UqbqCFbCzuczTRAaeg+HR/tAuAFLjNPmVn8HLaFo8nfh/1CaRXHUIEmIN1YLZGhGjWTH4CoFr6xC
ckuuHQ3+ytOy/nTpcEOgp32WLSVsUoggNdgdAPueQNt/YnNJTg1U9TL5A1aahDiittOWKYnC6jyA
dFwXwFmwARaEsRrNcOMZQTTQQt66XInaMTCaP1oG8mju6QbyfqlP5elMO/PF61A900uznYj3IxVk
/wmolAnw668T4S5WGrgc0tUVhBWZG7FRv+w/SMKOmRUX6mGEF3J3lEJ7Myo8QoN7JU5ehL6z6yrb
nmjC7wZIpPfIsTlLr6yYBGViDxPX9f/pW5+p1r8z9UZIZ2MZss2VtAYsLA7oiYWPcSfA/zHRuwLW
ym8CdFSwuoim+rB3T1uuQSVX6FVFkoTl/wXRIIvBfJ9dMnouyPqrqOWyCDe5/yNYUP8+viEjwK/J
NXjsHuxdOoJkUWaMMkhPlxuZN7wLzg0Po//bAcb6voE4MnsQOSNPz0NEpP2z9ttOUdSaRUaZmRMt
g0n2mQBFNPE5R9raQWmFpJAeClssy/Dadqm+wDijwYlnw2adTxLdjvnOTUC1z3xDLEE9Fl0DTmlH
T7yKMLQcQ0kXlkVmmN7avzTs1weZ8GcZt8G3KdRa8J0Xsx40pfdngCDi8JNuAhyF/Lue3jYuTWvE
9cA4mJOszcygSandmY3skZcf/oW5TnZekiDBXyy5kOxBXyFdGsq5p+mhfrOZTqnVZZaTo+gyM3eD
RQWYqPGE1Xa+3DAjmnQJmBDUJcDs9CgJe/dlyo6lEaCRmQsLbL2cank1QibcN1/sXS682jEn8n8X
FRFbHFE3Ptxl5ncT0Sv2reViRjxj2Kvatuq5d3slN4Bkw6ItGRVMehIXm8lPX/Ve2U6CdlzPyOpc
jGTn88e8tEBVo+ctSBvX4HvE3EceAtvKZabljZGsdZ+/JhcqlmMYjMg6j+8QZd8qLwDhJLP+P9KR
an5ywj/81qfWo9CZAdmOxD7oHGvrh4ywt7zFMqndCPmsobomqRWaOEVqCFWxgtveB9QVgSgTe1LD
Q/0rirhG5hrl9AkGcv56x4md1/X43HJieVoTg46Xq549oNy55rDdrSy5g/Qx6bqfylafuXS4CU/v
NYG6TyNWq0Rm8fhYAya53WjPHYrC9HojKN9ARUq+fc/gA/VepN3J1/2eXhsXTtK8LWtkRXGdH5ev
/WxcNbF+Zu3YNTX/B/Iqh/FZxEua+d047DPR2ILqAOhOzQ2R+s74LuFBm1wtgdrUeeWiDku4ymse
OuduAK+uubyQ1UypY8/fuDtYWBfd1lqwbt2qm/yR/ZCGK/F3YFbnID/m8mtLfrEIPXb918uUCmp4
utrOzF6ElbuXmM9mQBWwvO5DYjCIe06diHiaxZdql8g3Ouhiwgyypoct5L5S+faaaNhGNytsCUNr
HdpH4IigJ0TOX33DNKwI69u5te8qNaQoculz4qca/+klwSDwffnbwkPpXMNt2p9A9FssSy84aAgf
03wYZ81+9D4dhrHOjgtw2OGcjteLoLkGDzgDRIU5GZXvWEJBC2kBGK03eIcuuinXXofvZSMI+tGV
kbYxsXilL8/AfEcoGPcK+gzTHi+QEkXPMbaACAMzxf9NHhFNvmK/A4d05jihIPp7cw/xBL5/XNTn
L1OV8wPzwUyoLWnZHGuaUGtu0ZV/o6FNd86FL/kbX9bMZVne1ASV8sliptJWno8vlnvqB1TH14C/
rB0qYDwIPrVEPwkKdm4JuLSTazHKrgI9H0YH9tWAcnFSNJXZbzhiNTWMw3+ixk31hAWwIr89phqc
1M2do4te+QLWNJ06GnZajRTXVqhPy3v/13La9IC/0wKaP6d6odwNZQ5SOvnoLQR+BXbyzWFV/0h4
Bjfxf/YDS9y4IK0a7o4/L6qVqaQIs4qNcpMukByhgYr7YjJsGpjYIGSWa6SS4XALHR1AflVJJ8aQ
jqbX6ULhgB1n+mpDQSamKobUEETFlrZa0yp3Y/kpdZwktkfH1snn55thvne4x/Rhb8zTo59uQzTi
pNnw688/2fmOJnxPSKbIfpXUbatllU1KW6dRvDo92Q1CwDPTAvCCnfyb4Fj3MUPgeFYsOl82uVEn
a5UKNZL7XOkX+8YouD/jlCLMcwA1uFg1f6vvRQP9v7rl3jPQLbC5vGqA0APaTQGYhyhoq+gl5JPD
fxRYHDteC7YRb8GqZoDISYcz+J7/ohxfywI3RzEAs5iZQ9g3cSvVnNsIv72Kqm4BCUwuT1QbC79U
FElgar4bH1eAfzgE38YFiFdrof8GHUzLozaAC4YHAeUN8aqLBKkepoFQbokWw+85Thlm7faFPqbi
vzTgj+yNP8mMGgIRQjpu45x19lzvRIHzPDwYEy2Y0MWuXyjru2OmbbmTiDB1k1iKnXjaS+NJCII+
cd0zQQqQsdUS+Yc68Sz7k8nka2HX2BAHHqY5IuHDPs+FVwmupa6w/W5lPXztKtt5gbfoSkXT9MuH
j/pkKMAUJ8MaRWNRjNK8gJvzAPSm42rsWiWx8zMf/8xIC6Lgss+vdRCOCI0sS0LljqLh9641WWf9
Om+fQT2RcBMQiqBr5ocESWR4hnMSFHhUKFu0Q1fYntLowMrCkUp4dmJkJhHjQZUmXxuImu+aO+tx
RejuhDtRM9XNtbbq5zPNA7lt83uHL54/LqdZFGPcFbSTBy1zY+ofTAsYIHy4kWPkMd5uYT4TatEz
DzE2zN4xRd8+AaGz7zXB+mJHz2MGmulICtUNWjY2XH7gZsBf0em4pScEeKk2nwndNOhm+5w7BHpw
YY6eWFXguRNzg2zKp8KBvMtYylEwYxCNq1JrFS6A6/LocKtk+EafMnvTSVX9j6m+P4fpAoWWkhqh
ZSov7uMc4Pvd4qgLUpX+QWEN4u1iltCP8vV0dVSsl5L3ETgGeq+vPVUwxaiSWyPgamLK0lNgEF9E
RlH2yEbzC2xwYclla7Jxb3u4Gd56xiYpsPKPZWTKStQRSidtjvKRre6ZJ+pUIxcKpsTFyS5ZNl/H
c5ZGGDPbbhTz35LuqT0NGWFVDuFCGWews3YQtmi85VL8fr9Uq0+RLEwBlssWetXTfd03ruMzeCBu
vuCzPhDA7dmdJ82rsjMd/OLbo/78Bp7xr1FZOtz0mm2QAWM8VQNnxXJQz6Mcd17lcyiYJCmc4Y6c
tEcy1TwqPLlDjbIzxHd5ODjpcojhZ9qw9IP2nAL9XYdJ0lN299CzNcUFB1V8dJtv5zwAgdoF0QC9
Tw07FwryuQ3Z1qQLiHcHdpSccLjqbG9rF73VPejkThwqeGvTIwbCX/9aAV5ixBLH3NdBeld/eidu
dVv+39xzNPa8vLG9N8h7UZIaTdhlYL5sziogVA+CJ3/oM4j3qE86Y0hAHe0IxTvWTog9wYwtMeG2
okIeurFTJlNs8xPXNlWoE6moF52dphwgPJyalnmJreTitQkVcxRKWS4Y0/zTRlAE8VMSmAOMJHtc
UTzAU/2w566xHOhxVOBVCuSr5PrV0+grv0vAR3WT4X2thcMJi1uuXAI2PqTt4ugKk63f+kqFJY7/
DMsfHNMqpdMmjJD6Vu1suN3vraNDMkfVds9FhpZbqQpxTTBEGeDmdpBLFAMhSev30cF+FnbXcciS
CrccMcpVHgqZrva4jHpKd61xUW5AJhUgGcTRxfJRVzAN7p8ab02bmwUwd3VHZKz9ZnzNYn2dQ/fi
+ftId7K4haApburUEl5OmCyolgivTt1T7+eJfuz+f4GnqaD3iCgCFOVKgaocdPT0blky/ALLL2Lo
LK3dvsH/7mZYypV3bOG1SgUpb+PPOsp4sID758Szwwhwt4j/5gK5SJk3h8INDXv2Ob41xNDCW+nG
LzJDWu+ItjGoZeE+rUI39Pliy/8DB5NV03Bb27eHanyGB36J5A/6UR+1OUNSbjnETVBRBh9dTgvl
1mBDiinRcw7+6pzEAfkgPzHw+6M7qS3GqRnz5kZx+v5xcDF5F2P75pCd67J10rQDnkvdoIpE1cki
K+rZaCwfVQy2F3TCQUXG7fUIAe+nXH9nKzprKfUEnXPMKfZLtQ4pgTsx86JwEB6j9Rxhh3bxwpmr
+zUM4eWM7jEqCvL0rtCmP/qX2FFFCrKJtS2hs6V0R0D69jTmTDCV59vO/uenh7uwXOKryq6vgZNn
d+qPRgNcRTM7f1N3avCthAsUNOAgOsFndvO1B6ILfIwD5wyuSDdYozxFvFl1hcb8kxaVHB3HMF1o
o75wYCQeHUiJRimdvbAqGh+7IqQHqeWlLNLVw/5X0PFWBpfmDT8jUeEZhU3uNIeblKWhEuYEet4J
L1NKD6ILsERdMhRq4hjcHe3Zr7sVP5jPFanCJRs11f/3ZrWp815B71I2/piQZOs0PTtT5mVWAT3A
uwwGzLld1JUfJTXjTLXUY4dJNSV47kfhAUwsfGk+urEk2qNcJJe73ObbTbZS3RSkCSsDKKQR/cGR
WnQPtWhY12rkQVafpUtROr9ssjvYY7OVTEAjEFcMnJBy5vl6aS3RJXnN4eUa+vAg9MI7KUIzAEPB
HIF/jZR/BcF+Dh43Mhm0vtq5ryidXFmAIBIvL87A04/vPbqDRCtdvv5PcK1LIDIaszDKfmJqzu/N
/o8zBCw5Y9Cpt2tPBG2jPzYRNLA+WgbcG9tg039k0DNVUO0WcIiBNwxV4ejrghhOqMFXcj77JeC7
FPwZteTzNyYIV74nZwrDY9R7PsHCLEVvcHoUabA36JqZ++cQ2VlxAap9gB37JQRQZyLNX5F29ZwQ
UZFPOnRGy+HL8Nrfi1KMEc3Gb7empfeERn66ptKOGmQ0IQ2LwGjZz19yoqMgmPrvODm6gBS6AeZr
2beEOVClAkniWH7C9nbkbNROQBBZHANE6yPtCFZ/XDf6K02cNxVj/BP1zCpdP1+DxHf50XWMHeE4
9q2tWOq8YyXpM2/rEFnrsINKdDn3x3SG4+Q5qiYfLay/yfpkaIeSN4TApe+RGvU+cTxTIJZblMJy
5BJkz3NbkM4kzaWijyN6xI2w5d9BH67m1D9DgqfwKmr6/arXW1XTm2FApycMkj83/vEflrKgcAqx
dcESNXKRhSZ5fnBmrVT6A0SD4bs8qzJPpWcNDC2mQIGSmFfv9zMreEkX3IU87ba7ZzW7ei0eyju7
X9I7UL/UsK4EjhbJVa9GsVc/XCETsQK11GFm/sDSkg8PZec7BeCC5caNSz5VzK3WUHu8mrZzp0JL
vTS0zPxQgSlEciDsMYZcTXaj7Kbxlouuke7SA7hYYlADyYGW1YX+bbkHEZMRcrmm2BZWhwn8X9/4
Hc3QAJC+3RIYOszp9WUL4cfx+VB0fnAnjcZKqzRux3cRFR4NoXyxJ46/Zk+veC7HAyo29c2DZ8XI
RRheSNRrp4OFeSA0M2N9A6MrbuRm+CAsR8EnyC4jaTB44Qmd9+Sq9yJMlFsLCuNxh36xyE5RX0UO
R1n1HN/RRKpAeP08e60Tc5ncCsQfqgT/KCT3QSFbPo44VSoGCWyCA9M0qF5IPM+mNXHLOSVOyc/X
6u+LzRIit9IF8yzbFkCb89VTD78F2uT1mR/4xZTMHgnEvEV1JHortTQtH6mUltT/qr68LcST/tMB
zTPIDSdt8HVzpOnOSNkDucoKm0vWuxWXrDNF+oxpG+YfPXr3jv8NstMu54KHFHjSnf5FJkdDdX1g
Qb9gFI5qs3EJW69s8xIrRJiv00DCBsBfYPZ1D9eR0skH2vVhMdECT1DEmcUC6p1jfrEs5Aa7LHv/
KqfQtL9l0YkGNgW1i/Ui6xk7PRScnCqfXuuSTOcBMQJiE6TidLjRb/QlVEIYF12+kJlm3E2BeMZC
dJ8pYJGZxhG14FqAKZA1qfIoGn3jYvX7eLVGa5qsHaJnf4bMeQQUGfWZnK1U9gok0NBBCeEyzpY/
5AcHb8ZkQhogbD2mXODU7RIUipMteSkXY9xToIaXNJvc5Cah1nJK2COFDOYhjADvIrtd8A+/H025
E8RLsH5YueaeQj2vO7PJRLm8JxPoeBV1RpWpdzq83jKyZVKsoF5Wau4rCW3D1etyq/1Cpk4cOUTX
dOKZ1imZWZH6adX2gK7ykYSGZwsLqGE8PLsyDD/q8D1uuUUrjXQGQ8bMKf6bD5G8UFVBEDbB2UZj
AaDgzwo0GbsunyS7ixAcDzS078voQhgbPYsds5WHAcyl4spgpalqaJUc8PKmFxyHwYLSsfBDeQ04
Q8tFpRBFGYPZwrcovJM1tsTCBPsKccIz1xdiY53JOEXhXjFtDu7MTyYREFyMiLQgkc3h6MNmWRYd
2xarXEgKVLwVqenANk5n6NEz1AWDDSIswBV7Tp/0CsvfMXn90KugxpG462m4NZhdlLo6xB7OeyZ0
TUo5YtT0SuYr16jiNH5hAD5w4s4lWwoMl6pLRanLlJsu6/kcOrD8ZBh/ZNfTwwVmOiCQUTPtCjeC
ovmEyEgx59qpXhwEs4HBPLATO5SvHneZzfT3Dditw8EwFuXo+rm3O0tysBsCo9gFzqcEB4VyT71f
UKXUcY0A3ODjjXjjHzBzEqqT3NQE0F//z2hi9nuiNQ813hmjua/K6Oq3o1sP5wg7IYaFIUFn96eK
gmiqkQ17298KG+MaDNv7jRtzjrS+JQrWQC7/JYOlMGzge7nWA8FLeYmm19/vf+AjpZ+eO/RUACai
sMPUfWSMA6Y8Cdr795nw4zSeDexxbZwQyjmH67yZPm0KABdHdeYnjDBkKT+tOeObqXIUsF3kMlm0
uqYSU7GaDrl4lpThBaoc//gSFG0Hnl9XWaPyohtMQxv0/h89SWDexjlWsQpFdoM3Q25hrYoxe9tn
zRttAoVH/0UF9JhNqYTndAjRBxYHVmbu8COuIqJ4zwbZU+ecOQcFDzLkdMLzbD2tU+6XLktiNMDI
NueVFnpRQTdD39BHiFNATuXMJp84/1IL5sH8bqTDsEdpXDIuLHZNA14jJMrF1rjGOik+/K0OY+7s
hiOTcmuYle4HPH9/ShBnWK/ICvInwxzTgDgpo+aA6rbQhliEnD1ETHTpB+WT9XAwhlAxFOf0GqJo
4vgnq/GZRR1UxFWQvHzNDxLkJxnNG1fbfGPwVM2TuXWwH7chFJFFawPw0hdfdloLIR3YNQcl4Uwj
LKwP62u7YgNCjHQXGPyAHahkQNhPAd+1p13R7iELLB/+zvVqMu/MFSbIjFX154GA10PHxcQthckQ
7F4ll4yJxX/VmO3C+TFuMdkaJflTorl6kRaOUuLziGbWPIGcSkS5c0lDPxhPlZVVmzQRUpRm2xvR
hOpMYL5IAu1yT8Nxk+LATml6Py9o5P3ouHv20LNuTgQBX4laGKv8XkUnWWXcEgHqjKFCcOe6Hr7I
EzbRMYsEwgL43YyvPxgpk70AJL7Fw8P5HeXkr0MNUcLQbhtZaUuTYRGpZhpla8L0T0yfWLJsMi+9
JGieV3LAv2nj2tBFPnH/n/MT2tIeG0zYL2BXyowVIEf4gV38C7cYNECoQETHRpyawCI017Cic1fb
zlSHwZ7wv0fXgzxGVygvaheILrVdh9nDdG7F2s6Lr7MDBX1JSrm6qZEwcizPBFaUMLzqtZZ/bly6
ljpPPti+nIZmNAvtgeJ8xuZjyt5d/4b+Omyo3iOly9O+2xTgAbsff3rvb8Q9n0ZwAhG5NAr/NgzN
9FboK3Y0oh73ry5a0aqBrfDeT6ulGLit72dTof5IuYfFdN18HvNs9DzorBltcKscstz4CSyN5GXG
65M3pwrJT2NCA2/7Uf/ABeI2f+GpzyO20f70g2hMu6m5ADsjyXqk8Ph5qzaRXD3GeTXuuMTw4AVF
9Naudn3QJVQHr4wRbCLfViMmQ61DZjR1wyehc21aiDCiAQ1XpreoJL6fz8H/wEHgwnmPY3zpcXLc
FoWplssf4FBqxkUAWMVuUWUBicFA9QXUAZwHpyU5pE0TGwQlSxD9RFfiogGVQB43zrvboSWuX1Bk
QDQu5zWgrHuEj4ZUAfEC/rlsyl3Ooj54/yfWS8aIsStPcjaQu2ptZC4fyuDQnb07jfrcHoUcBAPf
jl/gVpNsVGuxKmxFz+Lo7IVVMmWgToygCEjXWZ+o/f9y0QYBRBvPNlhX+wUP8qv6d22GtKee1n/6
BPfC5ZDJRK1ylemPLxybUjzpfDAcCI7OjhSJOlUpr1/jDbvxzN+lPoaEUPVDVrwpryXdjQzJAqLH
yPc/iOQcTnM+UVTe1/S3ukPruiSiCZgEUw0LKdeqg6RwiwTpWajx8nIDhHEGY0XgAWQHaHGnhQ8X
6I7XISwUwyMmUUTKrbREqFf19lfwxTUswT3iRaSZK27lGrZyya5KNicFkkIS3+2zjnhafcahco3y
Fv2FO4A4fCn1Px8eygZzi/VbMU5ZTohZmbZc7IuX9/AP4KTboXosSGoT7VQz4Pwg9T4Mx3HQ8grO
Awn2CDUyHA0nWeHr+oCmgxP+bpL+xoVKhVNS6Za+HMxBTONDFcJO/XY3z8978KF74xeRRi5MDMeJ
Aiv4JeR94F/HsCNj5BHRxp+fMGGA9ui2+MgYLQXxieJaYboqbgKRlmkIK/LsXmU0coUWbaRoht7V
Q8hRSdAcsKc7kDceMZoOQ/Z2KKF5vqdrCKVax34cg6S90E8rw3sfoNbLYOhkkpmf2siuDfPZH53v
Q5mgc+ZMkQoC2NivotidCnxMlqOATxplJrAbUaMyjKDQPAUbYLrbJmpX/aV0Xyq1U1Vke/zjCzUm
+PVLfYAVCqDKCL+eGXQBmfp3uFKqjsNINrByrDGAc7qS4yzdZL9/kQQTicSeCBfIQsGxXEkYmS/y
PUo9cTxGTON1fqsaCxDJkorNz18wq5OLIM66LCQT20EOW8+/Vg1rPROMK1ZnqHnWzGi5No/NyOZC
+RoQUmkPtKYv0kxYJJqv04rrS3Ig1OxNb/+al1Gz7hDpUWsiMyfdBvCJk8Bmsr9odRIis07RMgOf
bezNBgmbGcfSSOXrG/Get/N7Ay5XWICtAYy5Rw/GV6Ru1U3Kp5DK6QNFSveaXyxx5kVs1V4fxzuR
IhVJhQ5uhUItsfE3B+ARbrv21bvgU7q+PpKk1all3ZyATu1cpQsZxlLVs5VUlQcizCX2b7UKJeOY
bucsnWKnQ/pRQmO0VbDsu6q4S65wsY8dSabEhEX/zXRFOMsEkt/MUdt7tWIdGrbADS+mHQbjoZqK
Uy6am/qEqYnJppB4oU3VSCbID8IWe1CV0jNF/Z03GU0fCN/Z+Fpny1vsnwsJpSGJ+e0Ihfbx9kwz
VYeCvj9OuQWO+cswOdM5gbTOrUF+Hg3NxZOazn+btjslFR5567TnHNSXClDKJZICqDvR1rpCC5G0
acfg22pYg4KqxzL1n9W5BMAHrSbbrK8bxqsCHpLpfzgXP6x0UpuV5Vvqcp3Iybt2K3NAUkrLGqA0
R08E+2eebvU/WZcHPPu7mnBwLzv2fz8O3+4AthOFKP7pnG5BfIRpnhdCzKwZaYN5alj8cAxGKhIY
HE52F51fBJ7R3PgNeEvnVqwk0xfdZ5W1Dzdviy7yg/1fsPjd+cXFAlNxT2WVW8P+TH41XENeqyht
Y0guFXfY09JRMM7fEjsNOlUg/GNnuwzMYXonmjra7Dr3W0DwlEj//tROgOxcU797Pg7YbgEZA1r8
HwYGetSi8PE+AY9VL0KcCN89E8Hwvozl7kzppgAJepEeU1iCTYI5qnLSt96jgwc+2Bf/yu78gnOm
cjR3btgkdlO+Zw2+LisHIcvhVEA2KHVUYLTefSiUvao6SGzIvSAdlZubCtRqS3volDB72ZgKbkI/
7MAmcqU4btso6xEHKuJd0cQBfKSSUQVel9aPhheKZWPmMjJICEae4Dm7/lKNM8QqjNAW0x/0PInY
Voof1+Mivcr4ozIhAzRpzEroicymga7qiqylzwvdN8CyLGPtqI9+ZY60+xUH1JOmtbMSJE6XfHlk
Dfka5IdTGvq1gShOdd8BWeQWo4kEnrj2JuGG/LWBkCOV5jpApz7tjlwpJDwocATsps+F9Xy7muLO
A+HDDbhAp8TRoXUURSaBWLq3vB7qI3zEAPls9QgNY9OeV3M7EF62/cZ+bzTDuzrP2iSoShQiyA3e
1Z9MR9lZjESY5MQsP+A5tE9HbI2Fv1F6R8VX/WfboSJ0eVqQXg+vdYTHOaxObGcKE5WnwPeKeZMz
99j/wmNzqV3R4K2kGcRvcwq9CVDigfUYEy64mbeSXEOnO0VDMTm/3Pgnk/UM0YjIo+X9aB+6TRQ2
0lvNiDNgmUBsXAEFJ8FYL2ia2uw5mhNWF/TuK77/rNxzaIorkdTJwSC7ZfqJfpaG44v3htelHhUW
HF7Un1QQBQzTzDB2Qa3q2AZBPdAeZbWGRmKaTPXhyyh/NSy7fJ7wGhN9KdC6u+4d5eIoAEaNcxvi
t8uXPqAnfWCRZhRipz0tdqk/cUOGPBwPd/lGQXx+UzG1CQPMpBRIy0zQFuOidNoC7zPAMKfelx8y
VfFHmMmctQeIIkc2c/yI9DzZZIsCSe8V8UQSSCs0rKwrjtsVeAbT7tCG5R4MB6yYNYHnkrE7iXpq
9tZ+E1F0Pea78fHE+wDGRfQKwspg647j8S++Zo8rjSyMM6MTskbBL2s17gkbVfEXfX/GS5FA8Adj
UGMiZP1Gqi4/UGy7cghzdh1FBiHOh9V64IxICj80owbphJ7MCzATQuNunSk5HET/XJDJYu1qS4oe
7YpgEdiP7oo/qPHKEh8STncgGc9AOm2+ZFlEE3W0vsiG+KMzpDykOcfHRqIC9hsuuCSN/YjUmNUj
vAEjAmVfXONHfBA+K70bnSp0+aQs8LSp/U0MLCfLReVxYrFCZbQ8I/3dnEIIoaI1mNYUebC+7PK+
N6xYmoETF/RSmCVUf1CPbx/ibnw+YhWwAbcJJwricH2U0s7u1znvOqO/onMUcTbLF4hxY4VG1LMF
X0oAKdZQD9TFbnWFHWViHGRD2FrTQkCA/dEJjJIYvItU7mJARwGupL/oCv+gkTIED/Pn9nSTEQwG
oDLdO4eJZHilHKaN8nOQUUFcQkVzQPSAjo+kKOiJBFRi22BUfjDXN4F1BI6lokhvlfQAwHISbaFz
SW0oY6WjWz+0wjkxaWHAHX7PA+VzwSmK11GqY6doJfkz+JCbqL3MJdz/an3hsktA3Nvy7xBvIh22
YgQsEGCrspzOhNtoY8k8dKukQVTG8Eq9vNyOyfjeY57djo1wAdfdJWaeDkthE6FNzihj/dxuRLQz
l7ists9Q257dMnf3AUeq0F6Mrz/OxhOVWOR/c8+P3eedVeF+qyaJ539t3v5+0wRZqiDsbGm2U7cr
D4tSMH3bUTolFT6pL98eHD1LQzXKdzIkpHngWCVKjp4bCqE1lTd3WgPp8lz4Ng9gKI7O4CeOdDMX
lQIaxrGVNxZ5a4co9gTLnLpwT8P0WWBO+S6Yssz/nWIeIzvwk9e0dkuvrExBLvNKHY3LUwby8PlP
995r1jiqntweCmwDcBNnTCTEFANco4KvsywKSUFfycSEm1JhouQriNiRQoyoeX787lEMNhlgjBG+
tWT3qB5EK72CZ7y2KhQhYnL0hacz7Hr1is3ZUPc3XdcEaiLynavu5wlQt2eFvmebArL+kIq50f9t
p9fcPlPvr4hoSylwNUVrAHioQu5PxFSnp9CDrJSi0lvBHg9NVYCfCvKg6OsgvYz0AKtT/N8zY9Od
higDWwK1DKtS3iDuh1/ijqOqeltylX76/cjb1awP+UXVQLa0g6+q/Sa8R/y3vzhZ0E+gPqIgojUG
Q5pWlRTBkJevcvskq4pntJb60Rbq0iPEnuhTkCVbEtqSGwG1vLgsCIQrnExYWlfNDGIDZuvDZbEh
gDaDL2RSc2wVK9lrVSLSqJXSO2+tgtQS3pMJx1Qs3rgLpeGwblSNOYe2i5um1p3CR2vlePVA0/GB
2P6lngM4onPB2OTje/5HC4Xdmy1BKeNnVGKb825WkzebCCpfvjb6vHD64ehH3rWw7aobH2qnmpva
deWK+wX2CK3HZtgxAkSDLNCJYnp6m7aLnT3OJKbrkDkQ9qC8RggB9Vl0LrgnUdk6CMrMLl7MMA0V
aG/n7DydZBnJ7nEhsAWMsjOAuIjZEQB4Kq9RLznrzcdpIOO0qnHBJUJKfb+23e5sJafrxSKQOai9
XSq720UMgtjK6uhYe2Asdnf8Cott7cS9g9snHuP0IHf6T9xcJoV/qSoERJgx88xLYQbHFklMODlA
mNRRsShdKWvghIiG9RSs8aX0rYbx6+78urTAMP+aeDQP8wfn+oh4hb09nfaS98BDRDHfwvLNI9rm
eBMSAexxH/9AyV1p5Jm2T9tea6YuZdMvAQJwsKS2DXfOCX4YhMPWwGzU7xKRJvOEIa/b07uIaMeq
otVBM+YL5H/MqzlL485w/Hv/Up09ahgosrht3ENkAzfBjz64Hnu/3+TVVwATOEC/Tq5GBxNORKFg
i9RzT/nCdBHRuutVtmTAPQTmkvZwm+TChzyfbht6dqLKXAskw4MgfmuF1VYYiMOlzdBa8iCaG4SM
jhkgpYYYgkV47oMieJkljbB584Wp2Glr5vNcWUetETiA50x23FYAoBLnGDH/q1GkA4SFI0uThlf5
tsoSicHT8eohHrAQgo96eUYhL4muFg0Iz7YMVH3v+p76i5ptU33Gd5aZog/bokZ7gan9WOBob5hY
f2jaDVicgBVzc+Yy/m4Yf0OUcCyUnRfezIX8QMSWQtUHUq+LR9NDRfdSJoi/S/H6kQhd9huWHn66
s/eVVIhEU66qtCBU5A7E67vN6teK83nRUasjhMEmntZao5pelM89wRTWvF3KRJvHZEht7HGhgSUt
0LJB28P/SHFmpS5UQXCnFq9VKyI5Z9QRUEZVjLixygGIx9zpLMyACZ+4BxeMA8qzlr/kL973FS0Y
ovhpGuU+Zulub3bCLQgeTXZTuiV22QWmWRqCurgo5gOeitHj2/IFKKeDv3ts8nn7REEUsVeHgvid
5fiJ7JqJeFunBHFAkn6chM/jPlwnzjDLyVIB8WkvL86eM492LqvbqaHId3wKHhqJGAJbtnwSWe11
1WszsG/xgcP8KiaZLhtFToGBPRvZ8rRlbvLjJgAc5nbfulb9LMzGrka7PuwR6ILlsrveGnkJw4PB
/nVD9HydB3ZiGUnZnTQsFjF7gmeKQ0grQs/+fdAcGI2wiR0RbGX5t+bkxy5G6l3/f1ymd+SGx+2t
3ZriRIOcTTT65JdUeJRYrqNPZxb3qmFtBvr3bz/PAiNZotYLKQ361grq5+Jhu0EOGxzNct9I3x46
/vve37F7HFmjnXarCg4N5Z5BgTC884LJL9rX3VO3RBwg1Y6gdlAUiyOsLxBkegiw2Yh1x1go8EFY
Wk6Z6PoZJV4hPH5IGO4Qyi9oe7d7UKWonf0c67F8+hA//yjDwIZLdGz92t2bdAt3XcNvreEABFpk
5sb8cOjncG6kXXwkkcU5QQWt272w+QJsmkUXnWWMX67SJTinR1VzEbw+JHNH38co5egQow9VlLWQ
jYafEeVcuqSAdEcLvkyRFlkwy9jeZxH4rjMoD1z6rcN11VVbzGXVchpSKHXmTiVMuQy//j5o2iFe
C2FjOp9g/O9XSmO9NxbCcXjqBsOeXGus+wG0p5ZyC7z2EOdpkwYK9rmh99AK0XXW8DIXaXaWKYgo
sLWsIYa+j/lk4YnuwQwnxpRGgLnSa/O24S4m/WHxWjQxvJ+XrPk5hJz3g5gR+YLQU6NjPZ+L6HDB
Nf1Dg6IdY951HJNzCKIIgPPntzVHiWy8nfcs4rR48mim8MPS9TU3YYUSmyXEyZsMkdKyapT3aJXx
T5u7NLrdJRetB0k8tngof6HsBj+7bXDbeguCy/YQ+MCDREgNiW+dqiN74MdbB6+in9bm80Hp2AVH
USdN4OgMJ21zWjwGO71WC1QuuEiVd55mEBSjvMO+xhBHfNUPGEmdniIXC7heLXTFlDdc0JSYG/Gp
wjBzS5CI+fBsWLTJNdoH2zxxmqmFn1Wc+XFBHu8ehCsfVcFY9lrrreeZ23YAcr+apqzTEkvS9iW9
TiJ0wco72vGRxHqMWDEFwqGDa82Dje+II/CauJGYZtsKcwDh/lemL2dkjttLngQuxa3Wka1mX3e/
XLdxZZZUZBkLUmrzodhE+6BCKCHkmuv9Rs7TDh2pqPbFcCX4pCBkSJjMuOkBnJu6+tWOyUbXtpCL
Xhn2mDh94ImymvT55ovQgyHj0XP1uOZ+qNhHB5vNfPLuHpaFfXxpII9YzONOAqFOHmEz23Fv4iVt
5gxQ6x6E64NNr/crBolmdNpxL97t8VKCsvPIfpmpeqPBbQIYT5NsSUBwazxBDL2U6TBcNKHnvMZK
BNyW1pYPuI5w8Ue1qpy/KE4D/EDk3F/2fkNDdP1I1zdIjcGUYaQ/WNwGeuJYazEGNx3ENflyvzpB
8LI6sNKZ15lOHRuMjFM8GzdQYfDUoC+5Ie2Yr4bxs0ID0YkOvGUfUOluluIxlwAGlhQ7amsjz4nv
S4lx0LTrHOZo2gtbiG75XXpMysEJhcUknNIUudEg+4Yc/OmSpua+QT/egi2gJE2aG/Ff5lvbbJmf
CaPMcls/5M8M+4VT4Ww4JruS39uLD7tsyGRvDRq1IYuYeayQhV605CCCDrBZzNMbDsLKPmmK4zU6
cGbW89GSjj3YUtpVq5o3gavxP4QNKrKs4C8Pehp7tgkPGEkf4ZPoIqJYv1HcJUcfBwdJzy0Vigwp
k4s9FvVxybP+0NsZ2OxSbmPEbic1ClyLUEZ5wpA5SehIvc+KxkxNMkUuqhqWUMzcujeP/6uNcTRP
GhTPd0lln5RsHcDORSvkjsJ5LiluYRJMJFSfY86ipWl+9TB+sYOSkdIkpk8ilVaEPvzhcUVio6uw
pOdg/i8/fibS2C00n+mKY0JNEfplusXMswifQ74nsHrh3V3wvlneMywd1qFJrLsEqWWO0xsSkrMl
AJpTMY3FOFUK5fXdMD+nfKGRvVGxN3xOlHUHaouCNXAUEZrVWd+4lJm1D+LEa9kswYtImF4ofnLo
lj5MARPisk32t0sC73XvKc+hfYzVVHn4hzCj8aoF3/wK/p4/bV1i2uR3jlPmh3iztHbgLkPyK7IA
CrsN5Sj2M4qYt7C9b8xG6ptl7/6JmwvinttAgPpA/IWsP7I7/HpDkm/r3BeWmZVZZ3rC8CKrx8c8
+YYFUsCtWMZ2DikvgnJMY865fMkWHjYn/Q+Z8Srq9I8LYnwvjRvo24tBahwB4KnXEwnRlIogW5ma
F4IuG6hnrTCjzIAIyNKXqn1j1YuKBsBxFSsVCW2uZwr9+8e4QVK6LVr58rJjANqPnHqdw+VmNzVG
uYacSh0mVYcjs5VwbxgdJ3VBukRxmg05QrMpntr1ZsYsyzmIrXcvANBREHLL95WgqY5GDFkBc08k
cyRw6AJDrF2t5GQC7iokSFyMNg6Tn4Za3qf8yvRdoT/TClmiKU85lf/NkBwjvG+klskWewu1MoCW
me4p+yKJQ6jiQL8O+1PQqa0WFa71CO/kwmU6GT2+YA++se3Gh0h9fAVCJSOKkPPAugv7/C30RcPp
Ra521CZ3BInFmJ/IBcn4XWtDkGa1+hLWm98IMC6DHS2gJqtifmkvpXBf1A1AWcg3x1XrWOQrpPXA
M7ImtFw9Vyvg95xqFRTgIMXCSV/PvqVtvn9VKhNpvJvipkHmNlR0ljN1q+LnT7IecywO3vtcLp5Y
OVZ/qXOUTiTtqyN5ET2hyBOpgYFfqQG6J380JLL6yOmRgU1c8b8goNY/FOhwAxMYEFA/Aa8sHQ7B
Ku1uhJhG7oNkgGCBQ2qoag+y9kjnYr8ykPwCU1St1t8+nToAvAsZ6Df0t9apOExWy8m1bvkQ5NYn
rbqyLl0vcrgEGAmScvfeXk0MYDSTZbmi2+ruMtbq65QfNCakNr+pHJ+IStLWGx7MyP1FDq95oCR0
W5SKTbBBzCYbVhUJY4HJSG3wx+2sv/L23nPSyNci5dD7py7osAO1WHde9wbql9hgWlIkmNV63t0o
hcW4+0VSCMg4KC5TOty9PFUYk5VDgkjwhaOZ0VU8OuykClaWN4RX1Ro5eWC15QsCMkjJ/m9eBMDQ
ncSTbX7hc/ex+cpsC2y3Amp3WdMECMFGr0YKntnBReMS1QhinvBMBxfQcSLeBIzkVCpDi8pRtaD5
TIPygwv3UXFGTn/fjuQf8s8o9BeAUJI0WPEYrykpwauM6vYslMcZvSxM80zBK5J+SYWECjON4+Xs
RxJeVfePTSlNHrmSpMw72G3QPsrZD1xDsTfYdbcq7xWp6f/lSnEIKF2H6VTTeiyCpHohPJc/erLY
Cogk9S91gRB0WqP5zo4kfTH0h+jCj4cg+Nstch6KCa182UAJUl9yYJj5lFDGBP0CvWm3DIVMq1GP
S258cd5uFvDr+j0IFwrNxA1YpufVnfsNl8hWi/afiE4jDwj+4rMgG+QdMa8BRkjGq6raJSeNApYl
OAGtb/GuiYBizyUX91DjS4R+fZ53lwm98hMwD9lUZbNgBuEDDkpGh6wqC7CCUoQHtF0dXhYNtOJs
6YdqCrXi6IQsbWAQEsUVB1R6TahHncFSkRpRvYF6VH3LTGPEc4NE/+MedtxgfKMj+SK15uYnmoe+
Q/ZkdvRPdpvxMvRvI54IibYAYjula5yd2llzl+brbGoet39jTUCB7zIHFKwifJLvpsIRgF6Nvdum
i28xmMEH3EPfzJIYSlJNj1dIrnd9OxLqhWVtdxCVLCOW7di3L5OonqYBySMeuXv3yhEfVPATB0k1
IJUCMJxIkX/Ml7Zq3WoDA5BPlRvZI4OLo0dwcHJCk1xPsDmWS4GRX75xYcV2TsqFURadj5AlZk/u
4I35aewe+NT4KG6e6PT26o/jqfOSEfqfX3iMuSWlb2Pwhp+IhYjRLYaohkGvTj/8ptBqb5GBjbc/
E//p8qTZnGK/jxsCECudEbh88hYQMIqdN1r2DXnTW+hpIGPqbOu9XAa7Zm2PNT59hp82ZrvJ1ooc
dmhD1L+Mh73rw41F4JljFshCYb4q7ze9UEkpkDowHANdlRzZf+HGkfha74GajRH1oEUqn+YqPhhK
NN+VRFMdI4/wytQ7hjmznpuf/NY4ZcKeOrp0ppudSGHIvBoM+FX3gdvMpTROjQSHMxz+XCjI1fM/
QOgCLHf2AgYlODfxGh9Qe9aNsxN6plHrUvAQCiP6vuXVA52dZ6gRJi0SG+k8hx8EyxAzs58wKXnU
1GKvDs43xtuaxb+kR8Aq/w0aJhTbF7rfghuzDLMB2ZCr6NSj6b3C3Ss4+FmHKyGMQKkPSkY9MBk0
vf/MYPyPDCCQqNEmevC/qDRE1sOUmrNdkKcEKTskARlPD1cF7RMRDK8oqhXkbGHdnAhvnBlalInI
WyAvN6vtbTsE8EH9lqNcskjeuZQRuvr7cisG8NYhBl33e7s4W0fW9Te+stCIBwjAde4CIlyfzT9V
Go84br7SXjsdT7YYBE+xLu05IZ1jQjDDQ3YxGL7s3LTupvFNGFzgFXkWslcpfzIiKeo8nmkeOkkV
9UCMe+qdN2Yvzvf7Revo72PFTb36DZPEVdvydZJIpfIGhuetxEhvM90U5BakznXAYVCA4TpHk9YO
x6aUbfK0nCp3AuPAZLS9dqrwXrYnHWHTZasvTRhzhYdEDps445hxaKoNPMLaIKwaOQaSG2UheTD+
jn5zJlfJo34ZRvdL8cCsHft+tBQL9sCwDghNK9sFNPChxGkUsUzlUPRu2IQDWKmaTJAwZUWb1aCU
uLVTA/meS9KyZP4cO7eMU02ulazZzguiO3yil8yX68WBXyQyv350xNtVMVQQljOt51QT3ZHg6UFy
1K7Qz/WxgOdcPrHOPyVkkKKgqkToah5rI182JatSr/e4/yGiHykKzFz9sWGe5FiieXx+jVqrPugF
t+pH6PFnbRmS2zzl9BziQLPPTfuufoSNmN8PfY4g9HAG6IpjIctmQ7IuSyr+KFOm8bXd0eS8gbkS
jXDVT7+BYyVd6L824hAGbead5a6x6vIT4hd6nUCzCwoWqtEhCxPk2G6ufrY5kteJG23evJD5XYmS
KtfpQGkXF1F17TpURUqt+UfhaKE2XS62Znxvc7r52Q+Rb2rynZvAQCD/6+KSQ/AP8OVzEqsNxzr1
WSYF8aPYWuakBBbMJKvmYI4ITU7T4nTG1ww5NbHoJDor4jYWGb/W9GIlAiHHdCpEcU8uQfKPCbsj
IsMp2XgbAxkr7HLHy0tP5yssCSiTm3fuSfDqOArvgF8oOtCBYwGIGt5yxH4kvHKa0f6zRFufUSaX
DACMRVs3pIR5mRURHSb8ITw5vF57DGsWIWkctyv8PgexDB6raXF904Jba+mI6eceFTJcUahcMqKZ
JRGR7LIkamFDULrAUTIw3WU8ss/KFuk3LdXEq04vUFhn99IezPX7OEgwiAC5RkcEZSX1FDTmi3vZ
C/Ibk7hkdOqZcqRZGaHC3KSEAq1L/HX8X+zrXcL6u3/j43UQnZufVkYnpiqq+xu1reBxP70V1Wju
dyH7aRC8F7cQ0pgubAcWhBBOUL0Oa48BnbisYXaF1dpZy3DVxxZxP3iTKXFaQvd10Nd3UMMTlry3
a5+jaws4bY8aVVxNaDUz7xICjbdCE/VE0YqNJ9VgDa3/tsZF5MhtCkNBpNgTA/2dGzypbVjlv6gy
VAi5G48ggAj+vECdCmfLFHm8vyZ8e01b17zZbPvjd1uy9ZVMEG8nfcn6BPOjvOn+QeHpmd1XKjre
SeV4FGwGQAQIbhHvnehNwncJO5rT0TsIn8BKDsfVkQI/umIm7chaMXm/XpGvajFtsuxNTD+TF5ZF
it/TNFuEO38FxYbA4ilnHvpEFCF41IIttA4UWKJfsTfnAYgHsQPte0p+NHxn9NBPLoldKn1YNNmA
fztWBTdYf3DxxR0+OckRVHP2uc+Yac8MeWlorvKZgoipR7RCZaAGscmhKwkjtzYh0Jo9JmItsBAj
Fg7NO3wL3B+lo+lZUU2IUTjEAs+ht0cjOEnoGC4yyLVAZtSp/OnydbmEGOKpXcyOv9V17wmWuSQO
TnvT+nIq5cxxEk08pohPZSSI/CUXYFIOqSH6ksoPtj6alyB82zFpmcVJWZYy0Ye77ZHQFFAXiZaW
QinDs/aahrQv8mABkGy/SciGkTuUzezrRC0hf3qYHM6UBe+8+59WHwKT9YbWWupKW3WRLvRZ/e8M
4TdOpW7x4Uq1qlddrgEyeTx8WDRLuBECyAw/hhLSZzvtxAgTYJ6QL+jbvBWsx9gZCL7kTsSuDrYK
LzVxhb96HCuJXlwWDX/lqRvGdQsN3WgteOIhMSXcDVLiX04M3JGbrA5JVf8e3JUY3YD4TWyzb1Y0
N3kpKe3/gv4DWYhPoYEwjeP25aqmvpavXGiTtUDxMAGvswzA+f32lNlvA913PlTZgU4P91eGN3mr
iJ4dRqKPjn5ULMAxlkrN40xh5UsbN2FdisjkueDrULdV38XKTOp/q/za0YstQeVzBvq2nZFHyxCQ
8miPGr4N01qCVru96ncekX+RsekBxY3UCunWkIfX81wE2vVIFlLlutZMo5vmGzWle695B/s4fy+y
BtsA+iVSQ51BNBtMV+TzlmyRWJLPX90MhKYYOe1D8OWx3jvt8AzIcE/HuVcqX+qwbr4EQhWmupJ1
D4CiTOcRc87AVgEbxlOYlH7K7xJOLr7lVB+mP2bN42+CwSoqLJAjX5JfnPbG5NmV9yYwKZinHm70
+KhHpGjA18lq47YT1HMoRe0e47wm8CPHYwJE04GiPQvKfC8/z/CqBUGDUNVowCKa9l9xficr6iPQ
cX/Lz3/lJIWp2DMGxb/atpC+WyjIrARtCxpvq3a0YwYKoG6uGbo9b5noLXG0cmuZROAbb+PC11f2
dx3YZdDSyR5QwiSGh2BLQJ7eW2Ri4GpcLc1b0EdXe1xgUUx4tIZxssb5vzWmfCQEWLWZCHHdUMsw
SMLOcG8tl4nUQMtUOr4955UwVNhLmtPR8tVduJHcdpYoqNDwjqvafhKFGwubiS4emtXeaz46VnM9
9b6Jrw4qWDQ05zBC3k/fEyzW57sXsHLgV0x5kHj9JA5kCbtjth05JzBqChUYY+rpYnQjc4YDmkqX
gNbkyHfmw/NvokXdgnpR8nz7KoxCm5D5CjeAgyg9wWhfJgNedILVaQWVPFNw/qZNF1CBIfPhAMRq
nPs3zK+1Ry4CXPui9QFGDR45V/CyuB6JvCMcL1w6foBfMTh9BKFDTUV8coFlKcJgwkJsVQNeAMq8
oN1fXgrN7C7bB0QkVyAHZqBykpkz/3oDK+gO/p16SVM/8dNqz8MmWJCED/A+SYPADLPb2JhpuwKb
emCXYZXpA+gWJO591QkL00PwtFIFRMi6r/oe/zY0i/RRPLQ3aKaxMTV1KQIEeIxrcu4CI1x53tEn
5u2/QAAGm5zMbYZA2pejlwf0kGWo11aLuw3j08A1241Ooml9hm3WrnBljmt3P1SoaHRZiIyCzb6L
/7VZFspOVx/dqAg6VYtGVCfHQBW0aVOf5jYFoS+d10c3jvmlLTujaOB+6y1iKtl80ReZW5G+e7Qi
6v5F5vOIsfQjPQIB+c289PjjVjEbxJD1yrSsRicuRci+6AIxumGCXXF9KyAcl4pluJyYwJjIy5DV
4RlfQzJ5NRIVl/ldKoWLO3LyuyBMtGNWNqK9iwv7lxUk7X8i4p5Ezz4zV8Yr1PRgn9mf64lNFuxq
ZPepfCHC+AmGlXW31i8RHzpICPfJtPLNNITdK9o/+1bwBrA6ur9qaAZZoqHyen91NHHbquSMZk2c
wp6SBeaDwFVLC6m4wY9APPsUAdGc1QH/+8cx+ew187Jov/zdgZefU8M8Nz2p7lRSBAX5zd8VIKEQ
FZcAUOtE6tF8kL/9udR8URgVkX089UsOPhAmcG1D5MuVhynExXJIou0I0oxL1pvN5zv6XmYR/IRY
JCEclBwlv+yc20CdJL6ShoKlokyp8B13bqtOViQydgYH7ygbVO3Z/z89Y0HBqs14r8ENDfELllwi
GAPZQiX+G83Q62oKFaKIQG4XdXGMtUsoj3g05bFlm6eCVnrxjfsnvOMhnXMPlHy8cs5+hkqwp5/8
s1d1UEkLlDaJVT3cnbINy7xogJcbM1ucuCUPyKk61SMvcJ3GTu6Q7umEv49pboRLm5cSVL9GH2nU
Lb5PayDkHXGRfYiMRs1FlXLrV7tqhD7rx55xIvORZtvztWPSXIoTSsthIYuua4F+t1ZxZuaKvyPB
GSXtsC+Jkyr3iUxVS+bdqFhFzNtKBFUQVYoe77vXZJzccF24sDR0w0DFeRsipnAlC+1N8YkfZCSB
8WoQwIXlZzp8nQib1jLdPtYcJqQ5JKtuu5Lx8jQmuTuUSd4as0diA7Vg6UG7Q6ffk0oZwb80hQv5
FYw436ifsGucx6B2lS54/wqC3+C/1dWOhYoIL8HRMRJu4OnKsKbx5UxhXfch6oOG0DaaUSNbfSjy
WSp8jvHOK7fzyv2HKIlNtVGk34DcXozQmZtv51TBMv0HIBBkN01gUneByZ3hnpzBgWkigPb1CMZ5
tvExpGDIzY/gkvoYeBeXM34083PZNEHUAE+ILaZGxBVYuDBMoyZTMI8elWlXPxJ3C1OhANntpXhL
sZHoryG6Dgfev53t1/wwQMhpNRiNbyeaQGDEPnLuejFojxicyRDQGIqv/7R9bte6S510HZfMCJXV
NzGv4SBkUE8gE5syRAa2/e+aRV1vuCJmMNHkqq8WHP83VyTDDxSsfkWGp4YstRgbs/g7srZigTeM
RaKld8q+mPEItpre8yF9Qhd4jb+rR3B9pmFyylLokW5fvNJt0rNIv2ULLkzTNU/r0hcswksB3t6S
f80g/Jr18N6+/uFNEtjQGDzXoeVCD0CKyntgVoCuNSbCL2sfZNmsqC8gLLsA46yupyC2gqErRSi2
1uKAOMwdmBe8EQ8kngGwbku/chWB/ES0jtWCTmPpjXedFZwnkOQE+Rnd+EhRbU2TsjzWxB5RaF8l
AtowEyF37Vo91giAN56vj6x+zgUxDX91OrCSfs21DM52MKFAK6qhLdGs8vVHSAbVgkB5e4prnwSt
JouXBmes0SLWtvluCdwW1NlfaAvj+Ol9nlDrAANes1q5OYlDSPECni3sJzPRmD/Q4NvOuYUp9mFf
T9DRQB0so1yeL11mSxMT2yKB6n/4bnnLgEER9/kqlS8zWzNwG2onrdWkLlk0+icljL50KRCcmDKY
2M8uPJzAOCPfySxHG0h9tL7NI8Y2WMY5eF94J8J/K4PL0O/Ywu0hBjVSpP+6AuQmrS9FPmbgVcJs
+Q2x4dmSqJb/GbTLdcU5WpsHFgM7X9iodAPZZbjQEYMhFYW2z0vxyC1ibkoamEhqKNIUeHn1Xews
iSr2on9D9tjyW3to5dtHAjKEJ6wrmmUWDO6EE7SaNbOJe3UAfdqDUBq3KB+mHxL+bv7L+wUyc6Ga
/J9GiohAHNcsj7gFCvTs5BvsNzzEMEx/0n0gl4QecwKWVkUF9AQn2P14vFLLzbReZpbbZjksjFiR
h+lPGvwT/f+U2Vm4XezcRXxDuS5OfNtTO63qYcRWnBjfVVnUpuMnHOBZg17iZ/YnHSK8DTJScZC2
C4aKlMavOxzvadBoQys7zmyxPSNkLbsKQrSoK7uIvWrWClug1CMIoit3o206fEDnSAceMclNAbe6
LWXBkHUWdVHkGVSF0XhKql5BZ1r//UoPt/x84Do7c7ws4CgINjnbraWy1VbKm3ds8Pcm9p1CtA7U
6iYJM2EBnZ/ZNQW9CyN6DWfDwsdtnsAdJkXqKxR/r9KQDLTLWpnvCHlcqYdNcu86C3fuWzPCruJN
gCS0LrNWrDUtAx4TSXBh/wM4w5MFpHXwKAJhYtEMzvlXAZqM6oaNIWdk2UxVLSoDTNha9dlrcjqO
5dchsw2Gtm+hGRk9rHU2lmIloQn6ALnk3MuRwTwHOEmP0IXwk6jtQkdO8VU9W5fP/wzOx8iS5x53
2iTtmF9UgB7wF7dymxW+l8k8BTEXye97/KzTXoZMNJYy/eQuvEcjpdcSvGtC0OLYdx3W3SQKxHeP
4ieFAcdKEm73aNt4tM6pOvWT/FXAyHzRmtFC1cW6WIct5+b2r36fta801Xitrte9qP+fJmCeBXfn
dXsIVaq9iKQB/gmpa6fDqd44YIBzuxsQ89PQ/wJd8LP3PEpSfJQW+lBAHWuE348edrJZPWveK5Mi
mdMpnJ3SStzzbAJqNFLZIQNRwlvXC8Lqwn/f2aPa5Pm70sKmA/5vFBnXe+XDLfn/5eR/pd95rVCB
GuT7z0XOEoHxObFH3kJmmwvwIqZkqTTxeke2Le+4xlcyMXFB1k7uRQcfH2FO9GDVk3cHns0s6Cfc
MKMLpDsX1cz3ytXxuMT2tEzwNNg78JNoIcuSenKphXGeajl9RuJgxVA7YxOmuxMXYwfIAfCn1dmd
u2ZcXDAnzmaUuhENruyF4VYT61S9Via7/0MYdEiKAUA2ZMcZgJ9755f90DhDxEdTGrjw8qCLqHF9
ikNdM4Bl0xzCaAN2q8/fjbeW4KNg2Jym8ybxMNwWb1CYn5yML6UrPr9Cjvm3Th7pzyPZJOCQKpsY
QNqElIRlkVX1zme4EUNS+TX3NQ8KshTtBDdTOzA/hGzN2dL9zrqQ41Kl2W4VXiJMDhUJ5VobzmjA
cwg5nnk3tDnLF3SxCy2J2vxBkO9KopwBadu0Aumoo8w8nTf24O7F8RcSf9gaAEuwvCeynoINffyc
6EgvI067BGaDuevs+72ynpxP/aP2aWtPiCs08lvrFLYDAc00lunGLQUTNSDnWsvw7/vUZZdG16nS
mSIwC7qJtDN9N0vDSpwqgvUntJ50cPrBijV+BwQ4G62mqBWC8neV9poAKPGCbgDG7Ztn1kAzoF/p
7yeyDoXs966q0Z/AtXAy5zQ7wYsdE7FCesl7iUXw+TPtfkKbjjdasN8OPWvREkTORWwPEOfarroa
+6DSE2+7aXDHn84sADzxPxQ0yIrmDq4QB+4zuA1ILc04ezIuyinqaRf5zKnz8XSPbiOz+gCOh3Tz
Tx+m5VcVamKVIkRei4a2UJqws7O+Hc/Sj+LeuJ8ZmnTf0x3DPMaVBk6Pht7R3I65mxKF3QamuwWC
S1QF4H+yKmfycczoF0L6WaUQZbaLuZQFD/rYcy83TXclo3WoCvFA9Nygpv5UXmj/ywAlsj1OJk+G
00KtBzCdiTGJ97+koEQ3WxtB+lVzMSoF2DTNDbKuS0hcFKGWONXo9TocnhA60JIMy+d3OlT6Kmtq
o4fEcPSRTW2am2bXZz/dpeYyvHO5QvWJ0igt7f8Fz2f+2wvBc9IaQvIB5HCsRql1GAMpgL0m1BnX
+9jZAcJFRWgJJ+VBletrGXv9LNROxJlNS+o6DFfM7yzy2G0qw5nHKSd/VbakJFtK70woYmRdER06
kJshyLgvmafygRlSxQtFMAuWtpObBK/DdeMPIMaF+m8JdZ2+8AieQMmWzjL/5PxmWlyxGsaWcZ97
7E+yUN9TsDbKSazwJzu3REmQD9w3fCEDbyxKJ+XluEkajxc0f8nxHKCqHVQmC/fm01GWCfVoIigw
dpdB+FrwgBWTIfP7A99gmrgLZCrmgcm0oBCFxhTHEuUKuN+dJ4657hRaGo/qQgLd4Y0KqiHVNVoU
xu0va0G429kTFuzkvPMSjhlIWvefsRU/YIyZCgqYQkUU+ospHa1ls401PK648CCYxsgti4tsHkji
YqQwGE2z5SrSP3z6gFztOp7/n1tGCcNDOmhWKxy763O7MknjCPFljmauIPNUufThRlYzl22JPvLD
hVcm1VDrhKasyHpHH6rqhuHq0y+LK+8Ugzp9t1vfpbA/yFRLXs8jvWIgSBklZsq9pEqAV+uyws6n
jUv5UoItLmiqqxXUqDjkgh/n05x6Jjy1FfZTZbvR96ZV5e43qC2p+u1HseyK+nOxVzLdKRP3UoXy
Adlnp/qtpfYPG38caHwkwDAfARvWpMmsVTlqqCUh8N/ENwzlFyYvmvObfUjjwhz91drpRQWW3sSV
6w0FmbjhzX9s7Fl4JRT/gYoLVFu77FeAunYxGVGFv4JZG0FBXRGRUaG0YufckFLv7vLkPJIRVtuW
D1PsrpLQatHqqjqFuEsR4m5Sos5VYsSbBWzsTojAoaGkwXJAk5t5pNnFmbLZU5xTfQkgWNqQML0C
16A4f8w3vYwJQ7vYUraFRb93f6jgzX/0bzvdD8dss11jSx80AiQvnnGQIXHRwdk3zO1DVyap8+CK
eEBDAHcLKDjK6XItNHPlwFCM7SkcLdh93yHjnjFS0HZejJ5HJjFLo0Nl7ds9O4E3jZTsKmUL4iW/
XKtzRwVm4Ibv7lrwSwbFFXwJC4I7qvDjbcjCMgCTaEa1RIkhYzgQ5Kk3cNQhOFheLd0wHFeGsEKQ
ARrPr8fe6D283RpHboahYlYBz6hN31moocXzt6vJGHCmIly14+fRN4qcZRPsOos50tn9sIipc3Je
L7ZouRpCUIlyk94c+94JRm5GrL3V0EghdWjz3CxcZPCygZdZOP7cXfoS1UJ7HJ3lfFnU9UzyoVAp
tBx3Iz4geJyNDMCN70vA0shujphgSv86UAvLwkzBKtbTI81smW24kbKtefrglVnPemVJAa+YegLh
RJcd1rE6yNaC0D0Icqtx8vzlEdMkla5oE6K3zHv8xYfh6232lj4UzcnqYH4V2g1uAi44MZX5qjzr
U6UYb9/TUJj3CKqASJUX1bYRFSKQyflyAKOT9Crcubd9XqZyj5zQ+mpjc/VSl7wj5XYBlaU1urww
pR/OHOJKNAcW56mjqLcQSv8J1A1F2WOSvzhvKWPKIdvHxEhZLgKCKZSCgq7RaCJOU+XxGLVn+nSL
t+Tz0eNWV2X7OdglYq7D7eOP1nL5CogkrAJcYIRLeS5eUXHb9d7gn7HOp0/zaXi6JIP7ivKSUQzn
k7C3k+bY87gpGPtoWrNZCi3cAQpBFjFpSA65v9tajDmu2cWxlxKtz/5nYQEGqSI2b6/TRGihCNPn
F4ryylfAILromYJegfWQZpSjlAzGwzsesP8hc5PDec+trcQBDy+hU2S2ZT3NLNyF6+5Zdkgu+PR7
JshWMYndyMyMDD8OK4APb2eeU6Ulqd1MVF/MODQhhIUhkRYJDaedhrW8pxt2Kq97r6H1luC5m6LS
qGH/w1KizKu/fWRwS6iUJGwCwm8ooTarNMIkJiognSxt0V51fYO7aPsLDAIwS2baLaEuz3yJMe5L
f1mnQ3nHYXbgH0AMteZJHzuy2WPC38cmAryFOyfbs7MbMrS1Q/HWEG2eQ9axciCHcde7c3M36J3L
4LfI89YECGZMaQlTnmqgielfJC7AtmOWrOQQb8YjfWC8jJJva2/M7n6dfEcZ8ZAMHgwS2tv64LeX
RP/DG8gBiJrunOA4twje5Ud078KJADd6J4O7Y0MKMmQxQ9HMZoaSQ6FPGZUw8iUQkg7GovL4A2eX
3CDfArKbNH+jHKOs4vZ0HscqkCCgsdMYz4meEBVXV+3r+/ecBYrQ/4TSLkBwvV0ITgpyRwHry61+
kJfxIpnmNojylESTrYCGTL56p/PtYjhD01PK+hVQbaEu0ESL8fi4tCE5p4XgvN9oTszMtt5tD5zv
y/PvHAqVksWdp4voEEXgJ7odlfkh1xdBCZUcOOLO2JGQb+zi9JhrR89hvEf1Efh+xQqJKFJgw81X
86D2yWu9XapkE0HRSdMZzqDkm0VGPOpN2Ir1jZMsQGmoB1EQyg7TWvatLj2NPO6QZ2Ov9c6CHvMR
D9AfibLGgEBC2nQY0DDgN9WMHRe/sE1Eocsc577o1+/DwSXD8lql2EeQan12emx6iWKQT4lN7PL/
5WuC9HlurjrQep9LqGSJ9wxR7wwgINT+P3/jin7P/7hghctKAPFBBI4SbCCk8HQXSIMq8EJFJOd0
d8zA+btEZheMenxfaH1zWMNWZKBQ+3DBehkpxJIoYYsnj0d6yMcsULx7Hq35P2E8dJ6Jzj/DBe8S
bgcRo5dTSTShSmPgmmiy88h2ZKVgaBwPtGjGF26PH42a5Cz3g1AaCzaHJLx7Cp5BTwuF7dGUU0xL
Vj1puJjr8k844mXGyjmp9rpcrpNpi4rLYRxfdqZICAWYp0jilRmYRSRKxMrZYTlubI1n6gZrWxr+
wTzPTBw862NQzn/FJzWFo1ey1Dwm6WzlRj1t9wd6n2o81qt8cP+lyeNeKp2lD2vbMNTwtx9j/vE/
+3abFQq7MQibUvK8/rR/qEwNBqKyTO5n2ZqlOULOD6jmkm0xy/UzBFgkw0OFGLF9KEjP9kWacXhM
kdUKKsShmR/JvsA2b2q+Vs19JiNVhNy0yQcrh2DGJGpZ8rIxrBkcetG9VWjDef15ZwwSpFyowwh6
HSBCkiAmVrhCsMi0ktzcRbr6YVVRqWm0IMWrcdPP2Gb/bZhA0hoKfdDjXdSAc1RYSCKggbHnNobC
n9gNB/ZLbN9XbgCaijXDK1zVf/4gwhm3TuShMxdYDPnXE/hOPbp58NjPJFcMwPrivjjWnU0bdhK5
o1vdjRw+A583bANicDEmB+31i+0akBppOZgz549DR7KjQ2Dw/g8cMtlTzyVkmYN2tkJuJERaW1ei
vk0J44xp31GSfm33Dj3cUywJccYkEBOTmCap7YzSaMBX8iIioBrZ6j/vGrmFp6mmvi2M0IX1omLs
FEuBLZjHYg5Gmp1M+uzXPnhhf1JQ9D4h5bZ+OMPA10GfPcn5iXueE8dkc0yBoKXucmizEyONuE12
CMi5mkb6DF5ToRLFNtCe/s5U5v8Yizk3BCfO9M+N8T0o6rAucg4PtodB4oA+t8ir9lyrppf7jWF5
HYzaORdRmNw88j50p9p6dScOkusTa6QAh6cjAOPSaxz3TOcyHWPBaBZt+vli6Lc2mbXx/mEXa5UR
fwLUlBkazq5h1XcR4iYHv8vZJjIHA0OZtwc1Kf8LdzDYVaYp4uzAbSuAAc53DmDahX/fXQo++HZA
kum8Zf/n3NndwNSYvUrmvsPxMK4wHdGTUPAF+6xBPkEjFIgY8tujbrWvlZdRsxR+SF1tRwv3CcWc
P/S0TSjUcSbDrewzFAmKnpFUTmJGK2rHDW9LgYvzIWWkcBsXIcY9OgPOFzXq5z6B+9xkcFFggNNU
+rqPImHhXa7p73fsMpvwF5lm/20urd+c+gFdqXi/wzYPP+6vmgVVIJ/PvxjraPOZmR8IRPCJIQOW
41fXHNVGcs/hDulMIEvJY2jmtdsRNH90T7va11DFbY+5t5nR71MWI2dRxkelmeDN9kgmzcz/kY3/
mCxmqbPcgDreEC2xc8w/eJfEd3FBJYcwF1RhU+JmaIGCFARZN+BJ9L484reHtnLVWw7h2vTInE8w
wLhPlMrgifICAZSBxLQO+eNeJGL5KgHj48qKlJusz+JYwYcJAqqeX/7rOty9djoXpOtSmyumq23U
xawSDGIkJNCKck02m4Zg8ALBx6UTWRlp7pZ4QFCWdllB99JjSfq+ct9ypgQz/rCl6RhcXSjq3Wcq
8YPVXJYMAuSTsPBrCZQSOqSdc01Hj9DrkpT6PHRqVJeoY9ToyKLoQHj3tMNVrLcQn5RVr93HgI5E
U3RE1UCwwaQg3VorVtsQ5g9zIG214zvsWbQpneb+Bl5kv175ajVqPFNS+iejiwsDlhTOvK2rTJDu
xfj3SKV770pYTvQHKz0R84X6A//dkozmAgvWQtoO0IX7rCymUwOJ4m9tx4uY4hIIUpCaL0RmHJzQ
Q4M4dc2jHfZd38PtxDv2C2qK2rp4pPaH2/AA2QvTq0cIuisiyxiarm5P4KpYFJNbnUAKRGcYefdb
o7PFWPayqorIBqVXdYaNMNkBQTp2GHq+rIhuQs7dLePePWvoVYivfJZkuGzkZuXw49XeNeXLMDES
yyZlcWbfvwC0ufPG1/VaCbxK/GtO/7cMrILSMrq0JeMwbJ9KLX5+FfD/77dYgKYGLAbpFN0xt5/4
btxB0lX3UTG0GtV0uKMDNky0HumHG6MdjtRdX24liGRghX945ujOjfX1kw+3ToK2TUYF4Ynap7rP
jcL6BHASbb/aYKAOmkbOY/oCXE8qFTykWAtBX770/eBb0N/7yE/he7wCjO/2d76Mqy+hMntYhWXQ
EeQKEWUU+wleBhYLZHdN+EbP77F9N9HXjhevMu50nN0eNdA7lXsrb8SxpGGXVy9XK2PkRSYgGoZf
0VJxy7AuXu+6fh5QiR+ayYW/ETdmM/bFa+mx70LDdF3n/8Ja0JdBn2k76ki0n7ujZlo//183zaSV
6d5g9ald+bs90zPpYXo9CQ2AJksI6HepWmrbi99W6JrdldD6rOOWFtdm7R9wB4dLTDfknxQAA0UU
PDlR0EBXkOO7YUsAn+gPXf43EHLtKSmmZoIuloU8ev+OhEqFCjK/oca9RaBiG4CtOG+8Gn60XVFs
3HmTrU0L53KKGacL4a+kbRAK+jNt/Y308Eot8ZGffPHIsnKAH+1FmJ6c3roDy/OyOIrIvgx58jhx
nDeo0LKnUuT+JCKCpJbWhp+SG9AK/9PbvIbZfzwYTTGF1Sy0v21vvUKG8b/6w4k8mJBl/q/hHEvY
soHHTSgDpVOTkN97INX//hbQJH/RgoYaAIFFJwthkpl7h8sOujUomQe9wGFB1YB49Inv0VoqemxF
HlhgGY3kiCLxEOOMeBBSzCgcQr5I6z/euyLKDvw3UxmhGzU87qlc4RAceaDdmGb1+E6XXOmFT1Tf
qAFm1ei+hq0mIYPtWAjip0HBSYrjVS1rJJ4kFDF3nAViJM4Lh9hfsRYLby5/JhuC+iv749MjRnxg
ianhVaCh1o+AvgMN/UkyjJ5ZQzw6QcWwluNWecDxZFQsv07uymIeygqDCHw5p8zlNLacu7PVh17/
QTCUyKAIdM6LK/4GfcARLz7k196PZA4VJKOefQDjpxDxZKsml5sIiOiHwSuHqKmABf6FST1zmBDB
ANoC2f8D+Pt9LNlYftG6XiIEdTk+u9NgvVqAtkdbMSN+EbwTvOKvko2+YSzohfV5jij4JcvKtP0x
Cyc+aUrcNHzNui4lkJOZatmkqoSoaFr2/4Abo4cG5qsshczbcZA6pxTowCT/WMR722heY27Vd5UB
TEOMGbw5uX+GNv27RQKWQckkbLN4Bx54rtaTaZ3gms99n9U6XipCp01JGUS+qm/LFCoI7sjJRklQ
LLhOwLdw9yCN1FT0pLs77uQigzBxNTjnHLyl3y+Xe0MvFFOX6OeuSYAVW03QwmeTr5SNEv5l8kuV
0rheuCFBND0B17QTb0hUAxH2D0uEniWlNXoY7Kw5oAo946bw5zuvrPYaLDEzEtW4q4kXuyPZaVyH
fj1oI6KXfx/1gXp2LkmJVfF3b7b/5niiFEaZNSqti4z7zRHu5o8kmVMMsaHDYpwFfE0TqaeDn9f2
D3AcndCKjiTbR/Mf6QpJc/XD7GsPDLLOSH/xzqnPVKCdep20UVcEtQrLwAHmwMDiiTQ3QldALhgr
CNWz0us6TM59tkIvvgbzGnDy5nrhmGDd3pXr3DUw+hm2zh0BhKesGtk7R/oMU9+IZn4FZsJ6pmsa
CBRlWAqO2JxzY0hH0yWB+pEhd/yHg/smXOGrlc19haX4GMhn/onDJe4qsJx71nccC0PMeLhqycJ+
6TD3PO5XOI0A8xVEpjuyWZyuVamFgvu9XzJRRPTJmm+2Oxp9haYpUe0IpiKCGJD/z5VB0Au8Pov+
uLBrJXcjHJFXuHpqiJCgVRLS5i9OBVysWpqxSkskED7AjgmWGGA9mYYnbEgmjaA3d8Q1ePHYFj/X
aUz603JFtF8/vbjeiPOQHt18dXbh1JXyqEk6zEP0dX33aYw0tpYkbJIdyu/BkoOVPxiN51jGiKRI
fqDB2z3Pes/Fiq9QWSoAinUrV2cpfT+q88MMTMfjXqPTO1fZVoEv7LcGaKKXQtwza6T0qkAfZu46
51DieH07C1IzQRgmABE/PjSef1gJ43HKc0Kwh6kvKU5iMdjYcZqjpuC9OvMqnnRnIqALps2dvs8C
3OPPEzUepCshRZ98tyncNXFqAr9qlVA65dLxVgqBv3UhFI0PJMy2h4Fqf8LnEB6O6U1nqx5/YE9p
qfUSWqrkj6h4IrUf1FvUT8ZMhoGL3mZaAzoG56YhgPm4gtRHu1wF2sCzuhPzZ5YgE1/5NK/Miihu
pGNrvhim/YCcxdd94x6BSaDPn1GWZf7pQwdt7kVPLuYeCQHpG8P16BVEDzIJY7r+O57WgH4L27LJ
urWhdHGVEpOqEA8AXbWkIMdyCt7pDwZbRuYaStBXhPEhPJ4zmn7KxR3HNakTAjP616Dzt9Wc2q7x
EaPiXExrPKzrl0cA/0qYjOivfsNEmKsW/4XGwVBElvxjMEmcbeW5/Ysjb9efhQXOL54vmz7mHLeh
GJpN7I0o1xmyLuAnscNgOo3XNkXL+p6nwJRy3mY/ECmpyL8WkeGOEMPQDsCW1Gp12Aa5vGc/uyE7
JltdMzJm/xpRp1xAj1ki/gL44PK6Gdid49q+VLvNQCBQOgwracsMSAYx4n1lv/zb2I7+ZhGXUp1i
a0mqWuXbzTMn0hZcYyA10FP5tFG1Da4Ej4S3tcpcuRjJ9AqnTjb0PAeE2o7jZZLeusG++o6PWuLU
HQtQXLhnyhgywfWyfwB0Utikr7U2pR5bKcGecqX59+bt4OFUqDFuw1EBcdevATNRXdDpArtKhaBF
SsEaV/O+ZhHP9Y9oBAVsqwoiOsdfI8vULEV9bxllfQxfiSgh8K5VwluRWl7SQ5Ul1blQa/c2hmYT
HlSGrZdPC4e1F40v74pLJCle+KMnWgsjp889GQrtkALG8+NjBL7pDbkPDCuHAkv3eGXtRFWP86zK
57BYHqNdPvUy3LCnx1LKgL80bqYu+bNzFYqXRPBaPvqbyFfaGrhpKMToo4GYXcovgNWl+EIUuAhw
vzl1b42u61Mxxs9kgaiMZahmekUO2uOAJPN1BFzGvPAvFE/ruhctQH7z84DHKgYF2hXe4js5Bco3
huVJGBfZByrZyWhF6c1uHk2QPzM3n0DLRyIuAICLWdF1tuSLTMoAUhHdo+0p0DnHN+8b9UTvXyVK
jdhIhnlmqjA2DojtIAuiUYvOX4NhMstPBH4YqX4bo3jAEL05WfW3VHpLIkKg78zXGuokJXKFgd/c
CdZlAjyvahhf3HcP1uP9zC7eMOAcCWxmdPile7oKo9mv95FoSfCGm09f4BzE+CrTrl1tFBj3pk27
AotJmWmCg39V1PmQ9PR/Jnx4uXmUp1dKiJ2zijO8fOjEpR3AeNwiv0xNasXj7rA0Q229RchxeGRE
9SXzRxmR8deFw+KSM6H7j9rC+vy/Uwt0VqR+z7/P9avcSmpSvFnkhEcptNFVPxgZTOmvfuJgeYSd
learuI5OZcZ5vrxP3F6N+ugcQ5G8fdp94g8svlNZH0USwPTII5e9RHSV67NxoPHg8Gn464RVAYM7
KgVqKNONhnF6nVETAqFm+IPM9YUli437CJxPjZqelfsmnvd1/S/IJePLxLmXRh3jzzHcKxKoNLOk
pxFQMHopao6EX+gnNYzMLgWLwkMC3xH/3nmDlEnZgOaBjj0+mpjr/6f60ua/BmI8S30x2lIIjOrI
rYd1DPfizyuOKW6st/T25+Pbl0krXRvf1BfbpXLeX9PlR7vUUMynKe9QMwPwg3QAU9tcjOdzlgBL
zgK0juKeuDxpk7GJ5ESETmQm4vYX8vujqCPIvfcFVJt05fTbKQu6c5x9JDeg5cFn2UI1uoe2sIg5
1YaFC/DPXGnWvkybotPuVFlqxJRDYjfqwje7Q02VcIrwBrYHmoqq6NecXxA4SISMwbaiqXpuSsOC
UaX8cIcloiKX1cZvQp26Sy3K1HGV369yof3m2sDARPXiU5slOQ83meMKRUWX/YMR5rqVbMPN6m39
PL9JWxUXFVDHgxlU7DFwblEgfKdLHPCMBBwZ8HZR2fPMlo7OHKmulj+bqWB5dUN2J6nZIhv9F+rP
7YPnxkucc9SyUYWh6orpuqa+hmDhhOAQxbPb6qoBxfNiIer32Ryz4bqKCn85OFuZyGzlZSl0Rof6
SAEHIoH8u3JVrld26fG8kcDK5Fz46VLy1vd1BFTkMrx0oWBsHiK0dcquGgvVl03A8K11dTWbq0MI
5mbfKPeK/9vA47cZyV3HrrEG2Ee4oyaZsqBLH04sDskSIn2x9DhrC3vlyVp/iwXbBCa8h0aa2iP9
uXa5Qhe2kaAZ5zO86ZBMSGb1MXxsV8WBsWrU0WCaeGFbAJLIVl3IvPIRuS9b+yEeek/sbvxA/vx8
LiXBwjpZJeHTJVd1ONJbP7poKP2sQxaIIkNq4o20/+hcOsRdRUOvTrveLBqc2275hoUuNtnzUuwe
HsknZAG1fdIepkOtmYcPcXhK4qr4A9wlG04j65sF9WL/ERbHCy1a3Ligj9rJazB/PUpNRukZ/EeW
rLLjs/q8j+M2aLJCYMYynKApWMIEqA9jUe+3iHNpoOa8c58a4cpEvaJHutzCb+gYMNsiJlmymaNn
ftKWZqgPlnqh3UrwXB5OP5KAEI5RtA7jdDYtYoljiINuvCe72ntPtxhzf2OL2aZ4RDN8AMZpJYPk
sr5bzTFpt44aPWSm+N/DO9WMSbSZiw49iXe18LJQMMGZaO0aCoiCFRabZtvssn15BysCvfND+J0w
DnlYU0EWComjtIdDqzvkRa6F2t/BwNfmnPgAtVjIh1u/Kv6kAnVEnC2bshqW4ctwqgb4Tkyu/Pvw
5llSqE+3kbiAvN4jbAc4qSd3mAsn9L/6gKeArhoVG+OziZ/4VDOgnwtTMNYnNmGA96sUtDXSp0zQ
hHUr0FgL6AYeod50woLvO5bA7tsDgEciTtYGGfv8BUPHtx64pmQkmY70YsU1AGZnEH9Pwoqum+89
UX9LGEHOKbfmY6pqHAhV2ndtAg8Yg3XKoxCB61haySCYoPP0S5MfprBAm0lipj9TJR3eXpBjVcQ2
spKvrNhbU6AbfqMEexuNGBQlWDiCuTnnNUw6o9jFrx1quRiYchBuiUtiRVSambUasq3qYlqkuZaY
BV6y/ZdGn+SRtvwm+DiKsAfyLi2FwQsevwwTMs06DeIRwtXdIOCfvu3T3p2e0BkCkYqz7IPpGVs0
08jjD8q6w9J9RVLUh7kYJPEuF+/rxUNGFoGjQkVH8UuNOdQUL3XwJl0FjZchRUjstVecGLaVImw4
muvapKQCtcoSsPLrC6y0Yez80z8tqU5rclvERfyy1O1xLYLCXbUmpssvFGPULGqIRSatOhvgzY5t
G1L+BmjVXaskJQIgxM7htNLKkjZguTxaUe6sCX1wF5f3azRZRuQYK7/bPLoy7jhzqr67QE8/0I8G
vggx/ZoY6Rrs51hCZ85wE0Q9CmgwGRm9cdsGMraPUn+vH523eYHZuLRjzngj3KiVPqSzM+C8S6Ei
gV6SxaEJS4h3Z7hENRJv1QS8u/Wo9hIZlyo/6H+hRshrSjkxOYcQkqRDkWYGq9A/BSIFpEZVk1b3
lDKVDlM3i49FQZ7XYLktTxMTfYkyfEDz9+yuwJbnBcDUoi09lsp3jC9x+YCtC5wTajQLO4I42yoW
n0CT5X00qaECAjprdGjZHrYGhxlh9zh8+NhP3PzTwQDb4o97zJ8KOStJ/d42s8Vi7bWTeKfP6AVr
5NwSmsFg2U7Hjq4Et5lpp5NyI2f1HhpTaX7EvL2Nt/eDRqKehskHuUhkdsm1McqCpDdxcKcPGFr1
rY0OikvX/zauOPnYweXQqIdd2KzUYrbZjE094QeLd9lpcdMapL68iMAwLcuw/gssUIdmRE16WNxz
vnt2L9IGxbIzGVn1G4QlW8GEAUlzit8h2WlTv+k9xnXvjQexVdND5sQkHU+pDOvTtYs383IRswyp
uzPxgCu50A16orVPZEt1jShWvPeV9WQS3uuyGe8inFVxOZgJWuV3ZiOF8q+i/5BAdi/1WvV3IwQu
aYjvRm5Xkuog2JZctrmzJYeRfL5p/swN9Ok6cPzpgZOS39+XjXKVNx3dNy/8/LOZ8DIH/rAK6KuZ
p8OQ7J+odo00tvS1eSnyILxf9Gkr5nvWaJlb1W/LQvrJwhWUnq9FzNLElgaSGG8T989wHtHtN7gH
5IvetmpclhRUVdwosGWfvSTWlFls8UcyCXO8jI17yfZc5aVfVy8jjqC0DVLj5hNXJ17cP9kHSiCy
Cs533C9jffxD0WWN9GDL35SyZgXZP4vN2njygrJI/ZJzUg2Xsa1saVNBmPqQUVQOd/0puzSuBp8M
W8rZtbVe4IfzZ7NGjNMVJuSQmgWrIDYa+4QeUWIbxpKh90Sp6VtUqMcYAOHDstov11bTBoSCFVBa
pgPFB9vndT8F/Cr51XWAZxfkkB3wJP5vRLUWNtNEUi5pz/HbX3yZsITa6ZCywmbZtYsRjznGyASn
cla9q7Ga7OLXmQgX+NrwBzXRc1xwI4gy+NySaRGxqxowO/EGcUCi6YIVu5Tc7pyN3I2LI6OxaM4v
cqnzj5+wLm9eg5kzsNomhPyMAYT1v31Jn0Lz0q99rpgkF87X4APWdbHYU+aoVYK4KiLZ2/cZMg5D
1ZJkWwkuGlD8uzG9BsBB7QT2VHucVz4gsY8bRg4qhivDLLS5kmIx30pXebKhjOTGIR5OjUAlh9it
k13hv+gsd9F9tFgP9PMsXSx0ZRplT4+wb1bCNTupKpB1d/sHWiUI4ghVeONK0lF8CUUvIm8OtWGe
OxXkBa8/JTW/X1I07ZRxeo7O47rwjgDsl8yGkSBfxQnvtSxXpfmu+ttnsJEBBgMi4PS3ucKW8czT
YRXh5po0rFMY7Rz/vxAvoMq7xwpfK+Swol0C4I2a5mG74fJWJTILJrHJ0pwrcy43/1MVEscd/DkG
DOBRMlijRqtUzO1Ka8ox8L1bgJHCulZsITRVYZB1OhCgxWwiSGBY8xI5x0d+mGyx42jotbDShmy9
BBo7hTDx90kJGqwWZgKxkBIi3GByYRQyFH2Tnr3Nn9Uxl7qwgjWxE+/ZhB7EK6GZZzuThgvVqkpP
Zd24432UqtCDCC1C94UOMfGITYMlDz3qvlKHl6XVf9lQi6+iatP5IKqHG5Qpi85920Jad3q39phh
/uc8xdZwQzlWPeVP+plrcNEYp8xHZ9yh+9iWiBrtpbAl6jwCgwyaH4eNvwIsL9hHW/5Yc9Ngl//3
EXpJwZdt4UlHziK1X9bmTC/DMwR7cAj+rETX3HOaYYEYLs1z81DxRV2u0NlgjdschJ9aoB0JrJhA
OKdHYIWnEH9JmzMeWs7jdnDYD/48ouXjt/Y713H4ilvpUGuEZQEkf/RO6/uiD/A46GAe/FUG6HpV
O79NFSZtL27WlCQsyKkc/Vp9sghYWQym9smQ3juNPDirFDIXGcuKcB69fKMA+GXkqQ2KPUtzRdRv
9NugDqvY2akOYhu5iOq9zhU3GDbpEjxiSe3xZsytA44B6uIb2dyKPzdwNbyhu+ZvVioacE9n9/OB
WgMqMUSD/OwoHeotTjGEukzvDB6fjUuDPJ6kCf8Aje8CMouygt3egFx+0j5MGjEvbda4mPLEzIZY
gcDBbHF1dSfek53js2g3Z8X3oieah5iDUD/RSXQJsTiEYQMrjEmHXMuFc6LeSB28UydR5fX5iNWX
tRn3lSPsIKJbGl6PIc5AwWmfD7INBllIJApz2iN7tFjRYTVb4DKaJ9LxzFo1NfkcVaFZkVkItlfa
XKK8td9KF8V/6nvuq6ocaESOPTEc01os8Ke+McOBE5/nVuw7tcClghoTuOq7CTtmRTZV0srOgujz
78teLSf8keDaGVxRVLVwl7A8b4WbsIC5A/mFwi0cdWbWZjRpaUxunRZEq6Vx6ewZNXK4J21k7V7e
uIXaxWlHPkuIvhyR3JD8ALhB4nJHj9mlVAY3GVSPO8KVNPFFABjGTRAOT6HpfpPWI2i1gcpUyNI2
ctD4N6TICj931epuGDLXU0hboMxuqgNFtqmQtcm8ANWrXQJkYEPSw5G5bbPNaZPuFU8acqdans8/
WLCSBfZJ0BlN6I4vKLAJqt/JlJu4nnfsuWImVbIvnwVWaxYNmLUr+IHcUWzPSGEdqTr8wtPi6o+d
GVYKlCkwdE/PoFcPB+ZM2n/YysbZ/MlbZxsP2rRTIe5aUUnDDc1RieAVZw049GkenTnOIC603jGQ
K4fMkQhuFYSRgm7l+eS0TG1B6J8/qEtn9oWlSUntL4b8kOjHiQNLjKniAjU/0rGA8tcHiiWHmfK1
qMLXsLESxI9lN6C7pCol9teLcEbIMZvwP1y+78jD/TjAJaAt/QX+/+b7fBhLbQSznCNYQRoYST0w
dc8Qhe0e8XucwLqZsdCfxUZ7GAolMxV+GAoaL8s9UQLlvpZdMFs7cfkcFqAG42Kynj+wJNClJjZv
ElmXTMmpExqFp++n3qOPTF8pGbHMflJ0a1TpxP9Q/KDnRqhW6DP1D90Ik2zR8pYbhuwnJoS6iSVD
sdAvmnN1ddrLoGkB4AliCwRm1DPKxhLQ2joh6a3qSUxeU0kSvfvWd0huLqoxyzd8hrDyHmEgSSrV
nLLXtC6oC6qW2pZjl0aKQejrvyqsJTFvBlcMtOkhovuTeIv26I3ntJZjjtJ96sEtyznIAN+YPa/7
Rb8bnoQf7eBCbDKAx7jGt3K3JqW/BwgqXNNQhlp+XO4F3JMQ8fcV5c1grzOiyA0gFTwFfvWnCuez
W1UGKrvmywm6bWmrxSgQzwKvbrTsqLPpHu0RYg4i1OdvtHrJ2sOljgub6w2Me0ZPszLARwxdoyFM
bRzhwXhxisULh6/VJ04zB+B7ayPqz6RBeZuvE615UXNkU/v8zbMhbQkZTTB8DJ1yknGQnOZpXQH/
gMg/8E8q8qh1bigNo94P4XmeOal4pK3eqIhw6TkPZ190Fvw4/UL8f8BksBt9PU7S/imaZlr/GagO
31fF4cm4Y520K9GL8p9UQ/ImHgcg8Jffo89RVLLxA2mA9eQrN8M0OCfC9Ht6yJ6nEG3D9wAgUluI
saCiDYUj3Ibz1wVkLYYcrtY1sA7+YiW4F6N2kc18XsQAb/RK9e3W/TJraJAL91yVf7i4ECr4Gkw9
kq+z4gN5RaPh2qPwPm97ok2nQ1oe0eQSPujaVPpGhUZKvGQhNXABOawDf7CvREFi9KnHxsXRtKJo
OpTVm3mvAaQ3Jrta3bcTJGTMOhgn2NTVpyqtZkth0swq9svP2ggOSD29iB7B9Gl3+VYkJSkwigPr
0TlOKrXKmqZMJf4DBMaCN1NR0d+/36d5u285PB2/kI895AEoTNJUtVBvsaANyTXsrs82glkQVGHG
k3srWGbTett2kDEUobYT3uSgnE5ZTaMSZSnbwSeOTCdu/aJ9rPsZsjKxOKzJ8TBCSICT5xSdjfYj
H9Zo2n8iiLQfn3C7gGEYmkSq/TF0KpmLhVl6Bq+zGwXyTPgntQ0+KNE5H0FsUWQmWZeR4nDdX1a5
gr6AudrT15QPbdVg36I6zq1j54DqMao4VfZnEsE6H6KS2LHXWNaVg2gYr7KWKheXhyFOviDsOQuH
ivx98l3RBbvQudYIASPLPrIXbXw9TOXxOHJU8z18Es2XdX1ThjSIU7wSkXF5h33n8Scy86LnvIxs
WVQ3NTP8doAabNDvrnw8cn+jJ3iW7ndwdJtUqG7DJyLZP9TclC0yTBeO9Xov9X4X3vjV4Geg5wC+
pr9ni8gfXmwsApxxKGsjvQMlSQnezh+QANzz3vW2vhh60J8w8DTIEA+yRmGnAEWSdwvChfxY5iLN
Yx1f2afqOXOQEshCPKxgb3bS7i0SJ1BW7iIb30URQtmCzg7FFypXxLuNpZBTm+3SsZPBfFNKeIYa
Iqs4cnqL6+CNawiPLJJQuwgViET+cYG+DFC0kHWY93HGrpECZ6eah0PHVo27hedExLvpLCuVqRci
hP61T2SZl97KpPpmJMJbiE9e+17VSP9srUI/BHZrcCkv+dTDRLpgLFuzGIV/rXzeix5KapsCOS9K
2ezuH1xZ2f/MwD+qjf28olax8v/sIEqp9VSIxBBBjU4Ou2M2FQe3KQ5TeofAdYyaXb6UdNtx1FcD
Ouc7Jo1rxn3JmTQrNC8/UDaVowGAy9Okh/kmr+gXm1uEccsJ3p+daNJ+Tty0j3a61ldNeN9bkUhX
ljeJTe8WnEp3N+ckiBluR8eYjm8eZJBJ619chtfxJvqZoegaBEgc1zYcG/6l1M39jU++Ari1gcsJ
X04BRcCs1qlFeHWskwq8kjXy4fTYQBcu23RkBEdFAqNVuMPVZHUcIxunlzxaHzh1I3qqclK7Ib9g
shKhXTom4n5BWqUPxDSFosruiOaA0aqy4BRalziyxCJ4cz9Ip4+V88M3S+mm6d/+iuwCJZuIKSE7
ij49cS7GfgGmJVXf/kD0MzXAHegkC8yW7mVzvAOTraoEsPZ+j0xjEwnht4s4n8A3toGSrpvc1n4Q
ka32fEr/ATxCgRHQ9Zb9rJTCFcX4LAnJFqOOlpIOQcIGmaLY5lHQmofsug9z3RlhF4l7NW/KiMZs
16gOyC2LFImja/o9EUxfJ/lNA87xwRP2t7IZSZedZXnSrJvYxJo//KVn9EScjaETvvoMUlGI5egb
F/kJCpHWelx4nPZ6oD307Gd+KcUreeMSLtG2w3Wqe0i4OVIY7DYxQMNrAeSRKks9n2xHXYgiSoTe
IdsnmJw8fT63f/R8YZJIF8MijdDxOHfbFBcHlSeY9QOwFLqegChYz7fs/xl5scLE7CdP8nZ1nyRP
29I/9L7cHKL2FI682fJABWSH/SghIg00bCVDAU7KMrsbAIJLT4uSysDXQ52k4mlBjUKbp5w/PmrS
k6HFMs2sPdlHgvVyXr0nxqzlvLM7P9YS/AqCCSwFkA4BBXKHCCddeuLIl2BlQ/HQkVktuwW7Nv4n
EPkhbfGjCs1vYJTccR29ogI1isMWBPonXzpjP/XUUXGlL8O6wGJJAbGPU/u1xApm2uaeF8IUsGHI
TuuHoqmcrfm5I4sce4JiM1dei7csPce093ec2c0Xikr+DerT2nv1EF1haIJOqf4jeB4uLoSAYo4s
7ZWTINjibKpNcsOWQ5CZ1tnWULwQvGoaQddtOh0Uy8M+E3bdnzMrUurpamPruZlFobKub+TzBTXr
k+exchn9i2dHl8CnHQ0At30fAbsYCnCTvdxWKX4w/HzD2E0ncKxvhg0F9Co76DgxIEA9/dXfWO5Z
9blGokzvFNSPUK0J32boxnRDUQF4jEJA9PYeHWrFuBku2Y2svwKezZovcaCWGUbtHBlOxHipQMEP
YWqN4c1s5pjnY36md8wTZayU27K2brCJ/rgdnsrIRaxHl4XhiqUpEPhxBEu8zdGQSWuLq0LQAyr+
f6Rjiu1rnWqbUz4unPNuGfG2WoL/gv6XGrqXt5erOgiV4lkysve/43+8Xo7RwRL9yvPfMEHpq5QF
67ry33hyu+s5RwS7J03NKil6RQXnxraLcMuOaMC+y0lq4urw9WiXeFMeSgLYt3smqj1dXtFQtWBW
WLpJ+DNopHhgJmpGbOHrNXKve48YI/6AtjQ+45ERCNdgJE9CQnJiSojewZMaM7HHeVA/8iU48KaA
GJ8uIe5KK5wVfFp6lOJRn7BmJIe1+lkt0du8rhzY2USgakhP3Dl7Xx3ED0PMR0f0tDvfBtRmoE9O
l1hEDDaq3dYlHqHBMJoSc5qoqZiJgiNjjwIzys/MA83w7quLX7UOztB3v9RTtUEwFScQwg2NsuOe
pCjMupWwciB7TOTiwyXL+P87ShyU5STqZCzDdXldhNJCEL3Tn3e8GuxCXUnsnhPb7nUmz1zjlw1M
rVuhpEgBe52IFT5AjIFpDaRifVTK+MXLvuQ3nserpmIuRO8dYcRMvAX+MopA0IBtmPuI1O3pBwfm
8+n6B0RRhsbPcLaIaZUgf8G6VYTbPebwbj42AVQu1CdgZixkVhcblFLMDit6MJOSORR/vsh2RhiA
b6yHIA5JNUt346Bwb+8SumYnDjl2QrlJdZoangq3ekTMVqq0qFCE6VVX06UmoAKo2/Ce3HBTa0H8
kABMZMHlm16Kik6JFr8rk/r+kwnR6cHYRepBg3sBxVtaadvg5mmxW7piMOob1b1BNEKki9QHRtS+
B9+SEDZxbZ9anvaAmkTSX4hUNXXpVVQPlNOBq8CTTQ3XZ9FzFL4LfaRp3x8x0NB2m1CuKSvSjd+h
W1Q/qtcGiR5eUrJFS6pWa5HRHAdhJ8hGZPu5gcrg1yWE+xhNlKWo4QU444ViWNjKeQvz/atJzdzF
N1kHevrgqCF8BJcO7VAXzFua18+/T0H0GuY1Uk8r/EetVoq8g1TCagdKLK06swRUGewuE8FG9FHh
kazfzfsn0g5zuPq+zRwGD5BbXaen81DX+aMej4tk2RtNcVhBY2MRytFrIaMizIkar0s9xakqbwkP
jr345hRDHuTi9jiFxLW+SeH1HhnSyISfbx9bQDoOSfVc4dT25Nyh4X3RFEru4M4VLLLrxMJ3xOby
Rmd/0xhrJYlzitIMTE1M383mT8sDP7mkTVvpaYL/ymDEeeEsfPsPWnBKJ6lIME7HZt2AcaK+ZMYa
IlFc3id2DLzp9DEw8KGUT18nhKmVqETJ/QSm9PM928lt3wFD4wwiYeLBjsdT3KYaxdHUfWoQfOf0
2MxOVNHJqeCXCeYne2t1H2lr+X0JC/FTOwHacixOqLyWslSWzhBfxI19WiuaDqjVG5JLJJIycBTy
pIXn26zmHRMtRxFuSZLayfX/JwFJi/OomFcrd4gUuGlpHcGEvmIfiP61u6m9jE2xp/it7FUaCzxa
WC94Gn9b7czSv50d7HLh6IbsKlXF1EPskxIpO4ywVJExrHC8LYXcOkW9c/4ojSgdIn3MVNJYkeU8
UwgR3JqwM5QZAa5Kcey2VyxXtEzRHKDB7oA1z3sCY/Mw1mU1F6N9M2emkHpokAvcMWs0TUUYcfy0
F3vhyGr5NfYrR5SQeXHlhbl6UoCqAwmRHb7bZtcJwTK//KHlQg565dMBUWibsyrPhd2IeGXdowNk
c/iPZKTrCz2fc4BiemKn+39Xv7CnjbHIfmHypGpwM+0kmRu8VJiz4pcaDFp0gzUt8SyxsaBM4ILf
pFtgTa2VSp1UGwFsdxVqv7THAUpKnUaOTyQPb4IKikIfe1FhEWRqewHuEIrAGG5rTepgVEk0wNCk
eJQl41bDg4lrcLdlaE6HXjP7nIko9w/GI94UI1DV3SzfNeIUnR0Yknj25mSUqKKejvdCszZ3q3nz
nvjD0b2On58qYTDPOSuDRKy9AUZgllJCX/w8foSFnp23OdEJhrq9iyiYK7+xnjpgOJR0JNXd2K7H
1x2XuxORKIgd+NDoqHwvLOAL1lDL/L93CoZ30ZpRdaoaYo/c6sH6sIIrKniM+E8PoU+tM3MOt1Gw
TJD9i5jvz+CpihNFYGC/ecfIQsBQQjGZ9F3PHs8Id5sviSPg0m/tKYew7dOiCppqjp7J5gs2KofH
MJnUDPJbRIU5Qzdn6h7BfIw1I7+wUlEbZTRsRgZlpVbWdEiPPNKAosneJYuheyf1BOcsYBR5PeKN
VuTygU+G0DEvZi/Vs6NhyZKnxzqZJhZtBzBjYUNSIBiefdEBAV/tQfqo3YF60syt3+wXXfTEj5tu
+4JNpm1hMOPaulrsYNUOuOjgsMivlge24wiybIVZNYK5/SRbGd5GMcZCoFZ16KrJUpl5PtKBaO5k
vnwKLKq4PLCIK7T1IOVmv+0tAQq2d3D7mCS2Nv7n/Pits+7ZQbRA2QGKqaJMYvSnKFVskWey/hOd
pydLoIEKQr8xLMzJoesbPIbUC4kZLZIKNeywMvqPRr8yZsdBRZ2K4Fdwlr84EinFvuQqwb8Acczk
U2FP/UTFjRscHdX+xGMeW1pogDxkjYrT+fn7YZQFn0dqSg+mB+vlnkSStf/H51MW8BFBhLKEXz0B
Ck66h8oxSPnyzejuXh7Worb7jJIS88lLbHtUKXv5ucl3vtXQLaZzg8PJKXcabvA68Z0qYPEIVRVb
nz98VWvkUBU/j1MEKumyi/bfU1Iu/VF9FaY1FXXKsq7+85e8+JPqiJ+hu/TFvv9ndXq59pyXvCMW
oGTu1gtsBzawJATBK7fulorpkm3/VSVdW7foAvALtJ1IppycM/sPceeDaYoGUQGsQlWIAQWM/4pS
E9gAW5DvksXPiw+JQ8h3wzCSpAZc+Zel+DU0mblsioNvfeJmFpKlBdfqNVJQVy1hCYA27zk7XhqY
D6dBPIFzIOeqsIiyDJdW102TmBvK3XbAp78Xl11EiyGwLWS9JF273yjaQmK5YvUOmSei++TC4S1z
dxRHJMjrcZwG37+5EqJIYJcwLB/pjJPjK0wXH3CECs8o02BrLLHXmuUagOaFuwKqlCgL0EodfCf6
YWwWxBuVpinPY8A2vrUNO06VajS7Hrn0WulAb4j7RPzDis533drS0msLtKIQL8wGqlpLnprRAVsy
vy8KTKH3WD9FZD30cOwZ7SCQhczMh0Mpz+xf/gRuWknfn5MfTOYTC7YwHHDjsm3TSe53XOJgB/wb
//VeaNe2ROvSSNii0ldwzqE82Ux9zhFK3lL8qzJ5AAAGCjRFP8jC9nibzh9BOIKlqGVDpdcRnHR2
tmfTh3yucV3UJR+03tctDrMyvuJX6PlR9Kn23f2L3yyVj7o1l1d0Rvcxkj/ZaFqb95O1wqqYTl/g
2T6rQX0w2KLD5+/QPrMMfWEugT4QrMzk/TTh1SlZQFpto7vQXE2pC+qgyNjES54iw0TQq3hvhVjD
42Ckh6ViMIvkn1XpIekJP3B4ftseNavnirDoLwTUdcbV53LROYNLmXsr/dwxKKJkcZNvfTTuvGZs
OxY+pF9ztVUFxOTo8EOGUDRjUf1hqPkmAL4vlBLZWDUvHSxPJsZtP9IcxYz41d7DjSfUZKhIswKs
4ifpRxYskvNfqWyv3Ll9rLCoy2H1ZPenlokWcL7ZNmSGbqq2xgLkg4O6SBeqVZ+AgfXkuUofPyEf
UVC4qhy+/0Xj/snATKj/t9n8cQRBT/B+Ke/UbjUMZxfjROF6nGH9bgUIRalXS400Y81hDI7V/4WE
Jebyib87Zh+8bC/I48fuF8p6AVsuO8SCv4ox05aIKITQ6bcKDXqDFokrY/a0K/4u8iZ6Kn/LFwoa
e4/a/O54VFBQQqn99DYsaFcRmE+kkHswutugkYDS4Kdxpr4LmI08OOSw44vOW2USyG3K7Ra/l6sh
ixTKu7seuNK0S09b3kMvoI0oFeHAEg3Wd3FpqscppW0LcoqtP9rtL5Y7buX2AyIJ+iYFIPMlK9yT
1yfAXAyeYayd3z3ZeeBAcenxnzakcTMqAnDTyjDogK+q/20McRBvLk8AYWz0lqKcUNMYSZYTqhfo
XIIGWnl7yPx2+5XFEkv6M9C2kQhgjBFb9e76RoSgpLHbA9D4juMKxMywJn6pK52oKtstY9EUYdzV
5Etfd46K+W4pJ5d9e4Mn+BLGCCVQ/m8+M+wUxd80ZUMyTLqwMIzWa15OztgTedXSpQEnkbicWIug
S95bPVTDJgD6CXgcWrOVw8ApbC8Tcn0CqD4OwtTLaV5xUH4jlslO9z043Rh07V8NnUS3E7f8zQfw
WYugmCYvUoQS9/otewpgPWR1p905zHTgPXcHbFEd9PIxZIYDWVtlkWGU5OHUqCs9z3qVIGGctHos
+h9Uk9ja9OY4sX1vLuza2JRLB3GwCMSLjH5GqDWLjv68+WYoMrrJu/4BCeAv1taAatq9NOLTmLiZ
j65McfsqRPai8+dFgBvuNUYAGh3Na3Y1Ivup1jWygeu9VoEfpLYLzNzKmNGUmkcmUXrzZBPW64zc
Pocox63d5o3WCJn5XsGtD5obb/9EAPvXDyAgoEOxOjdwM6toAsbugk63sqffHiH4rLzeZ9roj6z2
gw2Yu0cKw+YOQ8nBaHRZbhGTbNAsc87hxOJntJyYaeE2T1Jspt9dohHMyU4f9eZx4jstj0bgJrDK
24mKWRu0qx6sZ9ATO5DUoQQ3PLG88gj0VcNJcpijEAL+9x6clD+BEW4InvQsd1z5imBVGvcmRd3B
QgegI2UxurbJAYBrZS3Yv93Q7Kr84rsmcqeS/gBp0Nwiz/HPyHz0Wo60r9KG5HmUv058bPtBqFZP
+CfL24N9zX9tpYQJ78/STBmsl9EyNK+YE9JcLYdp8G4mCgul8l6hV1tG13er/8dUptKQ8S6K3Dx5
yqzfB34Ing42wqZypvf4YR3tO1fMdWpGtDXDC94YMtN7s7m9rSwg+NyGI6ePk2xfLwjSU5Y2u1f6
NoHuBpvNGUyo8snkhPiB7Go5WGu31lKlw0ILh5iEOLR+RZB4XTxSEWbcxFgpE6nv8Ihyo7xF22mF
4KgrOcObRDANiXfu5pBhJHRxvRfXcSCcGp+F25yoA3m/JTUMHWhPXaQ3LRLxw9cbzaVsTyAWf9Zd
unpv1DN2T1Y65exJG9QM9bxT8ymQfDWiJ1ur3CAKdyiFrLx0LQwQ646pmUOF0GcL05XNm0hWz2Hv
EBxy2O5RoEkVs9ULkTfvQPfr4dZ9ZVePHBYFlBPqX8hECRyg4tKcIpHDK86k+lDISajNG4oxdfeW
Wto+3GOQ7sfdXESlKnKc/oCFIXOeu2aCE3jn2AwJsVRrZdbM72yI7MODzGlkQD41d4gqCM/WCvJN
qmn1b1TgCfGJ5AW3K5M5aRJO8+1ERD7mi6sn/PxYDa5TvMAcwzRiRHwaStE+IMtHMsoovJ5AqqzQ
aqnVmz32t2fNt1sSatpEm8ono2zWqrMGOzFV/AXG8TlgGRK9uqKoglYPUt5oyxUi+3BsLYdCA5Pr
faHmdiAxjyfQZD0A9HnO4zNQ0sDY2bhCRVKMWXmsMUi6JBctvTZypr+yeu8YEfSOjfb5yz9EYXQ8
CMZTs6YvslHLpIco0aAVqgRferzohN6TebdyzEFR0ECqKJjmpVz0Geev0QECSmBCeuKEeXOvlRgU
ufJHtaBg22Ix6br7Eu2W+Wv4couxs4GbwOFEcVor/y5NSVQpn05JeLvxJ21c7SLOMlqjmEQI3UhZ
imOZ37YRTuIOjsnrbnS6m401NI/kEJwnZb9ZeqX9Uu7oTHmMGqrrxw+Y2b8PxG7YbxkQER1pK8d+
bzyb4JZFQCyLE7SSFB8Qt/RtKbSF25samWts1xZIue0rj1/PqHZgbzme/5nA9vSArue/b3yvbgcz
3dXU2s6VzynaHBTdhX9rlo/nH+UKHcEKcLxYjwFZxnc6SGBvf94W4kYddeohN7aTn+n5eSaVefJs
Q6gjBN7tak4lN5orEEqumn3cfeDPcmmLbAF1/UDLU8Z4AfiodPCUSYy1h3aq2XS9GmxIPGiM3aj9
6evwIaTXGS31DbdTj6i1peiUSb2JJzJRzuzciOM/rTPvEWIw3bGkn4HeHCIAXhrMvQw8IBp65Vuv
eh3zdPTbC0sEOuGalRrulgVV42hZLQxlH+tMgXvFcnrkLL35aKyqmXyvlKVhxxM2M3uA3mD0DZmX
1tyO95mCxU0RnIHpFLdbfoP3ufldgxkQ7vh7uKplQZ6WrED/+QkTUsxHIRIDCG8wjgZ6pjjQUr1k
wfHfN+yVwXvOBhpC4RlOSMOSXarbXqHVBB6M0+9hL0x4OoTAqgmtRqtnOmAhmZTEZMh5Qpp043e6
mddeU6mXiNN3k+DUbC+m7CmeuGoL8vjiJi5DGoh4R67HF+rvy6AwJIiOtVKwv6PhVrCf1t/jEcgv
hq+tfNfH2wwtaB9ZPa4y202Iw46LrA6fuLQx25RR8DOT/axy+wV4WvWXTzmdffbtFxLHh7Q+t1BP
cJCcyBBHa1hmv/ksf35sN6Joi7vnwc7CK81OLaLIEHzFg4jBlNYVRqNIupc6YXSZNdzHK4LaG1mI
lmeV954NhOv3pOMmL3wqLsBjIcDwx7fgokGa0EqnFIBwL9KXXoLVWSUALjX3YAFjYJGJh15EiENX
Bd0iuXN8q5vJHq1gtx9j9a7fLwUKXdsC7CtswgBcvofHiwRLPXQHkCHjcDvQbhF5zljInGGOkIee
9gDDvdtMFrdQIhfTnsOQlAEj83Dups0O8y6lSnafoIEIxKH0pspv0+xzCDSyWGfRNKJJOFzvFaop
nagLoceSDT13U1zIfoUBRlCctDZkp+Xu9fc/x/4+n99IzK6dOifzesiCcLaZ3zt2o7oh/nxvzb3d
vB5xJoGWIN1BJZsu6MtrGkyjELev4tvCA6Wf5cLF1+ayDJmg8pkrccY981vMO8ZWO7X7Vt8Mr+f2
It2FnZKGdbL1ROQVLTiU/eMwzpV5SgK0l4YiD/C2AEgcGRwW0saWRaIDJDzXPFj59yQu6BAevipQ
idktKcTjLe/lSnYzoKx0A3iJqy1YBtkBXzn3ISxwVo2c9x0V3kuhYlfC5VeY7PetoQFbniqF9x7z
vagVGpWHycnP3AkqX9yKjOn8Hu9Kqpx8pw4XMy/DM2AowmCIfLwsfgvB+e11l13whC5CHEqBD9R3
xqWkkjd0sP6s7ZSMAa4G82cqVFl9966kG5uykN2rZfgi2uz9BZRpMnZ0tT2vp/bIDf3yCeB/R0QU
YABf8wpYK+7JKdQVSmHz0OK64gSjR8DHU2kSdBdg6NDiu5iIPiWhTh9QgwyCJ8At4DR9gsp9rgq6
G7FSkSmVGrtMrDsW6otyBFBbvZhrsISCk0hZn5xwtJAG0oPId6uMwHCOfV49DjWGyOhphNyPrQ9g
x9UweUkqkpUO6pMt56z/XpkLk7knn6ld8JU6obvBCgTSdSB685cTxBmJ7bW2JmaDoUS3K1JPl6n2
0ROUEL8NexQ88mujchF1x9EMmUttF+YLZL4weuZsiOc8UjWxXGhg7BmXRu4zyBXE8hs7/HGSd2Kd
PRexem1wobjoPsBoelSfma5Ly4pg5vQDjnmBgCKxSgpHOG8YN7mnpTdiPac5+zupfRqirTedYgYg
1VT/ZA5AxFyqfYk/C99syRyuSqbkxGwyneTQkPyW+pp0Ov0678d/pGL3pkugiurfO7w1NAX/bdcs
rd40yZcmuG9/tY+sdJUcXH5Daq8PCzaymeaQmK5goGFSxueJc37IUT/MO09Y0DB1hoSLoy4XAIeZ
IhF79AuojmKm/vAeoRnGuuGLSqu/1nCdpLfT5FhivKeVx1SqT1F7/0kyhQNfwRUT/KFTpPXyGmky
6BrAD+hSTX9HQqkIB31sgv/dVFWqnxlxrjShM7XLP5TkRs7jwoZ9MawU8bDBLF0hfbixLN/yvAVZ
9Juy6G3Po7mhbqsCKV7DqoXsIwKaaIy3YD8YHo3ODVc+nYd2+EamShfxi6JJtjqAunUz1WYCDMWE
zchAl1wCydKV+HkzkDhL7t3obbThhLAQXbMQwO69OB1WG9+LdKydFQaTTH4Wn48BhirUy6UCennW
pY5XcgkY3YIF8U084j4eCNybJyUxNeoCNuGghtg1HAFR2J0AUo0QLLXDdzibjaEd7vTat5wZDmIN
uxALF3ChgBMMfFx0sOgJUgBqGKfNO1ZODpMzhbQyXNj7gb8u9q31PME3R6edq2O7sr6D5yyh84vu
06S9n7BYwWuS2v1jZLXx6YH8zDch4A5lao4INvc8brv7jMKLbJoyb29iSrT4VByO8ZLX56mQXxuO
KQCQYCD2zoX7sUoiMDD/9b8nUgg4RNALcV4z4hK/rOXefVjFCYAj2xHS48tRbNsQHQeu97EbifBJ
mogXC4A5fBURYdzz89Tw2pTrLgr+Yrjnb7JIIXBgBuP9U/5/s190Q1KDHGx6CUt4BNa1kiTyir27
hP9cGrbVbfG53IGLzB969MgaLZOBe8n2LKmdKk3bXJS4udGn0tgbqLHA7wbQjauQK25DBRrq5gCy
FYYycGFrNr92t7ZEs2x61xCchKIcHrrWPZMPOfWUl5IA0LMHGDwh3bhHzLA64fxtiOIfEVphM+yE
mYylZJqyY5lpSIQl4TThu9lw1Zn1xB79qlBfxt/M7sGyn9M+31ODNev+xG2h+KR4+lHcNgH7qBYu
Hv2/4S/1c124vwLySvopcUrbyKkMqbLD8wFFYRqDFSRqBvU9lwiOujc2Sx/DujFLjRymNy/KTZ1i
/gK6K9jLMTku0TfKJYeEDVbXlqvTzQPQgYwYmY1Af9pzTeoDdA2bKenGEgsgB9U3jxqCkpk5XHjs
bJzQrA1cNxBQqMKq2ksRCHqCEumQw7176xXuQS1cVePfLQ/Ayj+RC6/UlN3BH8LLauGQCQy0HOT/
9kiFwBZWnHuXCKXgrBulywqWPVD2yVoSjrbIbvuzjhj0WSKNRVlnyuCmwq3r1oXpyT8P5KnFqPjQ
vIMBFFGbHJaZivrSYAR7ehltdo3sZPA8+rZq3ioAaPBnxLYcHiyFzk6wga2woZJRdwq7PTNRBMO3
4I/xiAH5zuDhhOY1NitaB+3fl0kobCwGmbMr+9XTNaXZXwd5L0sLLomniVj2Ovss1x80zOH9PvmL
dU0ZdV3lh47Oo4GOcI4TSb7Di0Ds3svG4ts8ieg6fxnEa7DbKudmzWfbYybULj5//l4H/d0wWk1c
bgnP87r/72cSCQMr5Wn4411rNdt3eXZEC8GwHlBLTKV9u2NPQIQ5KSSRy0UgkozSJaMOtPrXnMJr
ArhHb49uKkFR6RqYWNN/k3D1Er85r2NDPKi6mbd948OEW3E9uHm3rrDuSPHi1KkGFz1p/snN20c2
UuEZr56s7/DWHGZA3f7M1RZl+l/RDqv69tAjuVoutQZ3h4e/T81A1dAnE5ojmC+wCRflRvjxe0i9
NvyC3G/hvPdTo/lDIDeR9jeu4IvrKQuO2YkyNYCkQ+UyFNJgDSit6Qz+X1bwoMQmwmbACOH5CGmN
SRVTAckAtBc5LC3DGOdhLSnW2BmUaSlHqJyRreMZnc1WlgFtXeu/Qad+Hwvvw/ThU608vgtxW/gv
3+klT5bMtOa8FN4kBRt/nAJGEsFOMWP8d4j6++GB4I2Qzf+hYpozlTzbdqmVAlBgigw1QsyExTjB
KHJtX72FZFsIQrs+XvlgNP8CYDohNzflvtXq7O5JzV9WiXgsW6ZaqbPHa1InVez8Ck4FIOnIjtLE
GXuKFTQj/Bb0Aynq/yXCDNtkzjAdez8G54oLjEjRnaTk9q3SuN9E5LAyg0WQSAbL8ZKMQpY3lUE2
yOvjUWshdYYvqp9qka9hNSk++uzzTWYI7sHsq1J6NcKx97HeBiwseVBqPYMBQjICxkBa0d9FkZZe
uBoYOaozTMaDdOBFIrig6uhFofgTe9A1Luhp+MBttKm+o6RpSBsHTOk1g7HGasILTgUWPg2KYtjI
2xZEgoHCBnhDVcqlD6HOOQS1tnChBXO+qh05K2EF7Lc9xm9dd7soqQ/YKPs+6KFHi1vLttpe/4gu
Z032LSs/TBmWOb8hDRepv7828SL0NOI1aN0F9OlBsr7A3RU5WyKq1BNCGiOL73pJhd1GqYtearCh
n5Sy7Db1ZcCVEV9cxKRgBmuHXepmmFsdDXo4O1dv27P/PjT9jbCnPz339xTh3MKVpf/iKv1l5dGn
fbDJj53wiuJFW3HgQGw6eOpVqHpFjC3rxwtcgOsZiXQjEfIATGcl7DZlVHqcPi9udGdgoS/MzHCM
wTBg18EOmZlEEDqroNFjUe6NPiBRA1G5gRuq7xcQZhiIa4Sss21dPb3Iow0u83gKJROwXSDy79sk
ZrF5fDGiKt0JNKzoGOHKZxbAzWXs/mHeHdYd0uQxJLjA8T61UZBEJH6vnoJzchDXnd5w4n/538t1
6+TjKHaVm85OMkxTYznFuSZY+bDlZOvMkbdySGR20U6yXHcYV3tfjGHYOfpaGt7+mp2BTc4D8Urq
1bccLvhgfPM0Tlr+k/7mmcEalYy9HmPZkPkwr3OfgxAi8yUFdjdSYU5qGCOtPTY1NP2ujAk7hbFr
IAU/Qd8B83MeBWjrm5y+LPP52nFe4SaTVnfNMfQAbiyug9t1ckm5eM8N+iHeZHQMrJ7TKQWRykqY
FdmDGE313GmjbZnvJ2Ocza+d2fC5YtNUuJ+QTVYynXJmKsNy30xF4ekMFuSFFocNUjXAy9SFG06u
40ai/sdZoWGYOqsDm0rElWXyjk+lQ4W0n2mF1OzuluSI3YyQ68iowOnmIGqL90CbuD6XY+iWSSEJ
yK5UmfITLMTN6CdgSrXzIGuQBF07/WVt9MMv+A/Afvjq1K+GOMRL9dxNWY6lifqpAAKPqUa8yzM2
OiVnq/OtGuSta/9E43AO8ljEexEMl7quncB7fSEa7glQZ25wtoGg6g47f0msxT//IAxjE2JdDx6o
Ova2RVAlYWkoxauKfwvryQ7fI/4a+SdZSMrnkZ2QRM5OYPk4bA03XlqwZSztMDyikPt+OTOWce6X
Ha0Fv1P9U01UCf7E/rxc/Fr6HWsFxttQ6T+h4C5byO6nc4ZsiykcXosuqGRG9gC1JT+3d7KjdF7L
1eitEPTioWQx4/5O0XXqaaEopXQHd43Ot3NR6maDIv6DWeu7oEbIBpZAKf90e1IURI4+mzkUpdXh
XgOfHrxx2Kp40lEfLbfH2d3G0h0Ih4rwRMkqdP0pdhgA0KTi1IWvArE1M/PEsAJqK6U53yFb1b/8
bKy9lTr6kbSHgC2psq8WBd5cCnQ/ws6O+4Wt2IL7Qcf1HsA4uDWYvpGXD2YfAlFSQ3RSdMq84VUh
03QWDUCYpTKxYhPVSjmP6Ub4ocmUGH31MldjOoTo++4CdUV18x+XpfL9B4vLrt1XrQQr58+ZVE6g
r2hVUP63QUOukbz3SDJBP7FOWtGOI/R5fsOtj1Z9WHRJ7P9D2r+yEyBpOf7qU3mP4KR2RJ/Xwoiq
5g7VtBT2btfTUidtZuGS6E8CsVjCrXGxSHsX5d1L2A0vaXNUtImEz9O0axzZFixdNiGKFceFe7ty
r7xNbK3lOZfLSoZ2/+jY9b3J3sEgxoR5zzv8PliEMKLWx6YDvN2ly5d0wgrAU+X9vfEaiRHlbRmQ
lTbedx5Sl5utqjBQ5uoeXRX3GHbEZNCcvK3S5RFrl86ZW++FMJZ/acbI2kaH10s5v3xAxpen5vfD
gAV4TeZSGW5L4o6zi9Lm8eHSWTb7OxQ4cimeFVz7sFvLx1j70xY5RhKjLGSUNHBoDTX218DxDB8A
GbNSqYrmWUotNNrSq7g5rzZSDjoy/zBSMxC3xgQx8RpE1PA0ON7Gqk84oK08VbhjObuCkbfcQn0+
bEQETqJgA0TewjKFBD3Pl68ZiGjcfIxF8NMZX88+J1LYVlEyOCwhafHpBJZsQeCZZtrxQlbBLilD
H3HM3PkNC7YEfMRyszCxXn6W1VlQ3aOKe7G9/cGL+lDIh7dZArIakDeRKl99/DSkvuOFzOJKU9mY
buv9RRU2Cg3Pc8mEUp0T4/RXH+WaYEqyYnjUjqNY88litPoKgcrzVaZNMPN+GyCDvwzikRRranSc
O+TTBtUwVzcHRzrIsRgD0q+85bYovJsO1MnpFFS7gaP3agVfQkHQm4x9my5cgXLV/dQQCRuOrE//
IgR1WjKrmeZ/00s+jgYoJhZHK9CjEMwrU+BwpqbHXY/gW0GWqxBLwleebQa4jNW3uzEx9dNQbKZZ
7iSkhKt9T99KdQBB55WTku/PhLhKiIdE+A9YF3WaTckap06+mrLD9nG3V8FbvIW/It2n4T6QqBTi
qGnrGZcu/BnZxjQHCop6eMrPeWRCene+dXyJPqWGOqL4ZxzVasTJ23DbQhlolRM+YXB4PGJPstdh
Eb/KRYxcPV/bGyy/lfmNYUqNDk25mbPoH4O9Yi13k6MLHZKayliV8vwhpZuU7LHR9ZT99Hp3EO+o
5SjNtLHpcP7skaDSMYY8fUn4G6XooYZLwiJepBzcf8gU02rtgeWT+6F13xmkrPPy9IwekbX/tmzW
Fo60f0bYXcI3+7GI2Xi3nYTmNMeC7tA1Rs7MabK4wMOqgDktJexLhrybNq3Wy/r59fkkaXC46m8k
35IW4RO6oJSG3rB7m9ZJZE17xFfz5XbdTAeJN1wk7IuQjojEEcePtVzEmdRPweL44HOiXHaxxqlz
+KOVFkpYPWTSf/lKPiNx8OX0mk+QGX/Tc+q+xpa3kZ5k0B7lGld5xntGfccXHMT7P4JfTYWVvhgQ
gjM3UFKaCoKu+rwOSzgoPLHbDPM89mEVNOhD+H03++jj32DLvGzN2+B8eHM0Duuwvwr0Q7KboImk
AOZqZHIUTOpeIuv3VAFiIGMRfGZk8Cko5jJXcQua4KrK4L2w105ej1HvN94Rito5YDJ7qcYH4jCr
WGjbgn2vkvCnjL0o30WokkdBREnLCa/x61sRM+DHjD3RRHC5bBVb+GtDRy/9jWfGzEJQllTsjvMR
q96q5cxWClZeDN5QH4N9Y2u6aIfcN5fTei4+Z6WG8cP05xWbdQApstTtgY2RTAmQw6EFHzyhxvFY
IaCmhsbpwm6IkTVIS4k6LTfEgWkjtSNrQFa/wjAJhP6riwcOKXheJ6EVQUntMW9jYSFNnKPG+xdT
CPl7V6Y418gpwQIlk2oNfuMeBngSns9vQno8jCykZRNHlFzRjhdVBDOTskM8cVPjjneFO4J5SOms
PHAvTRBDe00cD7Dxw3z8SRYnG8iBIDsjLmpxsJBUUE2HuLnXRDB4RlFjC7Ak9fY32X/fso+6+S3k
TQ6xqaAoTbah3XIyKF14qnWFNDNIqsFf/wrj2Nn80A0+wvNxTg3PJ9V/DgahjGZc0OEhjB0aB6t4
CNY3KL/Ru0tQfztD6Ugi9JqkxryG5OflmlL/LOMS075SYL4q0r5Qdd+mBBT85dPsLmtmHnfdDolQ
mkf49GAeh+o1JBEvVhy0jGr9XlYTcbWglkU9VJxlZtK/4QTVDwqDnPcFli13JtjhhJox7zji7nYL
EO6gqjz2B5VlJaS/UtjMX8TCRPUwVIhKjZNYCzcmUqOvv+2AI0Mb5gCZSaYBye5BP0pcdw0+/8q/
q33DnEmZQazGYJsZuCVi36UHmO8CyHuHU06NftKuOPOxEPEmWU2Is5z19X/4NgKfoQYRcr5xfi77
qWa7FQaXPO7JzPLCGZAPR1fUDo7XbzwsUV4gyNk3r2MDdmjZmc84qq8fgeLs7X9pdZrT5EKnK0/X
4ozQDYRxs6pmggzYWL5oQenK7weqkV2aqxHCVtGrgPgRzwDphr8jiCAZVqFIKZx/9kJXroHe5iZp
0FK0bvtUNJo9TYi2itQ8/CidgaXer8Z7nFan/a+zw4JY6/ErQu1Y0PMZSrX4dDXil1A+j5Fa/kRh
peHE7H6JPh546zvMiRNgPufpHMIzlO0Gvf9qDKbf5sf8Rt8qDyUP6HRIFzRB3VxssVqrM8FRI2r2
Zfl5DmyiSVmHbJJIUDTrNq2WR/RfE1F+m3ctM+qw1Bfl0Q62dt9kZqt3aum2xxDxnvHza++UKyzA
/itx0D/ZmxHA+9CKpQ+R7IfJiCDE3hKauALMb/ILcvii0NmA1hwtYTxyoxxW3qyFReUkW1STDQpl
kDhdqhNrLR6uysRbVz5n3TOVHVEGSFv9OxGsMvcNT2pdw0imdwPyAr6sCKY8ePnGpjdwzhk9zQPm
STKiahw++MFpglJj+rcGLuT11jmKlU4wmEZ4UKEZb+zBaCkkW/g2d5ujVqGqEwzacCduicy61auY
TlGHZa0omBHR7BBsMJlD+0YQDSASPd8fpKp3pgL2ntDCf1z6lVs/Oc9vH/E4lQD6y5/TdMaojK/k
XEEb5vBN9SQ1tpQeK/k0vbyEAiSm7C+BqxcegSjH6K6iPwZCiuJQVEwEhk1eywq13RT3zesxZbw0
79ix5irMdOzndW4cAwIi3NiI7qSvi/UPK8j+9hHjSHskwJIBJuRlAzEp3kuhksyR0PrUGoll+SZQ
BrTLDLZZc2+aAgHB0JJ3ZlOJmffO7WSQztjlRlkWRZ8iI2dV5GsI31fSjSf6tz4yxMlyicahOBhb
mM/L2gu5JCFbf9p4tiUkgtgfjXc4MFo81x1r3hLqnGj4PFVQxX1ufuWMDiVrPNujl5eqPWVioVsW
mjNCxO972U2Bcx2jVmeroTk6VyiiRCfO4vnES38jge4nGzSr5IehKCUpwkPNNHuOfozzGQVfoBxn
EAyTWGCpZHiMscJx5fW1gdViOOCeWwkrtxO7LVihf69MYpm0VwygocEOjrvrRdqGuNRc0G3wf92O
mxgDcqFNZInWlsEj5EwKHW8y3DKCAi7aoKoD+Vz5YwfXqZHWYydYzMUTdOTy+ppRGnCyRqvabmMB
7+oonunmYTLizzjSPCD+SJ3z+Dko1sbiTWhrZvBB3y6CsyEH/NGrNQNeJDVahpPH/cfX5uNlMHnd
4oX39aTTS5Wpv3vVgr1gvU7iDlTXDzdD44g2NyfSgtm9OUhRcDab2GjfXQiKA24ebgUcmhvepYst
LbakciNqtaKgw27QtPpPnyJppC8/Zbu0hjqGdHfapnUu09p1+/yeY80fxbrNQbrJXinGnQu5VYvl
zETMc79TQdzOrrD9D3C0xWt5fsCzemniozegnPpL2X6PyK6/SXmqWWaq3Wa3XJRNMI5+ZcYZpO1O
FVP0PWoppi7hnpibh8fhAY6uVk6ixpv6IDDN70+XYg80HO082oJEsIbuAHv+YE4U3XodIICbAyR/
el3W0QjLAriOjyf6z96M//L4wag0+iTrWS162SW1u8CAbiqI6wqrz24KgB0yfCZ+0mex8aMCaCDN
cn0uSSIvUS6D7hDXZEln6QGDn0F7doRRuBAz1OXvPrHvFAzgrOkV59PSYdF9chCTU/J2rxl02dCa
qJNcHtXWj8U3hEuzhoiXPKXKK5g51hMNPwS6H0OHlgkoD8wNykDGUmlRJE3mHJeMbzs8Vw+Ibr37
Wt9PsjUmhspvLRn/a8RAxaqi8vGM84Fn4hkP5rQZvuF3cTriE/m3I3ZoEeP1S1vvfNq4rYncITq8
B0O1GY6Lf/UbbDy1NvZrMs3hb496aRDKNT3eZ+8lECn8n+5D+Ue0OJg3hn+7/fjUMw50j6CI68wy
IvHSw1lX/Knirr35hmpk2x4pRFmtjVXlYlo2CeB3bQmZCEnw07mEH9XfEAyXu+2bJmKvYKObgVam
dtdVfBDenmCGzRy8Bm4uag7bqnQC106cNRka/AtHprxOh0fMmDwUHl/LTzSLlNIz7tlh5YP7AwLm
i01zWZFivc8xLaMNqmvqSQNkXgzs7PUNupU9WtjLLJcelEkal0tIX8GSnyj1nFUQc02rLikik/ip
/pwi+B7wmwAVQo5FRT/395QjAoAuA6qYb8KK+46vYmlnpuA+CNMRtpF7PA77ooEoaeojL5RLZpYA
ud+ReBNBmw2aMZ1vcjaaW3t/ZY2F0N4uzZI+KGfYj+w9+54B98K86hgKg0fwPkQjKMd1J771lNhb
jTlTTc9xf80Yc2+m3N/2MZMNxPDEhPXhUBmuMCKzAGKfl0o7B24XCb26mTRs9oWNFscowED5hP2y
q9+oh4jRkK8Z8KfqU8zOYMIqfmMa0UzMMEXWqa4c/zLfpBO2JXA0/7STMkEkoPJuZAKf7nETZfvI
1I5WZ1Alii0ppza5hXUl42uhT9aZxCI06XTXsLwQ16fBUa3Uv/6J8KlaS+dy4IbNvsMoGNOIIW/G
PPlbA9+k3sj0LzEwbzTTbw+zRIbdGz0DDvwsZxyE9y4wxJYVBjIGSsVtm8s4i+qwJbjD9cCvMcy/
8QSbFiwFNoWslwgVssd5+iDPjG3GR5GPnUY6ftPX1wDjFKRllClzhrL95GNfZWn80GOHgv9L6e2r
NirMWoAe5G5DBAC10XCDVaYCpJNkNfmfGDvOPo+3fH10w6VV/U2FVscUpWl+eO6ky4OYrGG34i6V
pC6VQcKwzZTzaMybJ0h1P4EMTFfZaXybMZGNCmoSUoIdbUlHlzvnNTtCFk8kUbQ2bmDNNbzDpuH/
CaVfhbDcZ/FRGZzfDAm/4DAYnGlsrLfA2RKao5tHqkoFFfq4bAzjiPCPXMfsbIBD9wDYFBcynn2r
pCuKCspRe9AnXAAe1HH4qNxD2eOV92lxDCnhotQcIQQSA7BgC8PSv7AcL9Lq2q1lR2pJVR6L/+X7
mq4T2/V2q8yx9cqe8raGy14UNzFDa0ls0CYkPA0vyT0aiT7328Jc83sYP4snGKa/LrBmn5DpDrTz
2defEto6AeECr6y8WJJWOE5gX7KGFOmmv79vMR3CoAU3momjW+AyUMdLag/E9XWpZfsVzSdyoFQf
IBNcmjrYo0CxWh04KkS7VJ7TYZsz0Ul2Glk1+KvKW7Cm2YTA9WFKsCo/ZSn11wZMPybgbWM2AX5C
tOiynA5gUCqb5IWaPTjYBK4GYyuc/Yqdee46odfUUIzDaknZfCdLFr3T3BWyTB+Me/LVmzy5/YsA
iQYaQCazncj3TUlQDfpLScDXMPtN80axyBvao7D963vvzEjJR6J2vERAINMDdfRwxUTuuYLUtflp
Nz/Hdtc9UCc+iUthE7TWgV7sqEA8ril0p8kLfeD4ZtJa66JR0dU1CX0bWmdTAHvqPwGX2cczdHq3
Squo2sT/Typ9wjx3+O5lC23gdu/uLvnxj5frUb49MAyNNhw7G3clkur6uiNiG3P7jLgt7gM4XsHB
16VkoBjViOXWqi+Df7agaolWwoSQtlzrTHEH6S9pmP3S6oU8Wk0YnovsOl534BdHc5rBuK/828Tt
4tgxikxDSqaZUlmnGK7hictwf2sZOLoHWnJvHq7KREyrqaYRgq7dM0xjJTHTU24hM24ih5hHlAO3
5eZYK7/qn4tvf5zLjC0k5hf/ew2LlzXuXniDYsLNiSEXi6Y01dZr2hEMbcZ5FxSX8DUusX2fGCCx
oGU8R+6OscNCLtW442GJ6BdXHDXOe31/H3QiiwkI49VOmZ3A7LQo0MVL0m+mUHvltDeXu+1OSUdw
1kkGKduZ2sDBdceqG/iUA8Z3Ek6YYx10sTYWyyOywh8wZ61DAy1OC07J0Oelsax54KCq9AiSw6H2
ivraX1XZux1ec3CyCskKqWu95hCTpC0lIiaVU4RpdhfTtMWlP750WSklhKcge0BNJ+qPycRsPKI7
1WGlrFZSZsX0TeaMAXWkx0jtHntyr+tl5BUOyz3VImEoetv35z9hcQGdOT7TbtJLP7q5kPM7znMu
w4MHvlpxqAOqXfORUm2cXFamig06FEZRwlnvYt781zbW9FF1OWhTmROvYNjuadzvgSTs0VXMpyBE
QG5HqG5NXMIDpod+wx5GVvUpWEWkjgKIDEN4Zm541+ibBDrOFoLeHedvx/rpR8Dq/VoLSOe6vKMN
ssDFEoEyHBIsju2y1fRwDjAcuneUTIK/AkFDheZktXaDL5w2dGx1Wjwa/nyy6xUkRiUjKJRVmH66
0lMj/MqsWoavoAgR8JrA/Hfjknn3iQsJFkwascS+t7A9GvV3/U8asnlE2dGdgyYPBlYvoltJvsCA
zuXMdrfm9BjoIAobHtENzrurbYLbOC0df1PyV5/b+7djdYUjYrN/jdniGrzCfbsgik28XkeRlYn6
Tvo8drROlt+i+G/utQlNSvGyilLhh23XqqHqOSL7Rthh013HCXU3rYcWVqe+Hsz0Wc4pWxfuZkuA
tWAQfcDqRZG027O2MCuphivHTe+ZKx/E/SS3DLbdYp2oFvXFhrjIgHDi5iZkxSh2sULItgZFTc0l
Zy21B/faUPWAa8rySm25LGo2zoEKQRxbR2H7ssvivVHvt8lSSp+K514p0AEr2WaGd9JFgirgZSB4
EcQYnifu0ozqJaf8PygAgYAGgkmLePba4lQFuFBTBhM3wcsAggWsUTfizqsFiop0mKySxhxgVK+0
S4Nt9kw4l35GdYCK/wqJZ+8DMfcvhLItUycmwWVwCHQVsYF6uaou/4vsLKJtyJKmfRSuv0ga1VNT
LQcakR0s/ydD6aUVmb/v9ytm3SJ/8PUEMsQJ0f//73Ax3DjzQStekBtiJvgbJGk7BqTlbfkngF/n
g8/62aGvE/5V1MKu70WqWaUAtOK5go1GXj2fnUctYybTVEMtQzRS115P8YADR7BLv/ZRdpQdZGu0
OnZ0YY4Qbl9afcRqWgkZsPBWi4uDyfZqnSwjcNCpngAbyiFDk+yvn0/Ye4RaDy9WuVNF88o0ofaX
oPQGmBhAiZTC8w/ohStHoRyqOv0whGKQ6DtUfrLi+7vK3OSdlDF5xdvU+MiUnlfdItzd4nOXNCSe
DQs2x/PKp0dO/cnw3v2l35FZ0c5L/jPo/apbJcTct1ee17emvW1NJG7ylF+4hNtPxOoaYZUMmnYv
tWUmwKk0UyA2duZU6+TmazEjDglKe+7pG84JAH5U3yZomMKRYfz3viom03gsd4cmPu/BZ3H3z0np
DJRa1xVxN68OCOf7sCURl/BU8neQzoQ8oQ7VZoEZWrGb6odn3PaBYE2syvgR5rW2DaCP74qQNjKF
Hn470FGBbG7/s2YTjrWF/Bbv+2wEjHv5ynCkjJJhECP0O/HSlPyh72SIAg2+CE0o9TqtVhyqvAhN
aRcvyEMQsRhap3/kUzTZvzJGJq2fAbucBuQwYdSfrkB/4/S0OJzqALk0OiuNPNtPKaO5tg4IeHhn
UDDrAWrpQN37rLUkq6iGDdJzosEU5pXRm8vRla9Zw5i7p9Us99wPH74xzWvhA5vhv673OgH6Aga4
ePz0jTnL5YGsQMlPetpr/JtVcEI5vZN5k7E+abpoyXCQpYOtMlEdb+PbdJ0yudjYqUdHLs1wD2ZN
+gy4qnzVeNCRmKGQbMWC2LP0CRGHvE1cVO8mTGc0bZN8QGpnNNVVDB/RbOkA6nF7ElyKBXdz5sOY
1pLoDrkWI8bQJVm520JafK4zq3xSluvdZdpWS6Z2eq+RtYQz66yGIcA9rhOYgcvunyZqsU3ze/nB
iSOtKce7ZhZPkwq9cMmLrof6NIP7SiG6Xw9X2vRUzMvcKsNAr9A7mLlLu/dwfyjZJjzbe9rhXVXP
Da2PxOyVQdjsnDnc6LV0mABHVz5WYCxT/B5yiikwOt1SLLm3U+1jX9GpMaq2M2aIc0Jr8x5lShA6
Fff3cbHlmL4Nu8YGZU0AMA40fxspScQthQsoQVp9mlIMV/ZJqxcI+TCySbr8pTn5TuHIW/QRQVED
8g6Yn9gMsLcv/xR5b/SwNCB5mCxMnmoYW9yyTOTi0h7dDkmGjK7sHG6B3xRxDtEMyyUdTxKskKiN
wejUkhq/SMp3AH7zM/4jgW5j4dEbMlAIhbtWRsq9uZb6rUiZcUHqeFLffoXKMSvoaZ163x0EcLTb
mDTcjyeBCp3GwuqixIdWoEVCMzIMlHu+wC9BbCMHmGE/xBupBMZunyPfnmYo6HfU0xfXXdKYr9Ih
VI4b7fO9TwOOvdoYADgZ13kxBNCjnSc8UDdOHP9kfJf5pllPb1T2ZVE09lF7AwSmj3at4WBZ/DfY
suXbQMiZ3EZDyukFeclC9Wm9bpirdpEl4ShEAYffI6jFKZkhYz1R+SaxDwvhz6qSz2BR7I+MisbX
uGrKODJ3DLLauaaYpZan5X6gJHHbztor+osftQiJe9dVUnrxxpFD/oQqYMgMvALCJPIJ/+Zv0Z0A
EEMTzjHbILiD8j80f+ASsEsqcpcC87gVRgBIx9xjedDZRvE/yv2BKeDFMYvbAoQ9WOhV6EfOF0P8
DU0tgMRHxIosWvRFB9X8NemGZx4osNMqrV+MXwA9eyjJnuU1wjhxoIvBWs8b4sKbFuMRA2zUppGv
6yajW5GTznqoo+fepiP/3WqiLyLE7hLY3VvJobYujLyFbieu8wHDoS2TF/hvngMVhEF/S6sRDpRD
D2U4gvmh8rMM2HjTN4bAwHqwVMKaQtC6RjnV+8Y3joXy052CQyg44MCHZ/I89bk5SLCNhUNa0obO
ayUhO2oO/EIXxxQcU5cTs4jgCPb94REnx6Ddgb+CaTu77ed8adRxstM0J67Y4WEyL/A1jfqwyrrL
e1PSV/sMbDXM8HwQ7uPhoZHqDBCsA484+zPON07Ap/YNNUG1/5QcZ72i4WFba06jZSvyvR7Dl53p
6OVIhDWa42xCYEgOwDslBIcViTCPPmEQHK996wCIwrlQjwz5T3V2SgqGWv86scSKNYJrMfNzT+sa
U5VVARbqk/sX0r7d9HazRKRjfsUq98LIbBHm5iEvWWMUO5isOvU+yIoaNXjeCwm1i2MCue2SVCES
OpZbBr0M2iIEHxno303ARgjTkxvNtSZHWA+gYzT1qwnrfkSu0dYbQQGQpmTb4bRDrZ8ftfUxPUGQ
Ilq3syZIfPld1hJktbLH6dRrKAlWYJmoZiv02KUj2YdeAgpHWY/2ViEruTDetKgSBiem8XoxbZvL
T5OlKjKTUyeRIUkWjfc+EiULKljoW77Py2PquBwS12/2Lesepw2k0EbNh1YhWiz6hhUnJHX1mu8q
ik1qNpN3qMlWST9JGt6l60AiFNqXqK+MAyT7tZ6/qpReotWVCG8ApAT1amtcty85nfcoS37QH4QQ
p4Z+cWu+hoDu9ZGYMU8WUFJntq8U3fEN9TpVuzEoib1HPTNstv0DgBIkvh/vxZqb6ddfzJUY5gEh
M5D/8pGMa9jC80cqKvvn2o5RtV2H3fkDRKMPZva2ed398tU06sEK6nVkKa5odLw2oV1usHORE7MI
eIN9/8qTwA+HChc9IFh0v4evJZt44s/46SNtpWfqvtak8rNU2lkfVywFMNEoaHwwUChMpuuM8zhx
hXyp7D/NbjopxnvJQVA1pyiPCHf3ZXBpt5SaZtFfVJuzKp7RbFvrVHwNq/Biw1y2zQyPyxsVBSzw
VMjkBLztCjXjYr0Z5Xb7l0zwfidMYJGXt5Hx3+VgC3N3pQM6bUgNg0a9myA4v0kM2Gzye+Ltl84A
Ih/ZfUTVabfJ1LWmmgS5B2/4r1/CMra3WYLP3OxRz/ZwHK4YLyp6BHjxqDGrwkMRLh3XfnfC1SUl
bwowVrPjhKcKNNa86XXu4LX/XvUDBscImKYjstgiEk6ODwyhMyajYzYFbK5O5OW3at2ldFPWsx9J
w40eoU59iK+MEVMIIdU0PPby1wODyLKyeJSQ6sfI27D5CL3vWpzlz1BCWRv5Mrcotl6ke1px1djV
Aq8TfCEkZBppd/NNqPaodwizTZW2FcKHeZTWS491hwVBnECXp/gPvixsIuaJRTLlb0+LJ6RuZdSJ
ymVtL9LE/04kyJ7kepAVuhPL4b21QWEL+iJ58UResr2jX9w8sBMmxU8K64BrbQBYlx+G28Qq/4x5
1tBaxtUi7sVx0Gcf5YymwZYWvAu8z3oKP46+GomJUb6oPOEjQqNCHd7UOZYdJLCN1WrJVifL4d/G
oLJ3NOifhb8ITFfkFj3pIq5dsiYeBobgxA1vzeXw7iqR41itjJuaQpjJGG8+53WIBP3lb1coAj0z
EVSHBCcOEtEeuSh9Mmk3/loWCsPu8ve/zOVQs/EH5znYpUyxUdhnGaR+xqlmxhZyGhTu9EoCs67Q
jer6HLsv93wqmFW/tGWQw9MwpczUaG20cjYQMhb1CyCE00ZpbpPUx93uI5+fpXm7kJ9OWN8/5V7d
cNAPu47aXDquD5lMfvm0cXyt6YAIOeS3Q9A+O/Sm3oUgbMBv1m0A4yyLzpa4QEm1cNGMJzQfHtTw
ZhLu/8U401Y/GXhmP5PLaTJaIfyX6OiidApbAfAzI0Mw1RzW/CJocPD8/yOCjo5gTCOshJHD/5c2
cNfYbhSBe2PFFLWKFTi6WbqZtsIlwhIXav2c3Kf/de3xVCiR89IfAHaxmkXdDlxlbbXf/6qJtW4z
22n4A2fBvlffR9cjsxI2pQy6Z2ejA9qpgJxXCtMBXpZS+Es3eqHaBmVhh01gQwypT/9UrJz6T4K2
UOnPzMtbESpg+oTCxon44bn3XaSne4L/b5etKbunT2mYK5hJhSRfWH1gFuFES+q08AwFIS9B1Iwg
tdenKhWHHfCtbHKiwscvS2PrtQMqwcszNtMFpXuJJj9q0fNJXuy6145yiELJlahMsl1D64ITEPyS
mYqG4WZCo0YfVTX5gyZjBJf5+nU8zRttO7hQiVTbsw3hPPCMtPOfgaAvl9906IeagIrYtqWiy0Ls
U4ijHD4zP5tpXsYBSkkZO0QRLjl5S2MnTOu4jYAsp1aut7dUi/Tx0Jf48HbHu8xEZqZm5ZxJ+9m0
mEfM6ckteJNzQFWt6u5jmKqHbvnoH0Q2J2QqmEAEUOGnXQig6oXViRoa2Ry9VHCOjhbIXSkUrGqb
h7ZgAN+I2A4eHKjuDzFmpcFbjsoOaUk8rcNjeKjfp86EwG+Aofahxv4UhrcKXuDRzNOQ3ml3wslu
tHv5Xdm+H9ryYBCOa3eN9+EyMSoEViJWXp5cCl7v/WIsHFp5ZH3zzvqnGd1daDaVgv2gkYAtKVb/
zhhcyUk5mdhMtqbq5R1pN1yJ8kIYlztiEGk7SMGcVprHaDeMVMuIHhUTLJts8XDr2Qt7u3upmOWG
JdYg6f5ITjjsbVZdekVIJcgkG/Xait3Yqk5p6OUrxkwnc10mIYqFok/GwOOw0pdppzpBsuJ2EfF9
/wFzORZavVs6FFowZnmiQZ8r5dWhQUWXZjI5P8mmThCI7yhcZay4KKx83GgkUtVzOZde+icF9qGq
m43tPX7aiFUhI4eKWoYdzRCIN49OzY/ja+vBFgXK/51urCN1q/kduTpDqsWKFYq3mmBM8fZk6/8y
RVRb0OSIFNkGZeVVmXRnUpKthzZ/aoOPsOZ39Bo6dh4oFd+s/w+sn4YDU5Bc7yFhCqGOKvuovw8a
D2eq4yVJslT+daBYMPgnkDqavm/7a1SGLg6SmBOP+9KsDhsYpRSNFJBgT1nLJfbmftqFUDSZwfRy
9DPp7R07sBpgvM/+BuJHSoUrB5c9SXwMuybf8ie+JE+0ZLhlbvaD1eX/8dNMhECpMD9Gko8GRvWK
GClz8dyleYe1G92ZraqI0zAZgFNvO9S9iZUZG4ngljCSTt1DW2BPUzUeO2BJPjDzHK2h6R4kz5/I
lXN1o9wEMls/vs401nZOMwmfD3d7xSsLijg2CpoYVDY+rDd0TaPpumbVoKtt+dYwyScMb4RcrZL9
XyEqz4X1nkmLOqpSBNz0E/Z7wXVL0Ms/KSQHFqYA1pyzB7p9SdyYb8BEIFhIw92JSX74W9EvS7mg
sLLdfwxGEjgViY1njqUjoY9q4seT48RB6iS0RZrv/AQL+ZeIxOyXIbmRZEacJb96axy2bQ2MWlcu
BvyW9IIHssHPRsXPovi+RRpA+N/8anFwFwNj+5zldgnDWnkOiizjkJoMvJF4hLSfqWJIqQjRJuj0
zIRO58dYxR1ddhnfTcHCQJToomgoALd6Oux89QE+vcx6o7AHo7jCLgcbrzPekSwRNUq6PcH0GkVW
NiwmoL0ZHpq35yQxiwol7CMS+G0fBGwkfS8xqFd8LB0Ct/HW94Olgfm2GaQtXriyMpfCpNOBtfeL
vaFNMZY5h55cfqGR+vX7BZbxJggAHr35RJ2/te6/kxSAtaxcuPa2FyM8hft1Kxxsvq+/DHeERg2F
KK5TK3kDXE4l+bICB3OOQrbBhvd4mlkncz8F5Co+PRclexEP1As7n2qgacYdQ28XaLHoPPJ7UJbw
4LiR/R+Fd0w799NNxaRp95dQf2az0DRWdkehK0jrSMPssP+W774ZM/ls8yG6KnlgxOLiSIMNDaQf
lp/oa8yhkm4mboEPbu8ULpepotRuDLirEAyM/5M2bB0llUM2yMiFx7+xPAjP/owvStUxAoaxmZGK
6bnnoonMyRhqyaHkkoA6khcj3VpxeV2MOtUGMZfRJhymtxyf+IPNlK3gamFoeV63wO9ITXttk4Yt
ov8RNTGf4B07sVT+3rkLv+USbNgnVlbVtJsg+R+t+7SNSdGle2nF1Q9WW6uKbhNSSwh8i/OVqWkm
8G2NSf+yBbT4rn04iN8noRaO/ukb0l9aLt+fxJ0pzgGk7MxrZO2iUHBAFeOPxxQeDrwV5A6aBOet
yp4l5b6f/g2I15vgMlIIRFCvCxT1HjzA2MvVFQcX7v2wFDPCUY4J4xujgOwH/Yy8ZPXHwpRRPwMa
KEra7FO6ewchQScYbt1eJ0KSsAKT8OFwxA/ols+rxmt52hxVdrEFGKp/f+coXmax1x14Py2dug6K
AHwNys117a3ixR2BbYnc898ckkmb1uD/9kocHF2gllZyccTdSHPqlpI8UQrpkXCnTFTPztzU6ESc
aYnGa3k+P1HkvJYlDQvIolelDpgPsyyx0umD1s+nY+3jLqerUSXAafwSGfv+pVR/+p+tcX1E8gxz
1l2fFMt1CuJ2UCd/cmBDUw8wQtWH0/rXGCvzy7o01bfz2hSZVBRsVBNKFg+zx5JCbqAiZ5s6S+AY
8x7/rxVv94HvlpbxvKOKGWiotpolgkFlwdhaDuR7OTYe2xiAyRKqjhosKqnJuTdoYnxKNl9QC68r
mjNWWOPvaeCD4q2M612YDcKXy4roJl3PJ/0DQAXUaBne4anbqJgY4XF+O4B5iA++OqSm62fQWclN
YIeQmA6Jq/DtawUkQZbD04i8LwdMYepUp2aVINIW6hVo6ewN9SWtAoYlwo4IzJxbmkSIjaoV0jma
SWUxWRADRTBKKeJWILcqRNfkUO5ja3/z30aVbE7FAF4mF16VvV4NpWAXLCdZhNEjuBmEC4Rq1gCU
6jdUn4QmaKfQcXsPdCFqLGz7j5Ix6j3EkHR2wuagOJK5TOdp95hsQ+Ku4Y37BcW7kDqpJPtC/Em2
WclLp+sxN82bFZauX6dS5Jd9y7Z/ZDkP526zPsTSpv9ucwsMbuaiIq1R1E3Z9JflgStTZMc2q8qE
Vzh0NtrrbXrzKYGmkZa94+mYhNQKXDc15UbYEIp1/rN/8Bh1qXv4ONTQ/t6NqFpQ/hfnpy+rygJz
lxdmwm/8VloUp2QttH9z4mRsiLPLFeI45xxAtHZ2yiGVa+AK6Oax1U/jvrErUljUlbUx9EjTNFC+
u9gK/vtgjzcyI+sDtczcmXl78dWdl44jzdL2BiqmDjkJ/gPVCQVMk2vL8Nlw63Cem4zr1HAhLqZ5
DiPDZS7rRj0tfDRB4pWWeWdx8HeZKP8e/+aYbg+mC9hXL5/nqpVn/V+QbJviewjQ7ja6rscPDttx
BWQlORpkGlEpxBAGFQXeYSC9dTpvQpcok3iTCM464GcqeGCFk482rByvXRECrQhbA5s/ADtgFMHH
pD7jtiamVl+094zwGKkVWraCk3FqkWb4QIHHuoJDuoaQwRe8LdBNy3H/F/sa9BvoftZpxVoUEig5
qBGDH8QHObyw/Vxwo/FiUa6wk3VWBTn02wugpkx2ZOeLy7DNEsD26aBTP/2MNMP/ryMXs5YGqbyz
Au6FzMDLUdiu1tywnZdP0bqCQEu1HhwKePMXamOzI2cACFy3jrM56seq6a34GcfnfFTm+EhOtvjP
g1Q1inHRfJ2nxHPay6s6BPNcLnnwDEFwc5f8t/KVaRUHdJRWDFH7zdF5hDFfNfTRon3Sl/DMqafU
W+FuvXj8w/L4Lkb+4KaYP+c/15L2iYB09b1ApaCBSzn6XBcV856KlB+QfHxE03chxhDOkMPy3mfZ
DcKHZUNZXqTKQkRqYskOK27ulLO4/TBT7uI9vHKEaNiZKiNlhesGz9wixZw7iTylsnQ1Li3UWprJ
NALg/iTUgPCGIOBEvnHrs0Y+Xl/nAZuFdJcpeVkvKCpC5VDhKHRsEvJN6QV/s4WoUiXYilV8sxt3
Q4hAQxS3sVXG9XGniCpdkE9MElRIzgdkL8jVvtgAlDoFCBUp51Oelk4IMfeMw4Q2BkbTGG2Mmq2Q
RkMh/fOrNqwuZ+XeEdHWyTgbD4Ohvs4krze9unGjpRufT1RQ9jp1BwW3VqsVvNC8051gPLV2AOoc
9rRV4r5I/yT+KyLH+IVUW+xRwyNyZZfR61DyU3Lzj33olTWRomVEzBOeDaGWN7OnZgzkEUH4HCNC
BO5vUyj/qX+34Ul9UCzj/OrnGUn8p5tPMNjoq/tgY6DKy/CH7Q04O02bX7eEc5czsoNC+WO+Owp5
CrZ+H5Wi8R6DXtQsP1pyS1WmiWXXzzhkJSVA0b5LXFo9eF2iSu1Xn1/vhcAlNdhkAYlbDjH0hs/J
q3QBehWHRkk+eV1xdDHA6kZkqJ/4Egi9vt1jloZJgJ7UfaNqG33vaGK//4YZsLGv/jKlYKf39SsJ
2PKoIP0qFEOUNKmK9NUw49hPW197aommWZ7W+iTLcyxa43mfNANa5lbQpkRRxgIcT2rTBYS79aYA
dKzmGxP9S1LKuthXeFbLVI46le/EWOBMnms22NBCMJOnmDBnWIHzKXPCzE48+3GTv05D7XoaLnU/
zB9Jd8ZVMhdOyBxLj2TCSlHRwPoFifEpwMTMcLRlVS7Prxi65C/MnPVWXkK3gUXjWnrsB0kbKTmX
4+eLtpHWyFV+TIsEi6L/J4eJQ6f3vh0BwcDPdK4klETE6hBZWkaWyCgIN8pLktE4lVIB+kqukJ1z
AsJCvzzSBEkbPmsgbQKxHIVvkPpa9m3HMHgbrKaGWZaS/cne6Z1mxFtLAbiPl7j1RUJK+Gyw4HJb
RMkUPkkwgEFAYvtO2eUtrEbMazx3OL6NGk1Kp0F3GVLukXt5iZ632iXp/lZQ8zc+/nOsE/4FF5aI
F4H4RU5bx3ohse5RlhYYO5Z3NDMnQTXJKcvV3+zsfJkRWPTynvEQf3wR3ZPSC0zTVZ3zLdp4Y4vX
FfGwOz8EpLjrDky8GL+CqFossIk282JzNdkphFNSv2/IVTGfX6govSsMKAcUg3grIbryBtHrh/UV
g/pfWU4MYXc4rWh7H9lbSgcQK+nQD/UAZKPwHIztI9ui4+UDlB8NRQK9MrLEW5curqWppzMLsc4t
VGZyM/24R4HMb/sGClMiMhuBWn2Hn4DtY6KSeA98KzFa/yleTNjf0kHi7NSw7EhHoBkK/9qvhwOb
yQTrkuDhfVenRsV27+TloVRxis98XfuFjD/3/539ZNG+axGqaXszCkNnEq9WL7M/9XCAc0+d7DTT
KK+c0gAlOOEBYgtuDVvgYmwLB+ODeOXSPxShREsbdWxHP7u6tWipppmH9WdruUuzWRcWt3J/hQdw
vXjUZhxFYiPb3GXAe8NR4O49c/b2i7TmPq6AX1Cl48ooxCjdoIanqnzkSyEO8RmqN6IGSUrkUwoQ
aI1iFqZXd5vkORQqMmE30uwLzisyRHlSDgFtvOSRn13kUooc2/nAB40r7mU6rQmlkR+0sarUpHJv
ZC8VYOAKLETIbctNy5sgSbkgq8nXd7lwZZF+iilLShmPgFC78/nIubAtHPe9rJsXWM1ihcLu58K9
mMy7AY0eNqTa/SMOtGMO1Gpf7PjEHJuRk0s68hXffTaiTbq67AzaUHMrDqQfN6HrcbeexhBT6iwm
F5qxt+TuuKA+ijv/9D3vY/KIWF54UZAqAfoAPEijjVGXRcFr/wZXFuBYzddy+k/8sP1iy94A8MW9
3ekX3lUvGDk4bcVAYOJIweiz6WaseqeDd9dt91rAtwa7qDZmzloLqGo41T41atVu7mAJ8nNUADj4
exI0VaDemIlEUk7q9q55Qa34fBJAwxu49wBpVKh1pdo0UGbjrb5pYkfb/KH41Oe+Pa2RffNcj+1R
UBkUUsYCzc4LSZACC0ICQi4fYqYQdLEt6esHgDmjf7p3Q40otO1zF60b9MigX8wdueRucg29ru6K
QD9Y9OGwBYyjJ16d0p/nVzrbzuomOFguo63+a7RfYt1KuUVBEsYBgfaTyqiNIkHsZ6jTRm3NAGr9
W4bxjjU5ly4CPSox3JsLiEclxULd2NQg6Fj0SIo7AcleZ7GvQdVlERvI3s07XLI+5F1s4szB78Xr
ASd805UAJB84E0CyvmUmlBBcO7cV610mAKcapJob7+AtXGgM+Zg4QKZIfRS9oT9Ywyhcpwm3v83T
oFcvBrScKHu5iVtVrWUe2aeFs0f7ej+gCqVD7Up4vrsYJb1NwAYUDNlLs3p8JDeYVVfAnWIkBo/x
SRG6ARXX+uWZiNadnpi+6Sx6sulj+Owt1vPyfCwwv3hX2zPgooTtUc2q/yzxivqMGouhthCVcaFe
iGkcOJ8CTrr3W0oT+YY/72uiUqvL0CrXNc+0aOeCLD5vFVQIW8/7jWt72YKzxzhVrJA4VG6OM3pg
JkllMwsAt1gPftdNjGOti07n15Bu8/epR0O9mvnspV9HIyYYHAXjp9DqaYGqxNGqYcp/73vZZGN4
8RztWgVQ7DZzJXTMQAhVJUyDP0gyT3DtGKy4rVhd5OAF5eID+pe88q2/lWEAvLChcdo1xTuBi/cJ
J/HIVYyZV+6c4dysUZdBtwU4z5khK7EiJKmkE5+0aVpm7vXed7YhMMwzrmg7GVjwaJEsLk2jKdW/
D8fnXO36OSlAX9VQv4CfJUe91gEW8e51VulbS1dhUN5zrpERkX9ZTTXFvPRULMTRop6+VjE15OSw
8aVmbs+Bw6ZgM7ew4XeJqbj14IDaQmhXlezLBer1k2j9UEnxw6c4+mq+XW2yoXTPUz9e2hx7edSR
PcaMjwL6RnVtazCTJBPuQMZr+QoVSVVrHp7v/zo/sSWzFZOTUAMJzl0oJYWlw1E/9fE3g5vEFLQW
zXrTe9dG84r8IAHqplfmIv+mISP0wvZwpCx3ztZ3TGgdmKkMfRxTSmlsamqWizPI5l69QKw3G6fH
PsHScxtXGkzNHuR3EXRLfk5nGl3WmdDM8f+Cx42HXMBgj3MFLKMj0CQ6xKy4Vhkl0IVVMmiCzGaT
J1hxEqeVCeWiq6OPjVMxJoFiuR6IoiLtpR9P+X2OEeY2fp2dzx+qNBKFrekz9G7fTMlWzbaWcOrI
HVdITghmSRNmsIZJjhvqAh2GQoYLDd7x632Sik4+m4ix1TEPi9ruREsKfQbkUfOv3LPCGUpgm6Me
q0NHtxXrPkKEB7+WS80YkYHCNOXUDcStAypuqUtx8jfs/UyCNxvR1hFHoxE4FPGLcMHh352hDxEa
vYg0sM0S/w6aKZdWhV83nvgjtr/ZURycOS2N9guy5NfbX9pOI6/9bf3GsiKni2zwoQ81qUZvgEFx
cX+0niyEDHIulB8u6My/3IC9Qc6Dcg5i7EazZ3B8ip5nDVCuTBLQGcf5brkalV+0QL3GumqrRTeB
IiqNDJvfnzWkGcM+rOTAdbcoM7cJMagRDgX6X378gHeSmM//BayqUVrX+XJPL4v1hkJ99aHwmtSR
yVAuhVEXjU0F6y9x6lxmnqEbWgRvI1KE606o/Ax8skjrd2Tap955vjINqyseZfLaYfmmplgfrCey
Z+OEY/Ye6/JENydu9vUBY6lCIxr7WpmfJ2KlLxrJdWryUs/8rTmE5l8gKLMsCufqy04BcdGGIAVz
7ZXWtEH0u+sqk6fxtLw31SXkzqNxqLhBsflo+9vKR3HotprQGVNDpc5aVJtOqmo921CE0W4niJTb
JvBKh/Pu8U+F3wrqVsdAgVR1CPfenlaD40zJoDG+zXV8GuMNgzUUazaZHDIGITbQQo7kALqI6IlB
1LIn5rYqKi2ICuAdWlAP0Lx1BXejC7Rm8y5LL2caY4aO26/MpUb3qJQ8Oi6P8uECqlbWe0mXEYLv
H+JuVnOK9mh7mlaiUh8bBqH3AJRnewUHJRUWRubHncIQ4c5fG0On76ehBQdJsdeAVt9uYYtF7I9r
x1fAdzHLhCyfcUWQ/UH9wOkB3Q3FSg0CC2Ql9Bot+81UKCuqFu3lWj9WkkQ8kkt9zKxtF12dRzns
mfMwnA8H3RKsGhHtNonVTfbtlGMvtIZRgcEtDGWGxqERm8lgQdii+0b6/8GNRZREYoSCrnTacq7g
zplLIqbL4OBLqE4HUN3aFaNBnigq8POfAdOwvHt0/+efEtkf4ryGaLWvFtploDUtiPyoGtb1HqXP
PFDmZMtaQW9xXZ1HmKPgB5guKSrJTxHQJjchd4ZvLxn+f4DQb695epdDesUPAi7Lpfk5J31+RulG
T7DCouv+O8KXMpTYS6l4VCXwjOvKhGm1GSDNfJeAEwNwOUzDmCCj9NY2+6LMw9WL2fHR9ssgjLXX
CxhyR+UO1DCy7keEhr7PhQ0tlTcuA/NCahbTrbpXy3VDtmix01r/manc5z+F9EsLjhO0WGjWTNpU
kTpK98N7eSrhbOXfudRNGy6EqOIAW3qV6pItId2Wx6/aBZW855PTl+gaoh4c0VfHTKbcDFVscqJU
Z5p9L4woMJeoByi+Mu8QHDziYp685jrJmd2TrnqKfnB3qdtudM/temOwATw3Mkni7MYlVtc16QYs
7rzhTu0PtPvQA8o2FBUq1jdGGHEOmzkdhTIz2hUjl9z5plVCeo7/uSsLa3aCkfSRxXj5IMoZZ8hG
Yk0cOj3aX1430o16UrisgaHpV6dV9WAQ4QnQFQGD3rhkmrWD943NNXkmq0OAPjOlX0AATzEHHNQ6
HY+sjk1K4AgJ0Yh3mqljxKNSHwowsyodY2e1wHsfhKR56DHvPJo+xQoxSlwAYyQhyEiZNLa1nJ7d
f+QvyGjzKAjGq1BTWPVv81yHHST6eK+F797CxP425Ba86iIznGb51IZ2sy1AOytYMbIC1NrXJjZp
zSZEuEc84lZezF9Cb3i7QwKsc5gI4sj8P43aKItwxKYASqIx7x86DSKTG/nDgCjxvJqFNj4SG3uD
GmM1zHt4jB4/QMiLxO38c/r8x/FztAUSuFMnds8lCSuZ61jjcqyTKPMCEzc4Zt/szvJAPUSVfaHy
FwQY9ll5mzmrPowJYBT9cH3UobgKFwAkeXsFyjyl6iiUpwiZQOUC9Y4KHt+LnthrM965BGsYOu2K
9tdrv/bN5vXxhp2pMRgyUlnrb+TSYUTiCyci8yKEVOUTvjies6Q57FevUtRBPKfaRsPTL5/K5Dka
uy+eFlCw1Yb2wesw8MSv3VURDjH6k+d17HFsKwt/wdwaAwDe1hayExYO2+Av4KDTAmfhvkMCYBC5
0xChjeZsSag3FG+RKKrqwNntOg3Q4g8UbDPjUKczKe8XW/4/M6ttgxxt+TJLn91nQD8F7KgvrmH2
tHnHupcCzDVTHXj+sM6MdKMaQm6Yzf2HPN1PGQLrMgaviYx6jSmbSMgidGfrebTqLXDYcY/ht5ZM
mEUa0fOXoL5C8qvW6/Dl8saUQZjGgl2OTJc1WjsjMGDBPq0CaGxw6AY0uiGkzE6P5hS6YLkv6Rfd
rr6PB2vqBzPLKPgTWo2op17VUeLYTUhu4/82ZlzLdcHP2ic/C4toGbirumtDfZz8KoNNM1m+2E03
Q9LUxUgLjxATdvrRoo9VOXy8o0oWTxNau1PX7BKYJBzMdmyzO815N/RotTwGSDTvh8UYU7grUyT2
r//PR7IzRjQR7O5L2sd9j5rLJp17r+cFRNJksWsKpv30zCsFCdE10lJjpr/XLdeW6F8iX6WTNkcW
lBPH3bUb01q99Izc7Ro1EKFb+W5FJNtfiJldmBI3OkD0K4ypejRTHgEFBtuK2SFhMja7gMxzGk8a
Yq54PkuXQ2ijxRiVNfrr4m/2TS8MCIPphIXO9vE66twSJseQbrj+AWV9hjboXemL2Ky5hyT0yvy0
DCzdExpRqBrtqtmytVmGwDqfUTBRoNORjtlxxCaalAQAiGiApzjwOLIansQG1vzXh2cYz1mm9c2z
ovTMMao+vHveXF+4xlTHwrANbCT/wSkdOdMrcrHv2nQeiB3cbZURv31kNP9HxjlcmSX4YAEdvxvl
t8iqEJjdsyToagWlYFznwlrvNwkAMaeFru3fDCDfYoyif5YMU48pV+FDB39Rlt4vikJ96KobLjYs
pHWyh51SpsNAd76uuj6+Ne4zY/MFGyoeEZQFqLHQv6eZCOb/t+zYTqkAijOuASNs8n+0wD1YI3kd
0XdfOuKHHXKy3n9OTyfUj20pPCGAP+wdbBLPf84HBgZkjxvKxQaCSXhv99QM2+RVM3EwOVELtN4J
cvn8dh9SpmVBwhRUFkAaTI0dj6GBo+WBIs9IjCTlTVwG6G5OxO6qsg8Oirsr79siJL6j6UC4xiD4
/FY+ia7mITPQb1xyo5VNRVPXs9o1M1YXPDiFWBLwULo2e2o3YTlAcPRYlJPxFWK3UsRNahqRiTjI
+nSOQso8Oxt4oYw/jybzRscCxWtrY33aIXwZtXn96Flcz96r9D94bWmIzfV3s4x++r5/jJyb3Xbo
dPfsGi9LiXX8p3ovIRVXAAtZXmZDKZcCEeL2yAsp2P825lVamW33SqHoEfye4pdIWx7gNjx35pEj
37ua8SYWQgxYFSe5oOULTl1u/bF6t5hEJmLxfdxgCrIDrV8Qs1KriasKB86+/b/NtOYXAHX9M5Bs
0xJPssX+02eQ+5FNWLXHK9mbhz40h6I16xxABYQ03mUEIrsPuGwJsUL/HPGL/nYOIbdl4NbZ0pC5
QKtpcN2sVcIXT7XtWfOD2bQ6gqMmkLw2HO4G712lhB6cbHfOmcQug1XdYE3+cO6jZiAVWbp+XIsW
Len5VLVie+bLyDqRnQdMTQoQdQtB0TAHNbl1J6EhBv8i4C976Bgd4MCzHe+qZL5oy3b48wGwZtp1
fTXIroHcylYvgpuIiJCsg7YLrjt1xJD2QTbMyG4wybnLg4jeiyZ4Ur8A5WWX4QtyjhiDR2IFHULs
dgyrc11cjuhqglzBhn36qXp39BXQsgf6VZ0awGjE/Lxq01p4XzhMvlGulbCZANU9HX61XcS3P7bj
oabfH8rwjebUsP8HWdqbOPRJBXqMHfQKX3hEKhXz8JJD2mJP6Y8o5LTH8T+AGbTD+lSHrlbMs/M/
ldrA30YsulY76bzlZW+5G8Wje6VQv6BNHq0AZVEuuicHgTpljCHTM5yl6i7dRUm3r8CPQemzOqgN
APuxiKRnBaU+ArTF9C4J6kgCiFx0yKkKodyIJYu0b3ppPhJfTdnC+4Sr5/+apxe/4oOC9UOpkmSh
jrGQZgoBBFGhbNZakuVC8hDvx21GUZf9YQQ4lrk9DMyQ7rXZC7S9hQFB9hcOPyEJYe5zmn4mzsB8
B4xK/O8n+98qFeiAriwGCQt9uM9Ou5DYfn5mYjSPwgsXb74maF2LM1J/mS43nh3ZCxpqgyWsR0ox
12z2AZ9c5yRG51Izw8FrgGHJJch7CZvUJXpLNMrf2nmhIEW5QCujux0sXfBi6JMxNaVztIuF3Zsl
rohqiTo8l97hS1bwiafDnuDgHSAHWuU5+oAxce5zqwn9iME9TNBhC3Fc4knfqE0s+A7W7aHRvpRS
LroNZ7Nux6vNkEu1CAVZHi372XfomctbU8oSlBxbrwvx3h6PlDOho1mOyD2LxF01hBgNTCmr7qKA
yAC1jL6bRhDwv+IdmuVTCknVDBBOAgcZaJ3+SrZOCgptiwLuw7vn7z1/ZkR4SuENY3jKVAsCdfgC
9SOp3wFKPneyrKDLlpMBoCGYg9c4A6Y6VjwzNN0F5egcvEw6CZ+BlGWk44lStUSLAI+1eQcNXbD+
EI3pLrK9OMKZ/SjCHw/BYA4emTSlgy5K4RJm90oqYbkDJCwV3SBELTgBWaU1WZnJKSJlQ8C7RNs4
InJ36OGCnaSs+zIqYped/TXKicGquTxaSDupIkM6+kuwk75hT5IyjNe2YzFF7j9/xkdj+XuPpp/w
vuByJkuOCon/V83QeI/ifjInDFOaNGRdCG/f3AhmDnvw16er3NykeEM2TqluqhUVrihnDDz4oNXu
DY5W9n91DtQqX4SUvbP1yxWuf8aa4RJq84JEZvD2SBMEgruCE41VgbgbgqaNRHZlP8D9uPeGBGj4
++ywpIvsfempOAT6ob4BdfuiQ7hxBKJiZ1M1jc2iSpzNFQYZ/GPt4C6RJv0k6bRZ84VsNvgr4rBm
j3slkZsca6TKJJv5CkPz4LPs6MaufQPcBbMcEsG2SBASLNZegTcz08KNrkxyI8FAYU6wfBrQbagn
pgYk0gE3lRFZaC3Lh5YoX6F8E1WRkrqq7T+lIkfq9SsNW1ZJq8M+xB296OkF25ODH11weipCVfFY
9SKrONhnsooorTywzUNb/Ck743+R6Oy1IH6nJZG3oEaP1rdVQ57b/Ng7qLXoJe2N6sgkaUWuifyA
lLmwLFMoHEMZ0DYacUXmzxjH9ABHX3o4ptqqFhS8A3T2edpOxFlnNCJLwn+YEKuPF7XFhQftTwpp
D4H30hbCOtSff9T2FSgI87J3+Mu0zPi1j7QM7n6010cfBfJ5T7EW/iORWTriffd5cMa3/JdnF7AU
z2eZtve6XVfegLrhc55kU/NyWxnB9kgbFAsj+aToEL4ZV6Mfxf8tyeetNLThgyAXc44zponfuS1c
XHikl8ZA4CC0CtBdUSGfkg4E4uQdt83AtYUH53FezqepKVkVH+wc+gEJ3TDZGzkuNDFlpBW3bS6u
WvF977TzbSK1mnvLvspJGBrcYmRf2WNJpXawEQ9/HDyU4KGZ9UwU7BC/wbcJy0n9wMNrXMC87MSA
ezztAAgewavH516gf7yRNQ4qm+E4vGvmJISos7GhOCwto6e3HiSm7rr1tKl0HxS6n/jQwugPhAUp
FLD9yeZUD/X5e5op4RpwHQx8qtPa8Q4u2LuoE78ZaKC8x9618bQNS7n2NINxcbdAISENHGaEMAdw
GmSEq6aAaIUfMi/2MhRF6+iywEMJu0Lk17NUg0fJEHim/EQ9vjKy13+vrTfUM6p7Xx2C2UysxXlM
38cuLtAfpJck8listIW8/V1rh4ULjoexbL3wn+jgdXGVKq2jb9EBqfWTORCKdZKCeBSmQ2fNpIQ3
ik/uSE+lkXAPZWuolxvoWA8Ifx/qzq3IhXxM4cMKO1Xm3uodYwrcGSF4SKuQPtADPv/Z4AoasWF7
cmTErTy+sQE1blg4ovgeGVZQhxP2oXCj54ufxo1JrS3iR+stLbzkJ/HuED8LZLnq2ugl+5uoFjhn
0xKd1uib19p465i3HxUv1kC/2YeYIvybt6FQ+L/bCIusvIO91VPlwxFhBHTZuEB/mIjTfZL6Awsj
htGz63NU7TThxIdnWE9qCbslB28s2KocMBOSAONxNiPoib1NVYfphI1AlGPWFUIfNe5vmmr9ycNf
8pnMM2+uuxED98l2k6vPqcQ9UcrqyXSedmLmwpobXOYVH2U5YexKogqlexACCaobsaXN2oD9ewZ3
Byy/ykSFuygY9MjXLgc6bfirg2ymvEprH62IFeIHpkpPnTJku63xRYjg5RRWv25ifTOGxt1yCi6d
of5BfG2mnO6RcMo0C2MkezVgERRt6ug6M/4cxOUqUwDopbbp8/Yp0+EVv8gSzm9Kb6etaaBVdqSA
HFM4HO1erARZBTmSJSS4jeoJYm16ooYjKkt5Wm6igAxOBiA9sPlY4Qbzfy4nvvjTLGCKh48Vk+Bz
5OqXDCY9qKF0gUnv0Thl/9ZI0I4vqvu7FDawxri3EL5tnt9DiE+5oOW34YeVpm8pkkZYkpDLVcdW
dBIkCwgDgfESgbbdh42YpBmQZg72KxqDPX1sWTjNs0GmTl7QYmnhbB/tVMNABU+JHFXacQfYAshK
I9RtQqV5U4F34vYwwybUwVvqH+ooi3E2VyQ4C9KhB1gmJ4MOZzF2Q9RbmZl/4WA+d7esgYtFtpVe
LYCGuLTVOqF5ovfPP0GLgCcHOEih+TlT1ObInIVJqyt0dCo5yDuYYMsX+RK8OD+8cJ59fY0y/vwE
oHs8zC0HAKv8juBNc5f8brC8c9yfXOv1qey08Y2z0JaMvDzPn97NRmeqzt5mycGOcoPJ1SPqH7Xf
FVxsbfTpJEENnJVIogtGq02+0mvnK85uA8PM/qbra8/mGFToWiomZha2dhi4n/tMTorJRxIpX0bi
JZtdkuqoL663e4+83UKhYNBqtdR8COkWR0eqNCaqi17OvLyZL1mr/cmvVwwS9A12EBi4/KE1u212
G1KxxpNiWQQKFExSdNN2Idgs+W5LBOkm2g0r5Zq/CwLveQZQDY4MEtyWuJ3NxHoN3RJjh0xriwbo
nC1R3lvd482E2JGyxWY4OKhLMgso6BJb0pYgCL+bBCGlTMDSwi2gJo9FLRj4AXwPETdlqls2t4Rs
r5TOok1X/52VC3cfhQO2oxmK1keONLR4U4TzLcQpIl+BP69if950fdImxziOx4pWRUbX2wpWUW/K
vsNNTHaBSrY+pVzqUaSO/m5cuctISASHt9iP8LCtuKReoCqCT0ogyYv71XehjyWJe+tbd0Nmrz4j
UTCRKTHpmKDeudOMuHNG/h5LTJkVJuwGIy5ki+yAUOTN8IdezXdOFMQmeVCJNv1pvd5wU1IDM+6a
9v3tNykQ4coPavnZygih7fApwmm03J1SSTAnaJpRaV7nWaPeJUP90/Qh/b/OmTsA0acKTx8mTkOr
sev/wiFMuN2NxO59+PM97MTnM80+zXvqQ73BxLUvvY+V4hiAGuUny45GMnm0mV1kb9xgWhkbJ6RM
qzrMWM3+91QvzBKhQ9IgCcxVR0vk/NHyPP9WZXw755GvFCMBSnJgMyzPb/IxKmsDnZ7WJmCmK+wl
yAFAXw8h1Rnl4HsHvVir50buwNMkcWKs7gGpagV17sGGCGqNNYWYL+dYhTx7Z/Ms/JROROjG9emo
VeB3OM6+SMRC2HId3reeFdvBblAGdwlyK2lzFh1x8ZGfBA0PLbb1w8OqTI2H3+arh1BTmikpnSyQ
fVop1zYJeMl8L7PvcBYID0sp5FgPGBaM765XnhOtH8rLPrbzu83EU8StT1LGGoR3bdWEBPQ4zO4/
/dR8+DNCYT1GG7nQ/FqfbP7okPdXxU0H6/52u0hsm3tOu3YhlpASQxHYe95cfppgek6BwX1jwWmk
ak2DUMZ58/shq7NJ2tzTT/XhqDNWD2A94D7DQKnchHqtlwhMxi/XRamkTG57kHiJoieKrth2gZcN
qbfmXpf+YhfjC3HWp9m0vXspdWRSwu54JpwTHSnGNfDuRZxYKbPCVNQBISl2apgjGpINBJxjySvp
NH7t44+A/SnVC/3DZoIAjJ/1feMUZZxGr/T7LondhAjBdUZFdvymJJNww10u5lIHXsKNHm5sMRRe
7vAnFWriHEB/vqEeyYPlQfH3Mod1wJhm479qQaqWr92FFY3hb0fTTRphAl1ddnueVRi+SI/Kg7Hm
0Q/WYTVn8lHRQfLZpt+r5LsKTaqOJUesTA2S6f42imC4dzXEeywx91+yH7Uwye90H4GZBWJe2fPB
39pDo2TcZOaVBWdW/lvOPyVBBn48KlUHeOw/kDU0EmHI2EzFBA9mZGyI4opd7/OmOTY7f3CzwINW
u8Be55R7fNMBffOnwvvJMYbSEpLg6nxYMyVDaSXT9Z0pzjdgLBv0rxrTCvI0ExW8Iuecy8kob5Xk
pteNqjqO4ER4ZgyJ0nQJqOFN2SHZuR4QwpDtZ73GNWkPwTyj42TPUjzmtj5KRKOLOCZYP95EI1c5
lw9JE7xBcmHtl3tWQ5Qan2sFFNrPhvDk9U3ePl0MDwPytjOdDnoruhia3nHImSdaHwMHJc+EM1vq
Lve/Yc95Baa3ad/0zZpjBpNp6BSHAvcuqT9ouc+fDTMUZgISuQaggL2w3KlGAvjz9P0or+0cLa2c
m3x7Y1pNV8yk2ZxTYaWlBBkYohMOy1gQXp189Ecf8Efcue7pU8jCdArGQx0IOH9UscCQbZtkQedl
CGpYHibw7PBa85ZlPH1Nv86FMYVbF8xqLjrBvyfmzQkvsU1gKDHTEyE/FhHve2SqiCz99vFIAPbu
uuq///knApz34tz7It9C9C2tdl1Lx4R0CsVLk3zanl5QsouQA1BUFCOYhd46uFIf2QkPfxfFbzpz
Crj5JsYc4lYcZw9K6xTuDQ+CYl37ZRf7ZNR/t6wZQH75VopgNlmTw23644q8eDeSrLKu5WCTW3BU
N4sk7ZXIhSnnj0VCo54JaS6FivCWqQRrnkpoAg6q5vERa6hVRLgER3Iz0skl8NCfcJlXykvq4fRw
z+w6l6LUZ94uOW8zIakCBRh8iLSLN3rWrk32+vchRHXDTOMzBz3kApU/BMMRk955gncxLSRgMWfl
+KuTx9l4WlhyulnnOACc8b0fw20cQJJrAeyFjGPW7Ztb5F7wItZhlbeMCIe5wi/BNPQrHpPzuyuP
yAxPpNlR2OAVuEoBJBQwW+r/yYgiSzfj97k+thbW3gCeuKgrQ+tinzxi8cjh1JateRMwzscLCSCq
tYmhjH4mGLF1XTBxNtkM7NUM3Jb2mpC+fWskOwMFbMZQkHzQL/3OXK9ZpX9gzJwm2XTCWbjjWUMR
11bas2Rntjyhr4FGPzjOvjvZMTb5IvQNRCbz7o2flEK6XKi1nxT1Ob82+9Q7YrssHe3N3mWlPdq3
4+f0QB2PnZrdHh+YjnwJdXAtDVEVle8IRv2Sz0YyF9fQ/TjDMUwz9TSfEvx5E0qf4Jt4eRqDO218
RqBbW7kAKehrQcRIHr3gondZkRuZ+GHAgEnrOxblYbZgi4Exzy6RJg2wMATjkfzYQRjaj/UQfdHN
pmnarlYjC7NGT4gdK76ExjLHavbDIeY0YWY6JTbRIfqmDhwFHxj4jDZrTck9jLIi/tT7kwTBKrR/
cexRk77wD6RMQD3aVVgAeEgwnHAqfXTsEPP/t8MdSR2KcUNwxSPpA4QPJM1AhmmePMuGgMKxMJce
3YPVZIV2hPUyduJAiyfNU46UY/jHNT/FNTiWISVUUcnPoGUkFjIwya4Genh+EPaem51qDa/NxZyg
mx0qqZ/tzwTqIOIKdINTiMh7skoRQXrWoKoLV0gPv+vAruOAKYmyzCQOiKhwH1+VJi4dlxdYUZs7
rOuravAxuMzkdNJ7T31YhCiWWNIHvFxSMAUy5BcH2+BQ5Sj2G7RPyuUIqaS8IO51a49M6gzT2vUu
rFcNaMli1PmT7YrSZDFPX7i1Dv16HUZwDqrf0RHqTJW7VF8kKrRm5cwKewnCaPz1F1NojWzcZglt
EP/g81nhIzYOKiC8BwA47nTh2F/FpMDgHk2NjhAFRQOanOa+FOGhDoynMYJ4jZ6TI9RH3h+Au1Hl
1UX6HHW0VPcLeYkN0vnNlIKkFylvudlUB8l1O2NIUcpbMDZFofY5731FXwqaulkwDnB5LiKizFsp
SqBEoYC1wT0nzsPxmi2X+TKimvAo7iwGkzB2QwzfgmNkwsBdSyEOEBNh1L8eSn41VNw+VoE5MvmA
404Z5/dACSFs0mZ8Q7LEIMgbxwySHYOCtWArorMX7HfXK9Cl+qIHHE+3dOPxLjl4/ivhxlvnG2rW
CfLVhAMC2M8SnUY2qNbTETeolGyIxzvLeR1mBNk5yesh0iVFcnCi2k42ifypNJ+M43r6cKWBDD5M
uQDmD5DGjex8SBBCMrUegnBSQyris59qE6zSigCg/iZH6wgJKQxwcg01ejllaLJSgHqwnrt5Zwe3
Ep7fqqkNg64D+qy3LRkN98pLH33tgqnCQSOHbZCtQl4fXCbKm6zTqscroQ28T8aRSsajZJkHuut/
6U+NLm6niT8p6SmglrzH1qQGGOXU3meCDUNIRIUEwP3dckbRW+kAH4f81Tu4IeapGZ6pD29CG/Di
2jo7rjnrauulbpaEVH/kp7hgppB2QFHKal2hdW4KLcWdDZpXkf3IUBvG4zcYGab+cbSQjrj3aFvL
9GsAMu5Wi8GZi+PdBl47rcqzQv5fh2L3Rbr+Kt+PCOm1Zj6WPZowY9LvIT9caqAdQOXvBypjDuBh
u+/OC4vHD7ltFBe//089HebczpUoIXWsFt0naEMN5iHCJKURup+zi2lVJnsYU7cv+G83XDjUnvUg
l8oXthailO5iyuaKkle2piL1U6MxKohumUtbSJyLW+PE+6ifRcjP99WWVFGhgYwN7fxpIDHIA3Q3
B/PEXTsmnFEtvtogbvEmilCvo+w1hjDz/X+RIwlQn8TT/5T/YuTVpSkpjod4IYkUm4QwklGAC8+I
reKsJKBwv0i+CUjl4Ny4Yo8qZKu9Bpoj+RAjFhUxxZCy5Z4okn/k60x94C5XauQNEYs+suyhyFS3
gBxV2o7tcMFHKP5g6azGgoHwVoHtuhqO9pLFy4h89/AjZbSJex/gAin9ya3zrYrGZq4dioxSZpvh
fM/l9xhvd+/3VFUFLuATeJT5tA2jBpOIG9IDYc19je+D+hUYyEQC6Y36FziNLb5nnJp7tyhJ4l7+
MpkH/ruRTmK0In1ruPRRvna3iIWDocqBaIxQqv+nYT4oWTqHphaYxJYw+MXbMTVHIAkdilnSWoZN
gMz5Xm7q6ZVFg0STFjuHM1s0P1mRJECyKwVtBV12Q0oA3CNUA6QCXk+xOnnN/Z44WLdnBNLV6jbB
DEks3FBJdpylnmmQ07D3oyQkPZhsIxOpM2M9Ua+xcthXDTxsVEJHPZ9jZ9M9Agm3c1NckE2vfvKE
q220r8iLAbXEZ7WtCBJqc59pBPtsUb+PhzIDCWmRqfyTJWEh6A7Te+L7aAziaMiRFHIf/UXRIdAy
EoQHwzBAEq/fKt3TF/OSD8F3cCSYOzP8Q7xVftTC/A4U2uCnOcO8i0KwufkKRhfDSreORENFVLFj
5o+aVMi8+dZoO7xusGFZw8wgitMVpU721pAuSgVgCCphbMsXV67yx/nkCq4x3ah3oSAd5PHSA1Pn
TvF5QY5GmuCGbaJqHmFMXfJx6/Nf7bWY6q99TTwpNt5uAYHhChSrWfJOpTzuxxvRUKlcn8gAN3M9
8OSzq5pPgYy0Dcr8EU07/lTmP3yTnVgr/WOI97UIW6U6uv0lUygR9VtaU7K0QDw8Y+4cnDrY0KkP
roHBPEa4MERZtR8r9a6Alc/96z7vrhL7ghkAWHw+s52272e5wehMCe0NhmdUKC/SyRfIFRsIPUOq
IHNL8AwpMv4uc0pTcQJKi3Me3wOYRuJ05YAU/vCzxHytfImahocspcNG3VcDDfmLMqbJqumerBbj
fQbVyaVXPxcOmbPXyn9A1nHmZaeqNZY7w7WjFqGQOq+9w60tq5rcKqcZWkqXIyhW3I1jvU69PjdD
E+5RRgV257SgU5L4hjPwJSjmCk/VuBx3W2RgPmR+Q9D7/yW/0NIi1kS3NcH3gobDkq6Zoax1GRNC
hDhjt29DnLpCyujgBVUvtXKPloKR5CoSVgfkSCRM5C+CHoS5iKBWMCYgTOpuGS49i+xQpwfQlELr
NAcnUIpkwYi4bJt9ENrM0Y8GiQrOEL9R/KSfho0D3XKrfSmR777exnVaxQ8ymAtESdpQhzuYWtkr
fZLAljehUvJZggd88wxy7aa5vk0DV1xYXOuNDCegmmZ6Q5mpomsM26whRvFfTUhHj5dhjQibAUZH
VThaDMBL9eBlQvqHr82tG6r3BqQuFkBTXao6O6JiC2gpleBzGqUygj9diNq4qAGOOHIqIoDejcHT
v7kmaWRaEJVPtHD9/VU0QN+X88rdwuno9r3NIwBvgd69gE0HlEuQn/IoL6s0qmcb0GyoWIxmv+Rr
ayMoVV2a6EUPPZm/KREwVc7IlrJ6rmhslnc3mdG3L0irs3O1fL/arQ/n4/VaZMjMlzJ77grBmnNM
CFEGEi9vm0GAkuiZlSk/fcuLhviDy9/iJxgXBafWXm45HZnF3KWyuV2Tod2XcuX1NkZt+jGyoYvx
Cc3nAIl+oPpxZGWBklb68F9vwcisa5HcatgAh5+pIUJeCt1k2zv4iJeDntAMfimptcBliFlfP6x2
zH15MNAM+401SfZvGt7n7dAJ6HLXUptrIznzKamRekcDVnkBM7PboAyGO7qnJhWrUp6n9kv2qTIE
JB1YA4dGYXJqrjow7ZAP3Nmqv+BIa/nX7pR9AJKur2tp/wK28i0etbfYwyJ5QNzK16Ob5cBaKaDz
sxxlEENqUaskIEPdyQ17hGWRgD83ZrCaeZh9+6+ArHUDQn9613U0H99XmyX9nXzxIYk3+j7ohxjK
v3veprxMx2/P3ngBACNVgwwG5XM9t85NLMNmmVlxC7RpDCX2DozjRwkfNxZIUUCjnhG5n2p1e1FN
vuOJpPAiaASSPs1fNk1FNnl6tWdZz7irOLy51RYs5ZnIFa2lIzbabk6Ao83eM5g9SA3LmapVlpq2
X9OHawmiO1VeLEMEiGx8AkASVtMPQ+7DgL4N+j99Roy2IX2UlGBriqGufBp1FoCVb9hEI+nxNJsR
iTUxPUHErF9ILhcBJFJJf8HU5RlSI4awh3GNdaN9YXsaVsTOnPX1rsNqbCpAbangg8+cKSjY3QoC
zrtHfq4DG2dd27xHOqzue4g2r7Dk9kSULDTXz25IMT6VrA9GDNILl2WE1uSDpQIyIXQUXBhL4ZIr
8s49OIc+Snf/X3iv2eMsumHpX6iRal4DdczrAoD1rwFkGSwiNXjb0+eTsAD0Abpormf/hQKZLFjR
BQ9lMn7UCm5zwh5b21dv/AQvtrb7j8hqvJq7FCfmDre2cC1NxFLT43MOZJNNGnKWU/qC7Mg3VTDT
7uNXycQa/Cc43RJz+N2/pkmRLbvyaemhX8PMAcAmdD+Aj4jUj3BhRAb+gKiTl66yKaarI3sIi1wa
wVHh8tiC0vkTlALkZ2eXRb4foaz3fZK9TEmqMohXyhFTWAW3MXHYxh6UOB4k2LqF/ZBOtK6bZwyv
yh/jMuEvZ32/vAWvwx+chbVJMF6AP8GknG4FDLXbCNbI75/FwE9hyuLvLiGOG7I/vztTml82t+PT
nYHHNWmN6EPvn8o5E8HXJ6o9HDQBTG3yDZdp7yHfwC1/8yX0sFIJYyk99EqiOGzcs4EH6Mw70TQz
LkIQA8SfvPMYLl5aL4+rjSamEz4GwT3LzjLJCLelFQOeSYYS96WvNhcPtrOaMxB3QaWovajEyKGX
1YxlyRL2A+Sh6sffVaJ3VpNWufq9A5QagqrRbIvzQQ5TQ7BQFLlWAjCklHR/U5y6CnSnPGBbH36I
uGvnQNsVUn719rJCmyFkmkYjyywcHCABJD3Wm2O1NvTRWHsLMesUA5sQRa9nzpyNSCNcgB2mQNQp
b0uL1Ou+Qj921vzi0MmglB2GWieUGZSjup3+oMtxfuIB+hKy1zG6Xr7mrltwzG+T0Fw6C4tNASTs
C3/SQI8VTpYH8hAIWMDUKvz31erOGVUu7Olt/nkPl5VRiKqV7qFflaKgSwHvecp7GT/TYdF/YFfN
2bJdBA3OnicBv+Xk4g5TnoqHuYeVTFfOh+ehWK6AAOAL41hFCXAXB6L5++qg9sFwDzgHf5ihlWK0
lw+xZQc5LeUWK2PAmpLHfypxz76hdC1ygnBkiqu9fL6bcjdpVjZdG82XLwSeIoILtEwyU36Tszu2
Wo0Xmht0Jh317m+h0oSCN+ggkLmEOlgObQn82RRClYzDZLOeVZmm7juz9hql0xIAZbur2JLrerW8
ZcXbYuobVnFic6SvE92+VHxoJ1/x/m2/pDxwWgaL3YpYQ6xzcM6tD2OJyVcymnxd1ikMvTUJiquo
1tpT78Ouw30dJXAW7H2S9I9bASw/Yq0296llFMQlHS9JxoVVzeoM2ejA66xxdVaD/JUupeawvKnq
2Mbgb+GCQo14mH7tplmQYjL2pDGknmQxHFowePXbhjedjRwnTsBt9OEzz3KFpw/6i7aACAUs2bjt
DbN4IdojoRUlnl8zX88KmQDMl716yO+v+4RTF6E5W2kUFysG10VzppieBg+vI/0U/2tp52nYtgPo
NrZdkpxZWQLS1/8vN1TQdNg7aEcRDokpub4eq3lH0xEjiCfvHupV0wzMkYY3Z1Eh4l+J4zvxLH3O
PilnKzgaMKQBxdBxQs626F/xbiWT3wfEj1hU9zG4m5RUcki2CkJYhDL35Cs4Y4pJy29/WHQPU/xL
td+bWqkITnfGHEWWy6uT9Lki3x4ylEXAhmOtiF7o4DovAJ+uktb/BrLMZlw5TeGgS/BMt8h8eYur
f6sr12NQCWrmUI8mscO5OtsOLLoZW+W8Y4UYx6NnN9qlwWxglIdvD0LHl/WBKpNIB2FawjdgcOeE
0Es0bft/3fK96LCfqCQ02O9enJtFPDvrLvAoKO/8o8hCaKhHkqqQbOX6Vfl6Ln4giffF+slppADx
qDAQJdxeWxB0feHXGFz7M+KzzbpHwER+ibLv7MQyjVcLvnjTlbOrJTGod+imAjTClfv+14N9J764
oDAoD1Vs9lAcEMRgLU/+CU4/gEt5+29AxlkVV9Z+OFAuwaziPFhO0gbUmva8PKIN+snxyRP11Qkj
c+n4fLB9ItpqKqolJJfKIMAzu9ZJt1T3DLToVykwFQ+AqSF4v92NzI6UoNsGOm6wytgdruh1bc+r
7ch30rhfqnK3Wtl6Y2qkZqjnEFimShVT2+0Df5883FV0duxZGPvU84sr+yiwRqHxdQJIkiVxt4xl
XIQMUor/tyyAt2QNX/umEn2ztY2iz9yLGQ8Ficew/qwkDkxo6EhlWdnhyTVNyHQ9ITXIFpLwMDQt
Hvq3rznO1xB2RYmT2zaYI7HtYrjDwGJB83jGeYqj0AXSLHjh68DCn+TE3qkZylHkYrg2KPz0pIUa
gLZbU4ca6nhw0OFw3bic1EOlB4J+Pd3LSj6SSJrCzOpEY9Y/zu+lE8Cc5O0tNYNNU9hTm+CynJps
m6XK/b8nvWNfN3EVkxGrfzWpzalIwefmddr3VKEZ29f1XMQ1vjtG+ilz/MCbya7x/0nyqWSKDyFX
fFWOXJ86CBrM+ac6/PrDt+uuJVFghLTS4Oc1FrP0XYXVJjml/sBquFhHs8Ma7tYwt262PYosOrY+
t/FhXV390RQ8lbXCTXKZ1sgbnvPjAjg1PPqkEe4Y88QC+ChWbnXG+Uxv823TYEfVwX99KIWAmMTa
DzcPu3XKyPBnHFjTDDO0/oKcR5YjyQytqpsdXQW7KTgwWf6F1aifEiM6RbD+P7W//4bg88HOqenQ
Z98DmebWXPq9S/niWJjTWfa7JbEvQfMhRAxTbPjX+p4r27JabobaQP0QyA/y25K5u93LZnLvgAD8
G6ceHlNKt8EcmroxHxPNKh1SwGXzTciV7WuxB6cD6jsex6Kl0jj4AlOwulePz3IAMC35R6Mwr6gY
gsFfJ647BZiEwXGyjVIzy2JZGF9J473ZbQ4VxXei8y3NBjMuY/SI3+bGzpPeaVZRsw5/v5TODs1h
vZBFAX0D1/BH5XAUcncsH+IgdZfvkXOu74u34+POnpo3AIdkATuy5hprNGCZPJGHd+LnOuGTY/iG
9+tSOrYsUOzWMaxI7FqoODQDmcBbC9keZBx2T6jzRK6KDIgRMcEAkAZRxdHwguR1Eoi7z308rXEi
7ZFksWgImrD5uto0EyWrwA6id57OfPxPyCm1Bcg3PC86BQUP8iVeD5wuqiVaHUg2ocdjyaf08VcS
05WNchb+Ip7dON1fcUYTD4RBkGkVGLC+BxTxNRWmQfAzA1eEmPJhrOhB8V+J85twdjf+jBlXd0tf
JT2mHhXR8RmHTcYBjkiG7qKlRQnAG7snqtERtyZ1YeXN1eIouBFOJgKTo5FVjCYEMA5f/62x/a4y
jGJS2sfmrQDZqz5V6uJTB49WG/d9TZKc4yJBd1gGbJJYfMJgkXm2OS1Ovm1Pyl1GXEUGq465Egbg
Pu2uvanak5F2ZygKrC7PpRlNBlE7d4T5OHWotqNSQ0eHhSpt6YyLAiWDmB8hq4La2T5zxdx6L0Xu
jHM6q3hU0CgPG4ukiSaKTMbTHaAljcwb9YGP8xErM1e1ltCHgQj34KN6VyfWNSy/MW+r9DvABdGO
+Y6IlWoNo9u7PcC0wQfO2ae2cj34CxGByp6qqLa/Eh4ybGbYdL8dNmaR7pMxht9i6f7nnVrbbEqe
gcZwudcSTuZmkJ34YONLja49dfGtskAhWFFzZ2N7hES2zikthCR5rvuoGmeId32C+OvPKXqtcvsC
lToQ8TeohfV6Sq6JNHMZU58Kb4XQ2ChRqMcBfQ6TRMaSL0Evs2+FaPpeFjOiW2XMuaYMHKnhj9mJ
jni0QrvDm6NZRy3YXJMRw7JI9BvpS2P8R2LPodhgwK4h37H0NWTDqWzs7y9S4VzAyUzn0ccsTGhP
MSdhUfWdbfRj9zwVHEuX3G5//Va8jGJqnWG8vZiBuPjKAIS8Aix+mVxqY3sjgfrZQNQ9Q2DZYPio
07koz1Cx+WOFxMdEPV72mEv37XvsJHqEwnFb8r/ir19CCbt1BtuqQgmI6nDwEuZxak+tFJQfJl9l
yrJ5w94RbCy3QtU9FKAWVqll9C3c8ldWo/bz2K5stfxiNCNdvnTReRBo8z/SQzQ5jRJrJXHVhMgO
KAt0LBifdUZNFScm1LtzlsARccpXIgOsOHSp/AS4KLMA4BUk9resIPbs2XeBKD5+OfscfBO2E/SE
VTK0hRR4yqze4sH713EiYnFww9yprb82B5rtAG1AHAeaHn1G7FRxHfwlSchep5xqtmHSDbtZyws9
90IpZfSfX8T/h1ciieasIBCmxGhQvhNCPiPr49Z6k1/2Sj9KBfIlplAgYyWcNTX5+ILutyeq7a+E
4xOgNmjT761ZqKYWeKhFofsvLOCFlTcpXFyaMka7nPv4j4uWUe7/ghdgjaII1LwgZTwhI/vLJdJZ
zq2v7qOlRe8eOZ2xvltrSqbMzcEkbrBgLYN9Y9+yhYU02JPSihhHEAb/T/9uxB1SrvM74KmywT31
mCPhuxZQX9EHk/xN1klZm0x4KNv1yqQXz1h7b6oGdPKMv+bhIofWuyWWwsF8NR1G0mmq6PCbtgoc
TW6j6/ayj8+PGlliLQl6adqVyGb5DrxTdKIHdKGh/f5/wsZV+OaCCayO8nOSqpnMazGuVZe0Np1u
gP5a4qtEf9lha67TH/mizTNM9y38i43dE9moNQH7U7y0FdJ978SxsMOQXY35E4TN7u4GUoZ+a+NW
M32pd2EQh4r/2BYaRZTqyBTm3pNcnn9CfTCAl/td+lojvTxwl2F4mtTCrkgPEFDjxiiEb0mf98h1
TuJSmFh2ewj8cAG2Nk7XIEEoY7+Pz6Q/LTbtV34Py2h0+sDMw/xwklU0UixKsuVoA4fJa7glIG3E
0bvoRT76lOUJNHCYz4vOdwApCOdYs4jzJ4U6hADMcAwE9dVT20kuK41sLfi/VOO9m5Y+kn+bMM8V
KOF6VgMmZfDhn9iOnuSdHXxhE/62FMk42Tjd3e9cc7Oe2QwIL9PMpjdy+x+Jz89qtXkdDfZEjbkg
rRCXYeSJS7M06TKrBmJ0oPt7P3OIHxELT4XcqI6ouzWqSR33ai+yDSOFG+qCKcGcgQAsHRaZ1Gh/
ZK+0A+wQ9uC0kJHuRx3ABqvoZkNHm/0KIjmk5N0Md9mghDN+4HEiLLJWoK+/FUn4J2VEtiek3dqg
QX0h0iUtiMFDqycOoX7VwjgOBSYN1CuLi/8CNPyLW4wcf23mcpDkl5N5I5FiCV9efDFWgmav4RnO
vDubYZrYiri33GjB4Sy4qmH0wrmv3uuEAaidIe6i2LOSb0ytdoGqbEI2iUjsDAIdlXYyxpL0rDm8
rBz816ME53JHurItoXDnJRkAqgs9OAUiEQ9g8OZgyDELNRdwWieE6OF6AKB/DngMmSEt/N4MlmVx
rCPvTUxIMxC+9+KoA6De8+ajOjm14JyNWHfACYL8y2+35quLZ4dBBqdcqErIKnvG5RofM7AOE91F
+Vp9Z1oSivOfXNLTHd0Vxm9D4F6x96HdTGOKLlSp6XFCCFfpLvyzRTYWMAimYa6HNMoN4SwoAw+R
mIG2J3QppCV34leCsDjGrRsAciZxAq8ke4k1lfUJqFf9tqdh3hYvlNshq2yfF5RaIgiCg4PBpclw
xQjf4vlY5oZ4/V47usW8wHz+1ECVJALMC1YodJq2ZAno5pTuo53XJVRMTLnQW6M1xF6nv74ZKVUS
TfdJiE5g3knZ3xCveVjSlFsj9Yi5pJmtE3AZb0PMD1fOBw7wUM2/GU4pj6ovVfpM+irhS1inLuM2
tr4Z9XZEfI+pN2g1mMrXIQajLbRoiG0S1Y2A5H8F5hVIaLgi8yFwh9BD93psBVOSv1ZL5EX1h8kP
d2Q4cKgWnXXS6MM3w06MpUAJVn0h8Az1ifiBmzX0VjSkXZRffoDfGVkjCGRo5gmb9QwORBKvphqw
5ovcZOjTnLNF1Bd6VH0zQj2coiHXCJAXiXlKuwlRjEheRAYXlpNVMIJJoZWgtr1pCJTuEWaXs0Sa
hCbmWHp+AkS+Ra7A78qx1aBYxZIulyOZOg29M7VY20sjeC+xvR4OZj3onVYAJjwmeABLbgYheHMm
Qz4Y9XbJ2GPtmvoS1oKj0CeV8jLfHcSjJekURCS4Ht7P4fK4NJs8qy9KPGzKHVfe41EHogbto+vp
5FxiExvS3S5NG4gDHXY4QniUNtBGRtWgDyiHLcqoeIcxVuKH1Y9Ntn3o0L7Vhh2ChXJhz6GineUy
uVCZ+dSi11NxXL3I1jo6T7Jq8B7IblNvjEOxOUduAcqLGLyEuVPLVmRYXuREElrZLAwojK31stWY
rIjXaxgcs9UV0sSfkTa6lOfdIuAdcCMB/Ag8VUCInJRGEwubp44oFwDukknGhoqOwUc1AzaJF8zj
/qex+GDMGWG0ewZ+Ma6Iolq5Pk+EuPXLVKqiBMQ2zxgSe5mTb4hyhR7b8GltL3fBlKftkL/JQKs0
ecc93NclpKO224PKR9uZAEo4P7ciAylG+SMZdD3fr7Y1180axyH36ILvE9BsxG+3DMw/Tc/Ux9de
LKUPo17W64CdlLxU46fO4k/WJ0zRM6pvHO90rvPaqcdOP1zfxTgNeov/2DHZ9TbTBmCPpw8wjiw7
9e0lUpMn2IPtYscAxj5GSsUPaHrD4vlp1wXkqhUYNL5bMTm3cDNeJL8wdyFJDegy2Mrat3NfWZbZ
9CTSwhNifxeQwsxzr/HSzItpStxt64W/LZccI8IbqiO8XnjKSRAfbrNcZ6GleVUyz5xloTHhJZle
HLZh5XfYrufSGQroABQiDtNuqWabAL2i0bH+lRHyeiTLd5v45r+lyN6QdsRqJQCgFagcxXoKwTI2
R+fhXz1F/iaYpMDCPnPbQJkKhVoDPO3Z9fwAg9pa1l0B9vXQ/541sFh17foEHxEtezVBQs868bcu
oZQ70NsvpoQRlgCBiRgrFc5ZqVvSnPTWmH1D6x3g/NIqyxSMJ6WEsNhkKvocoYDL03xSn0r2vVB/
j4412d+n2JouaGjOEXZm7X0Wnp+hTNU1CXWRPHECNS8c1kPreWh2EWJ26usiMNpPuEf/7zVlfGgB
zE/KSJ2KjXQ1P09kb4fUUqL3tCynA9wivhwbrJYriorJdgewpzKXGiyXYTf/F9jAGLEHXuMmdTcI
oLzAWr7UPr04As5JrzZrL/bczuOp4mZArtVW4mF2EsWUBz8rQx2DS8nAp2kn9cKZAAqGp7gWiU1N
WYZ0jygqvCDDVnGFNZNS6NRiHiF/8cQxpdOpnY4Q5SYIPrVPF96AhYi6AjDZc2WJpGk5vknWCBNl
3y9ze16WjSqE5fOOlg1muMbX7jrmd/cXK7AMAUi8IsBvaikkAvIu+MD6LlXeUOMFydgNvHy4zOm2
lf7JtYlO/bcVIo4EX7EatCEo/PlNVYN8d0XqZM3GHxIN7O4w6xxQC+Vs8cPLXzRy3YitCJmaf55h
x9L4bhjDwR3kYtWDpRdGLW8FsPJvZkS+67CPUpgeGE+v48LhsPPzqyq7I5CMIj+L6gXSmruaygqx
RPvBWVC3db4XzcoKtEnYnHdQ+CDlF+2A7IFR5EWqd6FnFor2djVzWEKoCa/kzDHjf9kWyvP6NhVQ
mHuSFRjytlwxaz7RONwlGP4fsLePddVXKjdqFk+2kyySMptHkzxPpsB3x6VE8AVb2emYfgRw8+Jx
BH4MuaMOejcLlRTYLyhAw0wLdF9t7zLHFoe4GP5cEQpZJAEm2KanxA6cz5MNHZsnKOt1PC3ae1wp
Vt9Qeeg/+Tqx2uc3qshaNsc/R7C19wGbyJx/cnOE/PTHXihL4MKHfMZYUe6xgSQn0kb4xzJkMrV2
+TkQh1PrrNlJkrsavfcuCk8iCFVzOL2wcD/sdFo2ucU8ldDCfDTTFXaO8IsvmN3qybNfx5paEGJW
iks26Mej/5IVY4Xt0OKRPWubTdmtomO3yrCTzGcmlJQl0slPUxVV8TrNXs0Q6xRSrwnY20OS5dNS
441nyeeE3j9uXwkgH3pPNCaItC/SRDcoGjsqS/lB7wVHv+hiFI/CUgnkvkgHscvOyXrjStYpSkop
y7bQYk4syhv7n4qu7y2w9fIVz44ZbxPVIxjYnOkC5YlUaqMIsqDSX3fS6PITXTJXzMyeUUQhHGcd
WX7neCLxXxL2h4IvjYpWj/dLr8Fr9ZFZzezH7bykftdeUxgy5GguhwPELWfdSr0wxqb0Vv2UAJOh
1dc11s9nbRvibruG/xrF4hoi5MPBkBsrtuUqBJyWvsCgeZpk+k4ionxd5rul8r2dGPEj3QQq/1u9
MeUltDYTx3XXvr/VLg8MDILdX2KA+ssGpSjNdgFG1ZXYFNSxR+v0NAgMhe0Z3DRmcLO0L5QL+iz5
C6fPZ/zsTjqjbq6u9F+2bFEKAQmbGhzXIe6DeLTY+rB9yz4qooYYnNqSX5fqUJQw2rKfYQNuxxZb
nP6HmWBRe5xyTZi/f0Pj3PV6mnb8JBXznLzhv1b+VSui2YocR9ZQxIvJQlz700FM1P6ST5kJPMTL
naKwNA0NcK2zXiSIG/lQC8TSCVe/44puK3XJC5C+rAxEvPJQmvk2tVTAw7ECg0t1WOWNK5irB+0X
Jno7mstJyByQo68WIIko+ZJEh9p93dOTQhOCOfWPsgIfrHAqg6RvzWDszyKYw3riUgUVSh5ly2OT
mx8JTsEQK19JKJrWq/uhXQ6jH4wqIMrgoYQxeUaXxGiBDVnn4+2Y+RzRNG7L+F/GffoM57xgwSML
7Gr79sDdoxl4OjUDif7M3aQgZmUL8w/DOepHDoLEzkpk9nq+CZGSoQEGL9ZVwBgydLitFjmssmn/
RpQwYaz3bUU4TBnemMlmomDnUbDl/43O1SnZHWvFkABY4/oP3rBXz+oWK6v0NkrdWP+pG5rwXKRP
76egfggGhu5O8BkYUV70s9bpDhnj5kfOcdb0IsUs8EgbCGmuPEX7gxnthYfbiFA6O7s4igbHaWJJ
B4BiJBcsEevhCJ9tqaiHxAa4h/WwSrCVmWzbyUkZCSLjbT23W85cLDIpZV5XDYhN0sbJlLIKmkeb
+DujsB2MMBPUTGXFAzGk40UAAMU02pbyh/Il97ZoZeiEn9qRD1gs7SiPSPVQWxt1iERg5Z7LPZE2
ttrpbIUPCLsUNWhLdUcw9O3XxtetIvOSxOnbZhyHAWR1+ZR7RnekPq5ewxISzsmzp33eURl5b1Uk
B/KdP282ywMbC/Z7rQKjiJs+q/7h1Eqy9u8cxm4si0BF1HqKZHGhW+oqxradNBdiUwG9IoF3+68R
NLk4VRjSdg++OCZ28PIyaooDzzQdUKezj/jfJukKEziXO+JfwqqGZRQ4j8xpHK0QSU7nRvgGYWij
XzD/M6NXlXQkUCmzjOB5WdGNwUEschiPSNFqVO6hKQleVOrX7B+Rs4dUEtn9m0qsD4MjC8hIghBI
c/5erI/6qC9ARsnu9jMvIoFKSwMer0KzJj3g+eWVkOwqXzggF9kmk0OSoExD7qs9EvMCKXBb32TC
jjqmUxqfX6wOkYkF+sCQ4oY9Wm7soi+yGXY8549tKtvwQ7S6OR71xvtTyNP+JF/F6fLt6NUcn+Jh
232rwHxMVi79m47XJ3k0a/Nd5qQqStH9l863fy+LMW5zfBGOJCNsik7SFttlAide5dBycdcRiKR3
UxQ1dh4Pm+WSM1T3sO79By6XnoD5joQLXggRsz9vuhv9hFcfeglYttPlD/bRz8qTL1Lb3tHs7AOa
v/UUa4/h10iv1QN/RXNmryAZNu7XgjhS0VsYrAcXLN29m7di98SAGHV0HkL0CgukYCwoe4NdlBtp
W8TvHhrX0AlaDj4KAFG4GaZH2YZN1buQQjxjEbravYHV/lOvK/MASVi9nF9AkLDcpfUwfpDYMSZx
1sPpm0uq0g6EiI+nTT1XK06bR4vBFretjr+XIjwKF/RMl18WUfLKZ/vhXP5/VoUhXQnug5HsyFBa
NtjY/MHMOhu4wxpij/DapatEvROfcvbXYglt93mgntwv3PbcQ2uprJPwPeTRWCuyzWjbVo8hxJku
p55jaV7eFK56zxeVuN+3yMLsFjVBpdXKLe4W8GEk04IrxFEgNktoYX/XN8OTxRSSDCk7o2cTqK2K
CpVIWmMrElyaBZvxLJp+GlYwar+pWxiWH/9H946alGXLnwC1NCorS+ObSlyERc2p036vF/wnjjHt
AUSIpxRkj9+DKjd6+BrsTOuDnh+hNEgus2dsWRed3ACHITZle+okENu2xZscSIHzNqXkEYOTH+bW
ESVyyaiYSPSRzPccp898GDZHtHTR4VfWNT931Qw/W/ZibKzVqz8zt//Hc4kmo7BNU0BxE7842Hr+
WyyjJfPpKQ0HuetONhg2Njo7V1EdQrSALJ9UHqMFyp0Xe91Um/gltkOX7oGVMcPMD6ULdNTtSSjh
Xnm7DC8PwkkOfxCOkrQrg5apzI0pIKw+L5dIWp7mkqkHQRa7DA3FsWyVw+HEj3kHBwjpCKkAOoCa
qaIAqGdnD+pLTog+AUWY/oLLxq29RVAOPx/jQZNchMh0hilHajim8e0lFzyJ8ds1Y2KwkVO82uP7
bxBEEJS6RTtaAgLknrFlVXHMiVZy0uos1b/ecBEP/45ADKJ/qiPl40QURBvUKMhgT03oRANCuu5X
oNcQ7sfYR6An2Ixsoq1BR7pDSTEo08nElF93C5tiqq6uCtQPnLqBOwUsSJABTiWSsaD7O1bjKXZi
cZ7gXe8K5B9/S2ME/dNtFzJI1MjD3BzM07IX0pRn3caG4anLl59AkN1YttR/v5RuDxXjVfcgLpCI
g1llpaUCojyMrPehqKlXmgUdjqrKV0meForOwtSmR9NkJjuUfUdZA3PMsuFPpUwEACisAaw9Fpyy
/uAn2uUlablDgYg8cEJTSU8xHX5Gsj3YpgPGh1ZnjddbVQZOYkQVEWSQG8dcbOc9fZitu2+3QfqD
OX0PfyHhr8TveCGcFTuMde+HrSBrl79OqfSdbWGzPrgHyjfSCejKr1W298/z0HjOW3DLkSKmZ7Jp
N2LPN9wbiRxVchkISQ4rhVtkySJwyAdnbEkIIPPRMHz/6nQLs5rVC6TT8Nz13fU7b2bfFfd6rm5S
LUXFfx/O1Phy4NMDHDpf6tiPysbzSKH5da9K2FxTF23vsBx+m48RoZWpxFY7rkzcWnaoO9H71i/N
sisz2pGUxb1JPI6IKt6C4GjpjTgZ90u1iAUIpq15ycChhSfsc4YdcQgMuPi8Hpm7y3JW2GhNzRM1
NYUJO+d4I0IPtBRxGt6ACZ+msZneUW1eziFzajgrST+g+SUresaZj/DtQ1UoL8DawL8zcmGMMeqE
BxBB0I7TkkpQ5VBIg6fBr7TamjJrgkSeEY8NSQ3SSO1+6xYTZMFHNjpJDf1V+4WHP74PmR+QYZ5h
Hzlyn3iCVXH1uGV8ZQNnqDv22GVC6TPnmBmBNPkQQawyZ13/DELQLiVwbyzWZcryO7oYELFoiXNp
ernOnjo0QeBKgHt7e6bKc7of9mv/XdIxZk1qtwqCHnVocXdtBti4OD8Xi4YO/ddbxBZXCv7dHA08
KAOj6mEOz3ZGRwXcalmh48yw+txQC6vwCwjaK3FyTZiyuhsljd5ocOoq4429Wa9jVEa5vBHfWpma
7DCsK2hpHpTH+q52C1FFhFFGcX5crO3g7KYE2SoqZ+d+kSiJyLjj7+wfWhX6PsdRY2lImvzVWiOy
mamntIm8VLKozpvMhB29TrB62sgcQrprlPCZdsa5bbDTnVcbrpNqx8WwzkSITTKWpuNGv+V8wnF9
3Y/4dOLNrWDOT3o8xS3FazuOJ+aYlNSJtRKrHVELSwIz3Li8kKZEaSx6vFUW4KwKzSBC2VgQOp55
DzexwJkFXui2vlV9VIcqhIg50VeIJ8qpS40uH2pZy2uMN7xL5o/uuoFatGE1r1jMQSR/OTy5Rzqe
BKDnQQX0bGZJWbOuwETsxSnLu6IJG9h4MdVrM18oUn4CP3awoiN/7atEuMHVO3VTMNn63gRhT3Ah
Hav0TU1ebob8Xq0SwMJUUMAW6dLwKGlw174Obia63/kfOe9eNbRXZhbVcRf6aencX9kzYUtZY7e6
5VXESFAs34tD93ciwmZfdCDXKITrN8OhSL2V7Es1xPt6Co6+VrcYOlC2gebFFD3dr3CJVTyPmsep
I18ncY00xmsdLVZF7zl2bBo/aWT6ztptrAfKcy2ooTFR2o3jzU5uhuOXYMyyRvqqJ/oMF527bu4I
3y0ofeGQOzO7Q/vKsbbOY7YgiemDcM+QpTNK7fW++NRNNSv+LkNb1Rlt0S2pJa8XS3suIZUVeaV2
QUsLP7n/fT4KWsleC5QQReGueVmPSqMxKcSfYejubNZzhUDXUo8DTQwHYplCIb5tmHyq2rr/D4SM
UrpwD15F/yCwAiIE+fprHzYW4hXVm/0uIf+qvJHO91f01M/0ILSmxQthGc+ojM9lmA3vlVo8xx4S
hNa/kb7BQ6gBGH0AbBqFdIpVVYm1h9e+/Ce03onSPyuCh8/kS6QdTfdOG3VKgVMstP9Ui34qa4Ro
Dhi8WWOhBRyQN+m1CxUySqvCqKke03eCOaQBZDLg6Z+zv6K/wiD3p98suj+o1Tara4r6yJ5ef3yC
C3pqvXYtSpZ6/R0RnW/KcFE+LEknYoKQli6plCuWp2Xz27J+GVionFCBlbtRgYPt0OCo98A12ZuV
krjUwK0NGOdzDNd0dWJQDmVNQke2Y6VDPVEnVq6viadPNvFSpS95KvOnDSVN0a7eUpJds6ZXt7QA
hBiM7BxpkLgyykJD+oFeTXC3nwQAtyWhN+TISossnsGLz2kr/pGQvv2EwbF4dTqdMokKrviik0hV
YzMKcxwiY62A8hBKDJf6AOCt8I1BUaZz6wPjZGiuwevF5jS6ucBx0akEBTMXTM+qlrgl0yNIcavE
YQG+DtGoPx6lr+F7L7eSD48OFmCaA1O61qLEU93RoR4/sxBoxjZQMEV95/pYyIb3Ji6tFCTd4IW1
m8M/PN6Ydnk2gUp87A6Xfvi5Zoq7PWfjWTzmoX+1GL/iiMgEz2ABzkgmg7rJa3ZUF7YYZ08JFzVK
RUyUeopQk13pkrLXscQZQXvm5jFMFSuM6s37DG/QPxZb9h1UT/k2PVCV9XeGd9pv/v1njZV6Uxlz
EyexOopXgN6Q41DRyDAtHGrQ6jCCrz76JRUZYRKqSF2eru8keTPN/VV0l6ioPgzSa5HBbUOSx04O
4XraavIdAJSKrMp8VArwoP84qiwoMx+Kmf1wPCN4OTczTeuYvjCD4+A9tNwjHvR+MbqpSKVtR+kJ
CdXPQgREtOMhdKxjW8GhOb0s7xnwBwmdUfdoVQY8FhHfvMn541C+KRwFsz6PlJABrJTVcXVJ6GA8
/g1BgpqiRFMfOPVyGyMYgDgpauacmGh4nTHqkkKsiBog9LQ73TSG2zckq08LeE/w0JC2lmu6pThh
kNjFNJ+a67WeCWnVcd9A2ywa8OKYNx+JIikP1ZioWHTfmj/htDxjr/Hfgb5UGvHv6rXNbr4+oVHC
QRorXUnX2tYSngXCCYMV/lS4nYTg69nPrReabffbPe5o1lZav818KJWokG3N74f4tSLAr9LvMIoe
zYum14I7jV6N1KdZaRKmlZR4bYFEu7ms1xL1cr07qdXl0324bM97lwfgDGXQFly6GJWydPhcxwjy
NJI0oiOCKI21VqCm/2TifZA1YIGkuU+yiLNYl++RE6kEAq6cEqlss0Y6USah+S/BGaN33OuWI4/3
4hTRKI/TVZpH/1304VcAEH0Z8FcwB7F1lADGjwwo0icAj2CyVGVQS9xjglBkurtNVQ1iilh/BLK9
npB0dOeoY+pggFbxjmeY5ftgJKwMCh2z6F6cr04fgP8zqUXtSWE7X02XVv1Ivf8rFn4DshWSVKWu
IpZDa3uaX6To54bT/tDTMi00QAullowIzATuTM6dqk/BpG+C2sv6J8psvJxznOktb8u5pRXHqSB6
j/CzFZKOUFz6Wf4z/UOrMR4RWVP4OIhW1APCwKyMynmMrXq1m1T0u6dd4e2nLuW6VSOMkgIfx5b2
YTwGrhWKZTmR6NNFe4hxGPhOy/YuxCDS9YQSs37URKLXjVL6GCQt5l6GpTecCXFNZgZYtayeC0ro
1x02bhwYPjXpeaVURk2NtU8/x1lx9kta9D1bC3+w2Y+4LYhee1JLFXey4vwdl+kXjZxAh8NE5VTB
ENVs2qmEqLSHpAj5YAKT64P8ISKmxCI41ofmiNMD+rZ4x5ZSXBaKNJhnxbHFBY6mPH2neDUXlZAR
gB0KvtWaMPmGJXg5a6nH1a8vteeInoOsMoLgYjnTlrwA4PzvPFzmpjtyk1IxQYeXKQWmZ+1C9pf8
RNmx0QKjwe5VJjwcNypZIGuGX/VHOIq5dI0t9oUT9UKUZ8cKV0OWBAJTroCPQnD93oWtHm+eRxFR
dlj2zNXXWS7nr1bbLwbfFZA0L2d8njwuJ02tLRnEY5c527aauzCkaDVDNfdHQP6Zt2PT+FOYb/7D
akfgs6Uc2NtZc0jLgb4ShcCNG8G6sMLx21yw9YxOyaqF7uXfvgXuTwwbFohhkZauFDN33UHSYuhc
2mw4CuhsO74DN9xzBR0jaT6PI0UZOSq06xnZ3Gf9GAZjiz98gmb8YQt/Ekb7sa9vkBx7JCJPhjOb
zymUNoLnta0zYoZPkmNUlX1aNMm3hHHCm/WWSLw2Ml98rMIyHy6Xja1z4kj3a3L/HPKmV+cnac8s
Xwg4+2ZCw8sa5lvrdCm9WRPePhVN3CvFZSCvcjqfti4yarXXqiB5mEQNe1ZPw/hwfTCFK2H9CGNP
ILps+lG86Kyxqh1X49lS2v607cigrtbUUc9jEkT/qm4u3hvw7/WE8jKZf+NWkV/KPzuIG3LTnNEd
iOvgo2JMWTCpI1q+JWTljzMv1OW8BoQo0mcK7RAcKY7pEhX7J0dQ/r1jqtDSzUoSw2+38mrVopYd
QkRz0hglXtOhUK1VLu69kqb6zoMAzIVIG/iZRVh7fTTs/cTxkGS/jtTDlaIDVGfo1TmQ4PbUIXoB
FY/SkUvltEUWxSAQzdUNzB3w1wW0LCtkesbIHfObOqZRjNu3k9cnv7yBhJT70HVOhqHVFYXyXCBb
ufKlGGFNCt2dnvylWi3hwMHCKM3sRE0BmhgmdiKq77ukfjs2gzjhIED9xUmcm2e/hsiAesJ1mVZD
ZhRqpHpx1zgemzGv0bk3egWLqpaqvu/R5DgGs1l965bUR8TzYnB9JyeoErlu3WTMioDvrNr/MIi5
rNrc59/GoDDNX5eiZRcEaO7jocNmS7pKgAF2G+h6proi+iO+I4aQX9PHy8J3x7cmNuqMMch2LjoC
ar2AdauqRVMwtyssvtQ9jUN0HftSmQDHTHckip3awM8KE0CpS3Dy5MNXFUC1GRotIxiCnQ7bQwTw
5h/XfWT3M/Yx4RgZa06Ub4wJxfomWSD5UW6K2YMlKmMpCkOYXEP4Rzn+RnEdcXtDKUVD+Vjjwwco
8SmU1Dwcy3FNLu4VueGRWPuKwkY9Kl44lgH4ZG5u7M4rL4JsUg6AKTDtI6x/osXcgLB7SCB36GAs
rFUSTBqgrwqIzPv5+jcH60VP/y6yb1r/XEVFUZ+KXFru9LiVjNa+WQ8/N65JuyOB/Ktjhf5Jph0Y
sqqlyD+QJhSP1Ss6ljpq/1ujLyYoy9CcFIyqRNuiLvPbhv3triTspC/KdFYlT0TKx2bsXW3zwBbc
2fTtubZ0E1KR5vOA56Wnp34cmXMTk4KVPnXlX47C7m5j0hv6X7tJp/kJsGR6LAzMAcJDigIdKk82
7VxSG/XBvL1Ti6qtXr8h1eh/cXvO8oMCIXcSbD6qvcgvNM1/H96m36geH+VJyeIK6mjvOJTEpYmp
PHL/pRbZufMCb1rbg5x/LPj97JBo1v35+zpnKLcoEGXtEi2aGtK4YEuJ0eTirdiuGo4rUJKoKx4l
l3YdqH4edZ0vRqDahcQZeXkz4yucEKc3Dbaq9UMhcYcYIVQRNMrYrwfd2hKIiw+8VvzQ7aM3K1Hr
cddTt1moBmbGSJpWZsUHnTKgruVUIjFYd5eelaED7tS23MY+eama3FkL01+6z9U5gaQlh023gFzf
Slt6k7nDVevHE9u4Fzu2XPLjmq0PI71mJI+pxx9MNokIxu63iK+QaEgcUk+vjJGfvyfkKIGxLJD8
8HwG68O9t3ays1v2IGBnUAgXhjwLBt6Oe5qT+YTxrw8t4QlLzaYfMu7uaMZTwuE2SLJI33zzrFw6
AaCzvEzs+PTmJ5OEhSbA1wEP+o1Pgi5eoXTIh6RQT/cHj97o1nj28zPPLunPY7M0XX/L5Je2QhLZ
fgHxHaa8hZRhbrlwy0rZyWxc/FoUCJjxihsbXsKsnfYhHCdcuPKqRT/6VscUhwImYCC7YvPYCQN8
TV8yOOWK/R28Iq58ctvEE8AghvYr/K6AwobVKCk/H/inoSrboxOzPc/hLDql5Qpa1MWeiuOK0umL
jgbhgKvg5jDotMkkRmTgV8DH8yHAvQeLfVmFDnWVXaI7xQTmzWzCKsy8nLS7tCpNROVJTFdaK8X/
fvs3r2Qf16ski1g98cgU3vaVFLBRLdcw/X8kU4GEzhMPLVCeMOsvZZE444fiJuBypwUhO++TW1Wy
vEB5jfe+uej0ne8BaOdQjtaQ9Hk/D4sKxHzK3jdpCA0+zOxQOn7sfbhV+CNC2qk8ZtRr/Rew+UuD
a8fOBK6zOiSb/7y24ggvDZYbDBZowiPvXaWb8ztpgdWMR6x0xB3dgLpxyjyiabfceX6Ye6icrNTg
NCQEtHQWf6zoupXOXbwSi7nhDlQdCaiwJIPIm34dRAYfk29vfpEHEOjNhrrQJ9lw4GD17daQ5hWW
w7Pz6a2o0qvAkFjYDPzKe8SSe1/fdX3qh6iMhjH2y+WB7Fkjbd4cxPlSZQRFJxkugclle6l4q4hu
T0ORXWgwchMUL5UHfUDy1zQauDlDzOtD18ugAmIrHk0Ym9szGO/8Yp8XTfNHoiIGBB9uV84I4VVe
PlcM+tlU7OdPwVOzvRK8s8rOZS8J1wi+ruenscNwWkQBB/L/yYLNywXRX5BdlbpQ2VlXb8xtGx7H
lBhtSgJOXZsPy7mmw+L7eGKmeLxxbk5tMvVY7XhjsZf5siDGD2nNRUzYNVFvtMvCUXQ4ypMW6YMb
iuN6kETgqUptwtuvvbz/IiF+5WbIi+TMWVPqQ8ZMi4K9XRaelpzR99CZEkdRT3RZem9Q9TpiSIPO
3ufj5+gvjqxYVl2lbV4zzmE1VSvKeOVL+vlcXb9WCtUIH1/AIw49t8nGVitPJRCk+TMExEZ78hSv
8YQM7AYPGI9NGg8taHtd+aNBL0Ivuxvx+Ro7TujH44tOAiXkeJnKC5TU+bZyi8SvVUbn5Hu5UHV2
D7j6Q7wLJCz707cPT9oXfgcj5CQUxNCABRLC5CW+rFcbs3QfzPy63iXiwA/uim80Zrbo+UCdtlH3
RdGUoy6FzWE9JkeVwn2/iomZQjCP3+zHXoYCp6Ar5ocWey9cuxlLfP9FbMKcYjzWS509A7NsHc3l
o0910/1okSw/B7KzzsylhhpMR8pc/h0zFoO4crMyJ738sDmSyZAsya0/+oqHPX1kg+1YjKLPymxB
QRHI7VAwGXOvvKnY6wJeC9K2kcWhuCXAQ6e/bD4riRZkjjJN8K2B3UfAvwYRZBTQFgFrSk3wNqe/
aHbiIkT5wrG/UFYJnLynajvgyhlMhF0/7w7Nb/DVg395ofXJQoDKRpjskXGDffzvLLm8ptyZpDW9
iSxYsMzRZd2ozJ1Mr3JmFCmZMk0l7VximZXtw/0l844k3DST1NYlV5ja1NnzOjYqnGDGudNXC0WO
BUYoPb3C8yIf8bRK6L7RjwZ0+4vTeE8qzEvMNkEOL2um6nITWMe1TB4Ryv2ijoo+jAHJEAPGfxBg
+zn0RlMcCeEf3O17garis5R4N3BzgSnldbfCsUlpjyInTSpZ5o/FWwVk5I+EQ5YE694jTNAPEyY8
LSGyPAjp+71dzAS8NxB4Q3R0R8n8oAjuCueoX0WTc0Q7egpBoQpMRBvyDZpDaIZF/kd0JuT0qGJp
L9+QvuggzB+W5z2I20GeHkioAiJ9EaPYfdE08RzUaKs+yRAbyh+fu1RaHClb6FrIDi90J8ONHe1F
U3ivYPYFZMrDMo5anaFtNEdPN84EajL4sd8TdribqYNxOkRvwBQNHYBxHzDot9WwEOvLtvuvHLOZ
35arNlyp7IYas27sV2h3e6bYg18o70C0h9FM4byX6/hMGoVdkVihUsu/MF0DXVwcS7CvuqKfGwWN
bl7PdgroIDRByVnTh3mFji4kWPFA4npLXDC5Mg5cLB4R5L+jNy92gCCRVxvl9PnBbS5XF+wRJl7u
taqSRdTNoFA8/+nIO41E3SBfcnxeCs2i/4TrHjGMGBW6hYh5E6GhqO4nrYoXsecYjoVRchvfwrQI
iConD9Bl4gBU/539NgjJjdniAkn9oHGcCC7HgDvJtQbFXRR03OO6FFj7QTEuqtL7dUsdRPV1cpf+
6jZDRQj/lLzCQLL/HdBM+HJ8Hh4CE1xHhMbHimCF1jjwIyDfuz21OUtI6wEYJm7zjeIW+5+txC82
BA7tGOAHobpMt0cXQGoaqRq9nnYZ7nCHCnRbTiTUp9pyvEsJai4r0HwkxjxR0uUMiSO2l2gLeR6/
G20btKD9yrb/P1KAPmpy2j0J0VuwDXuxkkrdkEEPM3buGOgv9E2tTKvRl3U97qqJJ8duxlVMG114
wdlEIthlzPcrTTvcZsi+ml8rD8/inWl3cNMliLQHBtGLniKx2cmsAgqIAAPowuPonTtMjUxGP3EJ
sVGdBAyTw9QfB6jlZ7jJGloyqWEJvtjDmnofJN/tZXRJH5ro9/jlfkoZ4Scz/BFrQD528f0L6YSW
pc3WNtdczqm7GS7jkHBpLzPzFE8J9nMw5w+o0ZecRhv30Cd/9PW7n3GQclWpSgUhb2kWmb+iLDYf
V9Lqc9jWk6gCadHls8M5XtdkA0xbU5dUihM9S7Bx6Mq+CjdmuOoqQkMA7hD0Or4OgvHiXlFoPCl/
rQJ08cuY4rJyV5iRLWIBpKG+eXbBXOTl8U+J0reqltj3cZPEthmS+FG741zfGTCfccsOJo0bzfiI
nDb4Nfy7UjX1RElYqEgwUkrb+1ijcgOLK4pckd0ognsjuZWs2gdanzkn1watLilCPYWv8kympo+F
8e7l3QGA/8IV3xSV4X/2gssp6eB3zI7JJWdBG7prOE2H2QrF6K4jaVDUey8jN3PmkUaphkTIMmeY
j6ucXGc2yiwKts+5yfSgUKpdTMzyvmhfVD9TP9jtZT2QyR0xeClRJaWjRg3NE3b6o6mAB8CZCPWc
NETfPS+M9ilaIHxxsw6OmVrZalEtqtfTXwtJvtX3cHJrZdBp7pfHJf9nhUJc/GYGeOmOXsa2pZq4
1N/ABqyWrvFTVqGEJEU3z3bW5xeh3Xnsvw3YOYWpsJ2QgoJRi3VI3MQEQy1CKQQIJHQUJUfugSDx
kxri67mfBlJHpJzzNdFmZjFkTAC54fkydPt+o7T3KIh3rL6rMxrFy/IQanDeV66gYlAPnMyWcnTz
lSMz9WFOapJ3UNQz9qlYuqB3MhEWDo8Uf8j6PSz3VW+QqQaGl4HMo4+Ye78bA0bE5obZnNOd1vjW
A0RpNHrwamDXLWQhC/hdQtiRYJDZGBYfW4fDRBUrb9GD2ttGrBXIKqCNZXis8dsNrh6TspigTA4P
xpTMJ5nhrTYaRQReZKlRp2AMGG0j3FwnPYyNkH9Qca5zEV+TohQiYTQnaZhfuKBM3ZCYOrYpebux
qgFHRdkjnh7sbvuGF5LC7h5eZ3blKw44OH8zi2J4r5ZBezwKRbXQVlS3zTnGEHYVXxkhiX47hGie
CO3HipUM8PnEWrDhw//RIbFYikyc050fTpgilPtR5JP/eJGQQ0Fp1+kTl4VR/Kk0oR5h7kT1+AMJ
AqVuV1gSBLQy68vWJA9lvJ69EBwQ05OVnKTkAbqJ3QWpHnVc6XuCv90izTON3rmKGMCHVMKo2yZ0
OpDvM/rnMw3ecSXCP6ZDobNLEMEJTs1S+l9/+Pvui6TEcNPvTCa8dbWYC2NgAxdVN42Xf2uNLelL
2zKZkE9ol5p7lyZf/fxkq1ns+em6JDGQvWg3Xn7/jiemPr8L+MQX4YW5WGUbRJMHZPs7J1GPmgfO
uldrjEO+Mk13yD87cRJyEx0tK3wCj/95CKdej6SJx+wDeJ7lSDfEIDcRIyfiMMwajELAyKnm+Ci9
+aaHA0q4B2EuPgw+Og/hnfLh1nwzYGpGZQlgc4DqYQV8xiRbA16NumG7UqkS859jGpcJZr4E/o9S
1UGjOh3ca/QchLTrTaYHI7YYRZUG7kVuT4LBUVrrdQ1TN60l59sqJzKG+wDpR/qJRl4R5SeiXYZH
uhUkc58nRq7aBa9CMnWWoDAoVz8GJGlYdbX6d7oyDdpUS8FpYurcijr9zkxVEwvJjQJpy2JUkDV+
7bkgitaJEZz5kIU6VXJvB3cioUF62wSRv8fOp5htdYrjWcPEuBVRnXNoIPt7rGsonPn2hMDN+/7H
kugAEmssZNzXCn3IE8eikGzhQVGHcDvhcmhhQrWybBCaXg8zBI+PoJ+2UZKMliEmWX2XUB0hq9UM
hwkwZ0pYkAhkt4d/OQcbeZhq1bdc6wTRp8N86Afu+TjCjGTk3+Zn9lBImDLGx3+prW0BLxKVR3eX
wIllGCR5/UVaKVkoJicjKFOh8AbCIZLsLyglboiSrAmckCuIu6TspNMtTfk9VkJlScX/dgsMOCBJ
Pn2m7nzeutIqIssWxxp97kak2ka3Flil2+9PaeFBQTQNNSmv2iNUCOJO0TgjcJwPgeuMxZczT+gJ
ziDMJWHO6OArVmTuWaSjCIaOTd4i//ll/6MKHWmnqF6wrLXfWWsouC8tbB4xmK185vpPWQmSejM5
4akTWImc+P6qehxJaPAfBSoX46BjBWVYw3AmGLpE5dSIU4dLpHpXWF7lX6hKrIw2EqnYKnetFKXs
uxu+20BE4g76UfX5hJA3ws/O69/4wE2fP3PPXmBS1sPgAcITxpAUypSDifDKZovQ3vzg7YXm+2MX
CHJNYoqWPBPWq4TuIfcssuZPAIp75ppnQ9px04oH0MmTi7C2985RN4jT8Qcth2aMq/jg/CpK5BZI
10ze/ebV5KNTay/CAnudtDdzxJGYQJcrcv4JuKO+/C8sqVL5yEW+LsmX3arsofgB4zUxKBpX6n8w
9uJOJCDEmcRsq24xAoMDjfIemwVNlxGZvfnpr79FoswHLLqLGXs+jJKJPnQr8r+kFsxvPphP4Vga
f0lrr2IjgPxx2Yh7hZ3qlByvDJ+emnVFln13pARP4c1BBma7yKB1EWcnpeQZ65N1KK7Rdsn8S3wd
pH1/x47tYJZd3Yt7hCEHdk9yXMB2Vydrsw9DXX1yNMfh+qxrRf6VLho8hZt30wfkVcjexaBW3vSg
bSxiHjqiSXZwo1CZvrOVdCGZS69087bLYeCPi7gLMmKCPZEGnK17uLDeJatlZ7qW6F6K+fgEB4mb
8OrCIiDfFDECQm9dbJ9HepwMEAfjqSSbyWMspxKP6CJ3kB4paEkvZ8MHtBzNCFItlZ7gE6nKajct
crJMgWx1oSfuyYLSuGtz8Wj5Z4LP1GnBVOfF4rY4APZ4wNzjcu2z2FZs4Put2uAXDpvIvbgPRLpm
23/be200wTIrzrA6KtzFdCF2a4aWy6/kvR/z0HZBUJRDWvLEpp+iH8zo+UxOuPSOxRnVX0yVSAMQ
yHQkgpM3emAR9cliy3In+JdWu0Wc8xSjCxawCIWw0fHLVUNMI3JsF/Z/hwCNbblW3uGpCFMTgNaO
pb96He5jXbwKzWN8fWo/tK18MVfko0BZtnFFj3IFWDl4Y/BF2yceT4NRsp+Rmiao+7ZoXRj2NMAs
n5wAYVOJY/7Y+n3hX/5alHtC1yCmyDr1U9UmMPQZzLyaD5uPQyqpULqnmVzZaXsnGe0+uBAe88gM
WlXinmWgxHlB5GX28qk/xY5KklmftOXiUT1EaNMWRc6yeJ1to/1noNsZWDuYm3TEu17H2tyUl0ir
GgAelYkOm9GoZXklrn5CIbs7EHbVX8DiudJ85rPd7peXynczhqfs3xC1SmDMhJBP17mw8OPYGVEB
SP0/ay0o/hnni42lRhBNKORpFxkau8L6OpxyAIwMZ/Cc56glrncn/s6rxucZ64KSXeyfgaheQpI2
pYbdG927wX/c2+HSCBpbnP9W2mThIZ6VkDWzgHTqcdCkukQESWCdyKmM8FT/vsSxZgpGarkHY61A
DNqoGioDT5eoxy/25WKhWFff4P169B2MN6XgLOEz9tc3B24W424P81YWf69SFCbRHFKfjHpWLrfR
IZtvi/ivSnmtcYx7p0QaWLrMSDhNTi71/tsRRUmcN78AUuoQYb6D7oasvKJVxUrMglsFfPua9CUv
2jf7JS0Al9B/x0rIfHXJ+7A4iKTCpX7/e6xquYj2Iv11x5hI3ZHiyaG11bF1HLLGdg5NoYfKOgEg
H5mulw+c/fe+qgK9k2LopQExs9qBl2LaQBErQyz5yiGISBvHmdGgYUekZE+U3DCbEY37PB2bHiRe
KveV/iAvYM4/C9hVZaCFISmdjbjNx7YesAftLpC1YzdV6PMCNpwk3+W3mVxQ82O5LZosfJCWm99A
+RSzCozlEw1fT6NMbeI8F3uv+T8KO7/+NiJCiTDNgoGU7k9gCwMq0ajCMixTt07sDthDodq/XT6G
+P8OQbMP4/04UY3Pua39Kk2cJNjuJqhqx8sLWrxDzlzvtfJTlLDJkkqW6yGCYukSm7oPVbf9REUi
9rBxeIC/oJPFG4cHJ7jXAC18puZccgrLJyWzjmZlrEAX65F6+JC8ONjGs0tbTivbV1vu22Ak8O58
7sm5Pq0oPbluWIFCUzS4jrYYEz7C6Set44ccjOM7LtO0ggF9xopAs+hIuYgrJsGc83QSH7I8Hgfz
pBFFX668amPawV9hivLaYz/HwVqrGtYSf9iKCyzqRtK9m4bAYa1cAk5KZM1IT89UBiiNIq5ovwJM
q2g9NcqwWPukk7RzuS6oV7zq9OWlYuOW4ax9lY6c5M6C2NTTOpljBnQfDU0FCCNZmcn/HWwhQP1e
Es8jKj0Lc9Dm82GdATSYDr9vMctlrcpOTanoCirRGUzvupnBqAGWDjv4AhFzgFDSGHi2rFksF0y6
NUA+gVulaTD102u4EUc2rlx4TjU9IqL0keJbyST+eUn0QrRBhk062Iciuc8TFkFi7yW3Bt7zF98e
hDeDmYcFOmM/smbDs41zqOK26mUuEPakNJgDPPupflym1R8sdSgbKY3Vluij7VX4V6e2tNgbd7v1
2d3if7B1tkbCX23mgy+lmhRb5eKsf71npGr2vUOgg8g5T2nA8CqU8w/66IpTMjzFE5JnjuIk/9aO
x1igPy7BNUAU1Vgu2JE5hbWL7YdLvbMEEjh4CtF1R0R6F3FAHOTg32K9JnWgf3bjAfL/bJGIlzh3
ARmoYEZFOnlqMh7B6t8iZFg0XC++YMjBTgln3xtwrt7AXVSnDWJyPSr5FDOVCSXNNP1l7VfCjUhT
SdZE8Ppk7VY4+6Yaz+aiomSn9Hdt4rO7qdwUDZEN0Iic6GeuXmblFXNK8gSBj3R+RcROTxcAtccT
03P10tpUlSTwG7NBi9cLztN6TeFcr3nkU/WkXGCw33diIpo7M7luBgg/5oaRjiK10wUhZQHoqxVs
3qR9UVw3Dw9kaKBlpQKseAxJxHN84hFMq5ZmSx9MCOhpVzieeNfYLBgOio+j2fHBpojx2hA69Sf7
gzBJgZuVsKBLmdumkj4SyP+ItUY9Ek/LM4f6UfHiZ81oF0SzIBekFFC1fJ+zS8Q4g2aH3Ug1SDjG
nkRz/raGyC7a5Va7BK2i5WOFMgnW1T7z/WOpuaFD/viIQdhKEyQgz5Ejr+TE6ouL467x29HnVHqL
FY/Igyspj2o5Bt4y+iJPluoKrx/1aSSlAYgAxGqJOT+c0jv9iSzbwzgQFGcyVJZfZNtxgqovXVzT
mUraD44wFBjiI64EZnhxq27d4dgZNXg1OTwAXP+Lvf1ISn4v0eTbXbXAi7RtqfYZYDv14YgBELMU
ChAoceVZf6tKcDB/iHMpEksDzJtvtgRsxVy3NgrPsUjg/T4LQwa8LJcExbLWrdVNpyUJPoWqO8UA
83ZMD5EmB982L4FvZ4t1VESFj43XLsmvZAlZ8vObcYT5+cbkQ6z7tP7l3/Ae/139EV/Aq7fOrOAc
YI61SjlLg2UaD9U2JyDqEKlicdKsY86UAqsyoScVSSFJgHeBEHbg9lHRbjmh57BoAF2BM5eSC/iB
xGeXdrkGmY0+Taxe3NCw4BCGvFdK38RJmqRdo6UCR40zd7U4zpDADiIpff2u9Ue5yq6Y4BHvvzEt
sKdEeqAfT4L6b3mPgg8MTfWIXhSKv8mprajySMUX8mq6hESXdMygDR0UPGNZJZzUp9QEMVmf90UW
1/n6uGYtZsGQoSL8k8M0krrML9DesUhDrVuBoa6LKI7mREnqKyMcMd6L45vOJHQLQzyd2U9/tKP4
HH8NmXf+KZVql0EbYO+a4AX0zYgUy57wj2wXLAzMCzycN5CHFCZniWHrXC+puakXhvnQIE1Vbyqn
Y/l16EakoWlXGdP47N0U+32vBhbL3MOUEdld3iep1W4c/jZ9mQepsXK59nNCYV8k46RkDQ8w1dfK
hYu1XzRH6oOg6Q1+LBw822ElSCKSEDQwqY+zXbbt2zsXZPryWG1SrhB+VtNZzfdu3hhxEwEMQ9ij
vFeRMOxiDPd6TPAxKu46HgF6sz5XAWpE8jZXVamsYq5K6UugdCbka6Z7dPdD9PAQxU78RypbKtl5
c5NlGmvUMJXcPC5DDrUT2SmAWNukXvIMwFbDV5onweu6hFVmRFRMsvdUpQK5MTH1vrqDA8NiWdBl
eeCaE0fo6RK1xlroo6QgINm/gc9gpMmqlwM/QvuN+UxR08GmgNESjiaBw+Z7PFxBi9QFr8KUWcII
SJoR0N5Xcedwxx6E5WeX4FP6Kxc5OCJlWp8UorCElQBmfdyubFH0+5ojP2YCsqGb9WBmmOMfuWh5
a38dEw3yHH3QOsi+KHhp1aTjSRXkw+i7UB0M5K324O8mssLsvcGQ3zmWJCg2yQEBd3wGo4dTaRfy
TrMK1kipOgoC7DOr3ct9Z0/KUAsNpI0iz5pfN8xO8HPYpmll4DUvCBKKoHYOLCz2AOUI7VyuhXJM
u/XUlKYV+Pk08wCTjKJ5FuPSUqOT2Ho2pc+aidTy1eR4xBni3igtT/tllY9Tq9nnBmFwSKBE4laL
MR72ZIIZEBpjUPduABDg1aLC3ASmjY6Y7zayyLS+5Fls96PzFMG2te+jpRtZjAdh1NM2tzR2lGJJ
R26NIg11YkJVH2ETQEb+7a0eByVd7S7d6rxWL1JiOoNmhWesFgOt5KQHl/HDOCQpNUyXlrEyXI1Q
dSobH36bI6kn8sfYWdGQ1INJgjaGzNETseQDBHhmpd7bQlU95Ph6qT1TEdOJfXmvTKr1ZVBMB8fE
TgB9zYXBh3bHwwKWjHCDsaAf5NL0Ex4ljZiVXfgDHX+ruc9uJdupN/FVX4Tnf+2fyrCH96zgC9KS
1Gls/Iyo/LvTG9TZdviXizjEfst//35kWrFt6Itqp8lVeYeownPyqxhuBO12xWWi5IGMEIMbW7+s
eIG0yYWXJrXNOy59j2UgOSfKncXglUgJ/Ij3QYYWz8ye61GzaPdS3n7TkYnp8GyDc0Im8Mzko5cX
9x57noYuvwcKMQnTdH0f/rQvQH5fvUzQnXgKVTfIeEmrl8uO6QtGaRP2bcrSq2s7JY0lcygJdmX0
WoVOC5DdxJ7zDTn9fHhfEjBimeBInZnwjvwyeza8NLdv6xwWj7B3hxqv6TyANlAFrGGURWT3GnbR
u93nqVY41k5e7cx+yIPFM7holH8QiiZ8icDZs8BdRmJpRIqro7fMIrAAgEveRe41NrtPrBLavtIa
M7SeRNZuroyLnsetFyWSxNnsBYSBfQ+8IhuZrDfsVKPrFzN1yXGJBuHg2pwvyWeNq33rCtc0TAKw
9ZLlCgiuWvXhHGf//1uMMUNTw/8ts/sYPLQJOClHytZi9lflqTzbLgcinwlQDq8T6w3KeWoMh6W8
d+PyDvL1l5WdyG5tntZiZ1eUt0mJA7FPnkpqmnvDTtbskW9fhj93yEkyLz7Bj451V+0w3mc8a/8h
FmghQUvHoGrjoyIFDRw7c6bS+uQ4fwTdbm18psuegyw54UbO3+DapZLBxlzgrLVEEeNRwObEL6K8
HB5CX3yPbfnxap39Gj+JG8izZLgTaXycuvEyw6hjY4S4H3S072WxDemhXiFZvvcaWp/K09Ay/ccx
mst9/xqwe2sBfrIKuoIYKXHjXAVzq1HGiyb3fTos2pPlXdTxR0pZM0iEzxS3PCKpzg10PJiNQQTn
HwP39DL9K/nSjMAwECdPh/G7t2EyHGS3ppTpvKzNoG07azqy/3rNGjbp6E2vYd7f1o/fd9HxhLW4
kykElW+jrJjGZm2rzUXF1bTULy6ZifMVvMuNgYXP5wb7O8UeLdJO7S2BMUaTcK+ni6I+dOpz34aL
eadJc7dR3SeN6Ayr4n7HECviSRMl9fYdx6tZgBqg5TnnI/PtYVmHZ/RmUTw/F8+1jvNqOxJTusPa
b/h3pXGXsrPocLVXpgDuk+QlSaG0aRuq1XpfQlWEcWiDZlIWy1MY7h9yVNRlRO/pqwyjVGJJgZdL
k/F0UctjpyW2gRI9DYsIVAESE3N7Kr3ocZwFtvrYMfko6xF1CytS4a1dyKbTKhn6446CJUZasUSI
hiCxx8kLLlCQmO43fUxpkSJh9p+IDPXFbWoJFmBNI8tIb/Gb+FX5X0NXjrS4IZgrACkuf+PQhaXA
rY7gFYqQQzWZxynmAKWeP83uW56HOzvfahxR+2+rTWviR05nzsHxFsbd4L1jNe0lf6x+poSz+XDK
PtSTn7CEYqhaY5a6mA15vy203A95FuDfQQb+IC03jPLtJI7OcRugyzjynkszk+3LJ3EQltl0ed5A
fU5JyttpzirV/YPzNH+b/sgg9ND1Rs7/dmPKXvrX+wRuqjD71PU1NFXN61QWxZ+WO6A4a8NTl8vF
myc+LYhHTA0v9IOeB7GJ4I4eGwWeCVYVMVp5zGOMN2qL5PQ8cnqT19Rkv9TQhn3BDneV9sd2yfGx
ncWJ3hdvvCFEwvIYrpwYGbCkziKaJZxhHPWjVxG0/XjB5btV1FYytT84HDOqTLbx9qTDk1rWq0fX
j5RVrkrnKCSnMHz1BqIYbVvIlS/SCBgkZczqHSJ0Kp/HRpYExpLx89zitpHIamc0NkXhH6Rn7kNy
kctwX12OQ3EkEqkSsb9xYgYMeWKpv/5AFP7Loxz6gyQ7EjpddlIvzskuy//Za9GToZ7c1Ed0Dyhw
CkE2wAYhWXERbwO+GCif9BmaSJlIkbOndzk1ZI4dQwbda3ubhQDtAlZLGJoMO8UMpbJpmf6bXQ58
/Y91WfblsRDmSQATymAPprl6WVkfsCVsnNgPUlxvYlWOliet8WRCzl0mwuouA70SyYUudub9910p
7G948qeNu5hshFOnUy4q4hdOlw73SjYKhkSb3C9it0CSbYfJlbV/OWsD6mPdjSk8JdxUJqm0T4nf
R6DfhwJ697Il70GyRam5tJ/aqIA7FHZ7pmf4MRBYLEwaF/RBDSGZ3bZflLTWEQpRN6tdACcFVUFQ
SEhEvlYySKc04L06F66YPGbN79v9BbVY4z1cJ4Q2LsNwzT1GxJd2wLlcPd6NELK7MfJanPXKx5jT
6HmfMydaSOBJ6PlN/bFeORq40K8AgY1SNyNpugg0wgvnjc7dkW4cdXx72PtIK1tNFwwc5wbxSa4L
SGiiwjCXMe1bcLXtSC7DWR8qK3dJ/jgGCLiMylW4O5sZ9rNR7nT3//z4uzgYFOZptyidic9xBYON
s2K+YHClh+QZV/8/bIqL9NImKy1gJWZYXboYc1IjwSNTcYyGV7sLVtn+lMUwzGt9gvHiAXaIEkhc
N64WByJ8ujbzq2rj/00COWyi5rIfQR/wePjtEfbNB8kE9+pfUHQkVdqIpfvdjJjtf4uifgauHOxk
BgnSEQk71KObctmIos6/AzdPNoys2Yf8nBHT/FsMqQqSUB0chzelBwxHpmCm3azzeAiP7t7VS+dw
6IKR4YCsd+cyelf46zgRNAPWOeq1hWcWa0ej6UBWDbPh5rQW8oX1KW/z+ybJFA+Ko8Mzb7kjmslq
tk2P2j2CKeVqXqKBaPOCq4ugOtijZKamH4ow0TY8l90g3GdYKG4YYtXYr0JB6kkZQ+vl6q/wEkZq
1osSaN7a6k66ZICylr/g2hu7YWy7IR2IobVMrvf4c/rQPXE3Pr86kxeLdvIDjhZ54RYmzOc0v4DX
4/8nJcRmQT3CS71ve1lotAgpmerbRm/f8GsEErNKU5TctlbjL8fs51qHqqhW40C9RKTfy4YUPWJR
7SAAvH1TytI2fiL05wojF9WEXZaHKPi5UryZLysyhXn0dYzJJMt3Loyq4IacZlvrGDzjBu0s9pl4
UtPoGi3GWCON3l7MSvrndDA43bk0WF+1PctEh4gYqHnw4ru/LruogNXVOqHSk4iHOfjjg5OCaIfY
P9pyxs74pOQ1W0WrocPaUYG/2LtwtcOZPXSFxA8kBBd7IFaqFopy47BM3gLqHoHviJP4jQeRDuyx
gn6g2e4sbPmUC63nDnU15BJU9teJoc1xIycROBeRlYIzmoAWA+NWfYkCOYmdWZB3cH/9sBbqY800
wEfww7k06zlyB/g5cMckJwxJP43vyb1dC+z4VP2SQilBJvv1Or1S7MJe0IE++wfM8X1A1MpVwfn2
0Cof8QXQ0FM26XFtzdJg0u3jQuIo8N4J/uv3Rd8KUIrz84JRu0Us8e0H0BaZSlnKkU/elf5meblO
1G1v8k4XHd9BHqfWTBM3ENVZeuETW3uPu12vSZUsbhvP55ZXWsrf/W7sK+W6gAu38x0wxNSvnu9h
S9U4667IZT58+ZAoUmsvrW/BrDyYgLG2CdLEC6VNEFUXA4z/Hteno2MQa7cyRsNf+tUpMSzK1e4R
lj4nrsMKUuVU2+jzBNziCikvUl8q5bIDK3V8wFhnGmaDNGJ7/YdlaI/zcrTfZxUPnNEzh/zzxfHX
gitL3OU5D8gw/H4X/qnWmPTYRDvJV+3vRdi6DXK+B+3VR8VPlM1GmJ9hdYEYD/l0OXYe8gijtxxi
cqpiGco6jKoB/fgFoTNy9WeV0q3b8mMJCkia3VkcJXzpTDy9naLShGq8caWCfN3kDCK8dJQ9L28M
0FcODK5oF7YlHnKwJTyma5MLPqv/83LwCHjI/8znPnzjtIqGU9urcCSI9gaPDv24i35QdT5yVMIm
iG9YN37rscuq2sS/VrTmnfbX43EIiWPO1AYdAsLW6RSt3X2tX3PvlMmluS2nukfamlmQHaZBy+Mp
wSFGDA/WpsuBvb5W1WSGvsb7/a4SFnhCRR8374OeWqzjHF9GqWRfAHE80zQzRa5JgX5ZAGDM+fL0
K/Ej/SPJ2ZLBempB/OfHHcbz/IOAQ5BSAsH91kxAB4zrFcfxPgOQm2o3e+P7avlhTq8dwW/7L4er
GLx3jaNyMo4y3k0VUesKD37Jkj924RnzzEAfJQr6cxBxKHHOyARybHdR6y+B9y4oKoS5ISchVO0j
PKIpQ9T1HS6vv031sAiJ9w2QNSZAXCeNaGybGxbzyJ87chzZaWPjb3yntdWLJ0rvZSd1ew3uDoa0
Lr7VTaefpJfhbds6Ckp85W2uHzSRBi5p9WM7H9DlhGcq+HH+5aP40NB8tBdHmVkoNZ3xnqTh1Fom
vtkwN1m6RkLfDevomJCDSc9gJo9XbvlLsU5IipvVc/h54SmqlHGwvPK85WaFCdHIXHVzQMGISuHw
HTJdmOA1it2xElEN7jAiaLfqYX8xo9DjDgx2tLEE0EawH8ATvE2L4oleKa4mWdA0z7fBOF0L+mR/
sB6tmGNbPedVvO2kMyGgR/TRqvepKdRQm79BYq6qm1OuUcDOE280ozzuCtBKKrquG3Qis3O8SqI6
rAIg+DOb6sRkmC0Hav2zE4a6tjWxVwE/W04V0s57bpVr3QMnS86ZuioiD3kjl5PdBNR3vPSoztp8
HxaI6hL+O3dlBV/ErBV7tHlp2oVtRS0jtQtIvhlUCIpKFjVKsNiR9fJquc3eR1eAVLKYcq3tDOuF
hooUcH8gfSjQs+x72IWokEL5A5hOeRrlBeYIRw+DQJNwxzcJKq802OW0DTCOpAv6WqHRV3dC3h9g
n7N5Q7Ly6r+p+xkWxeAU7OEV1h/H//UQItooVFQTvp8GwioPXcJKKJDpvSlH45/1pq7NYr4P+47b
2Z+QcsjRzAsa2LUZOjLUjrcTFetNrTQqV8f4rMUZhyefPw6fROEzB35IrXV9LhxEm+/yRuGdFPOJ
ixcDUZK2/qEgVeqB8tIQU8QDWa+Ivwzt+4OU9Ai6fXjWkBlPU+WS52mLf0m456XeJ9Cg2Xn7wnCW
ahckb4FHQ7yKzjcLjuSsOt5P2kFTiwvER2mcl8u3OqTxjhKfae7+RKWbdltZsMLgUiO+4/Acs5f3
/T0r7ot+cBZF3j3Tt3j/UTAkXoWYlwpllWltHBtijthhD0KCd3SD0CtFo17GoLTg4kvuMhVrLQYG
KqUwxsD0Aup5ImICGzsA1e/UA+phEXrSknqQ500NFJd7wO+yVnBmoAwMZNFhHVkeGH73jFYYaROi
DXcvJblgdLMk3oxLskSs2oCmPGGuTYX3tczjQNwej3GZhU2fgd73sMIqedrrwG97QYvPFfV5U/BJ
r2YAa2jL8VYVzy4HAU40BYeixq73a+KrIquQEyUXjkjPwmSdR7ZVOpgB6T+m0o3iD+0QC3xvgVhe
3rTSpoOhsWFFoW9NIYx70chD4hKIMBtF9MwQv0ptikJJo/eaTJoEXmYpj6MyRdM0sdYbgmN2qChx
iYahomKT2MdGOsVsd7q7BWU0InO/TTE0thitLDWoTqjXVPS4uX7MwN9x/MUGHD1gJvG7SUinCpTl
2pwoAYNadlOm/481DrENp8ZW+dp9JFFF9xfgcUrjZ+5Ys/btdJb7CXUPAQ4PVv2rjcaoIa9YPpPO
8a6ShE5KwPY2rgHm0dTOrG3BQeWIBQ1pACU8BOAFIlank4SQ4FJgEQ4R7PTwzgd/joGN8GmGfPQO
mgH5DGqTESLM/R8AJ7cV6y76TPswHhOFEax2nD3w8vTO1/bTyy3xx2rPzQ7OvEq5lphY4irGSZGW
Srgc6J6/U4KzVbq6uTP956FayXeuyDUOxj80IpkClv1pwEBQIYPQBtgSLX2oSp53yuUkZjGhwJqg
yrR44Y+6J03Cl8F5wOGLj4NqwvtcVHZzykuEtZAZIrv5367LYBGF5nNRBJc8Pm4pIE1/ZGsVAqCp
so/vdp5Ymhk8kE3wLZO3wOcvwfiKcZtYIF6Ug92XvtHQi17/S3BlGp1thmi7ui8+GhBOBkF1jiDS
CYoVj3mtZm1vXFq7TUTIVWfSAr/KwCGcvK2spFmJvGizePDWGapSqAaeHhunwqVSaBysa6avRGHa
m+IqKZvRdVbF59Zl6yVD7XBNW6e8adhXMO2X/jezFlBWEP3t11EDr6XpNTfkoO1V5CKMcUdElyQ2
frgvzX/Ln6luXhfPlPKwh7BqF8nRodZRcX9Vq/wRZ5YkgUWfI/+EIJQ8rExo+lHVPcdKfw6Fcwqu
obQotaV68ZNCqN4eJw3XMEAn1ydMvijQTD5xilJva8wmcwaZGdGnBRBTYwp1LgYK2J1moUYyOYkp
krvmAs3ixeUsRvs3e2vkXtchOUf39u3V8dBFpSnSnNiiXHAlBBP3UYDrIGZwwT+DR11WSMbKuLpC
zFZotaBY6mTlDaAV2NfQGgu9gNwE/+D/TX9gvikOJWjnd/CMc6UAz9lvnVitcjehW8H6bzJP7kx+
5dlNtMYYV1tjB3SoJxYAXWirJJ+An5LHQ9Jt4hSb8xsKrbXcLF8KBGTzL109Kr2ftjSSS/jPzau5
ztUTQWecZWgAWVaassm6u9oZYO9CguOGU6v+KAdfvdg9HKEQPH2IEJn6Viu3mgMi517R1uBEtnRE
RNgr3FSOVlBaFCmH4ickn4NSta87qOjTjmww3AxqbGDdRKGEIO0EFyNq3AZBdpydRVjK+am+lB6h
R97rf44EVTaT0LnFQIIHEbmRvs9glef3v3+lE3kPxDCORdhihgA1S++868QBJRqPj/fxHnZRZqoY
Q1iNIMdsSIKT4fGYslM6rBintXAryLxp8MweOIq/4gGaiGOKWVO41qTwDjZMK8fHLVmtBlbfmxxu
1PSkTGB4zAWhCeB+tGcmgHRu0LHlJQn7bUiC1d1/98JrvGg8lymHOaSwT1B+Cd4KB+utYDxLd7YU
7gluBRG8oQrzvJn34e6ZMFhTDsriC2IDlemHXdcA5Cv8HiIyh3OTbqB768TgxUvXQY6JSuSBesx2
Lu+F6qQQcXsGdYvYtkK8SKg3rRXZ+DZ2ANBO/b2k+BkttyJmypRHja6KBeUNNpoFEjRu5Tu9Uqfz
+3KoUvqsaP9NXhwzO3ChBbc0DtE9GjCcTIiVfNoMd9od1dBaMKy+BKtvS0nsx8DX3HNun7HIye0f
x87X/Shw3LR8ZKles02osFHeUoELMNIFo9REfFiERDTsS+5mYIDy5Xqvo6xObTuAnOZZR/nIHPj8
Pwodm7QuSFP0LgLfKdVEVAwJ36tQM9Vwl7Ggfus3or8HvMg/Eku5/GTfh/wUuyMmCD4k0RcMH1/a
5JzX+gggSOuobS1JOTuzDxB1ZoTa67zYGjuZIX4rhi+hN41D/zcOhmZNbyFHziNZyrwMCVdTelsN
xoLPUfdt54lMyER/n16wpy0Io/K3MTsu2O74hzZ3R5NaD86JIGr5ee5AeiE5Y6vaILciEFCFab7r
7XG7IaV/Cei2R1/WL+9BoWk3lCw2ljgHTWi5SSZSTEWICP83/mRx45pyJ4hg5az2KZ7Y7ory6l1N
Sm8k/I8pigFDKVtC3hx8B4dlLO9/yKtVssXJqIk9qEYOhWUVWbIqKDLzHDz3YPwsckl7/TkpknRh
/jA7vl1ZppEVSLLyjhNJkFGbr1UblKylOzFLZz7CioEXk8p7vV0xfGgoV0PNU9eeblY7JjcVu1fU
Zl+hJqsgh0wy1JzF+Iisxm1bzqsYyxvWrepgP2y/ppN5Ux7arR4btFzkeV1eVTY8aE5pKTA+SmUo
ux0gQtzCqwyomjPxgyYduOp42MfiglDpYyZIaTlF4I2BQ44ioVjyxRnwK2NIkDhmLXmwenrXzvvR
GbEAHC5VbGW2IZFN6T8cUyugohKkX0DQUPFOe3pCE36Bd66Qg+xToczicDqUOy2hvCoTC1ljYZF1
Vtnqmt/PveQtUSFfCSCec041ZNmHMnpZvAlefji7D1DmlkUfVzhwOBSi0UKPUUhjLChi4aveIunC
gmAnVMT8nx82Zy1LR16JKpIUtLJC5KNy0CBffKjENF3fHd6nKKGNS6fcKSZ6xx+X6ZZMtXe9fE5i
PdftYD+sVHiheyVHrJsyphXVTyKTcLWBGTuhc04J7KSjEkDd0ykuAgXZySk22jUq1fKC284r5sS3
X46yRRnv+8+yWTOL+25tDivPDvmWo+ypCdHmxXczdx5vHkm6NOVV3/CjzWYU1t4bk8LK8Fpu2Uam
P4rP/SxKKjsRRNuoiHFyWyq46hLLW6w0b+m1eFfU/dZ/1Huldm8wTEf+xrzf+s2mUk5IjezUFcsL
x+qYtnTrb6A8HX1t5EIA8ctVxnlEeQDtDX10BCS2uinJBArzxlovr1mimDg4LHHLpPZsB7cQALLN
ZQB9vTYxptTJtZ6CZwJQUbwYYa/XvOgorvu8PiM2lLFq+2vl3e+ImD7JwiKfa2StT0TtDkN+HnXl
iYBV/ehnYTXTjlLWTDbZ0BmkNUK1QnqT5lq+Tk74MOObT8ZwfmELz7d47F7pyyV4iKGPnTsh3oIh
6HUqCVIHVSJHUV9h7rNyZohhYf8uBLyFCR6CPGWdWEYtEmkmgZUCLvTRXbAl9TIx9KjHuW/I97ZE
6g2C70Z1rIUXAix5weDch6qHm+tubgZEccofBmEi05SrhHWz53PF4l02wfFhBYLbbdDMllVxploP
Xd5D7iK6Quy+5Oq/+/y3tdUzk9ONYbLdCBpgfF0BPkljAJ4xhY7yPUrDXIamYff4dL950YPSai1Z
eE1QN8DWcK+XGxcpOstqvwTa47gJQb9Kk0VgaK4SCqlrdFZTrzJUBP7gXtI9pbGIj50pogEiRE29
7mWyUIbBZCK5icklATotlokymT7Bg7qKZ7QkGaWAx/b6NPqQSnZe/Np2eCsv8oGOJaA99uGVIKkn
hlGoYE0bXO2rrlXWLPu5suzPgnwoiqvaur+xaxsp6zLm5oVerkeaN6SO4cvZ36ZrFUgdjb2mqr0a
CMsHeYQbJnxCPS7AnysDjqsO2MHN/onJTW0eTm+p5UISatXCGfrF2cFbtaOfOTqxRYj1wpCJqoc6
LLC9Zb8PYtTCZRUrouYkTe7u3LhM9/pKnop0q3850MR03NCv73TrE94/mdG8gq9WIUfWBVUSV9mF
Ux8OjyF+sOZlv2BijS3FQQ3ezJdUzZL+5NftO0VqO1sluQTD3M1OZEGSPo8gpYiKx3Vb3fm7IrCw
xnOlgPW9IAQWPViRMStjbVc3V4mHDaFmLsCOAAzSPnpzzpEsyQO2ElfYF+Zt4DQlIZutqbj5D5bx
rPSTxZ9fXPEgvefs3tv0Xl5HMaaM9YVYd2K64xrSK/9sL8kTfyWb6RDuq8ZjwiJsU9V8hcZwCYwb
Gth8op9PKpHzd8oLaAMto/p5ZyTIhraJHHJKU9bIO/dmHuhDQwFKXokOTspHxrXPC0hU0iF+lfuO
nC2zeTFnqcNiYty7hA7VlKoq55cWLU0ZjB+cy7W0heqOz7iLv0YMljrkFw5+abGidmN4BubKnNSG
7sedfttNKfhniEVhrlaNeYCIc/M9mgTpZh5yxokV6Sd5jDsogmkkVG7psTiDKpZ5/lhEmWSLoiy/
UkLI70rfSaVFZA8D/HtM0m55UVO/QlhYklqptX2xus/jnDtDAZkEkSBJIAOfyz8JEMVBxLa47ATe
xQtNbF+b13G6C380haZA3ChVn7HFWm857ImmR71ERv4I+yqScbB9mDmK+D8MFZqb2U2xFQh+qx46
16/plxmYGiz0zZumO0WV5KHH+UO5C/LiGyEdLQVyY63IfXdxOpASb56dVLD79n4KhOd+Ce6k7vhe
WmONsYYjo7+AS6ly3NX/r5XWCovTOn+ajg+dFVAwGXIraOHUlUVnu12WGCgxtNArE8AH7sUzVRR+
s6Gt7g41MYIuam7sWeGhKN+5NZj3nJPPVexA0PVqLFw2EXkXUZS3zPMugOEyGMQK9Fu9JNJCIb8e
3HPGsFreKg6738DWGgmv4dBtZxz6TJu3g6/2S5pWleacyPS9Hy7b2Mt4qqPD2jvAYuIHIb5GRg1z
UjLLz3RDQMYDsAVRd4+BgWazaJU4vNEH4pfMPvaEC3GFejuuLfTUiRFFihCTTa0cs3qGWEa59lCv
lcn3WJaa+qW1y6e38lf6qp78kTkl1inrdrnBXu7qWV+Anyumit+23+qJ0CopVNuyPKUq+B71FIap
4wYfwlDFgio0UGA96+bPUTwRA4EDMvm5UaytiZgxVAoJnqtsTwIhM1psEI0Qa7I01h71CvVkImZU
j3iCRBw/t4vOIOEXiVfiwMMXNUcr9zM0diJENJhoK+ZOLyO9LJc+ztlzfl4SFNmwtVnmQmiKpltl
HHHh3qocGchfIntTGlL/Ls5dLzobalUOa8fI9On8LG2gLp8ZCrAXsAL2njtmGh7NNYj+omUJahai
Dw9lxBNhLAnPdknqjacnK1a2i8i+JLe670nAqG1Lp8Flc3OTcmhQeki+t2BBRKw+PTBa/wIDgejU
rZK+mc4RU26CHBSPw4ZZTUtwYzA69hpR/j6JieYzewGa5k1GgNMPZDdDIJ/p4fBghwD6xP9rVe8E
hd/s3jsJOqxDXkD27i0OOJsE6QtfhWKRkP8YoFropbrKm885ctJPhh+tXQ63InYfFNGbRGcj2mwv
gfoNxYdsL0YWJx0IlQTelCXlrbT1UN2Y0r5KjCAEh9uF1FyZvYMcFpprsDBXJecJmB/XFBk+2+Ie
2BYiHX5/8+PfYS29hnukssYRq1XsN7OGBsJ7tRtnY8ZKd9SgX3+vNKDk5rPd5RwSidxqk0eAtHhH
XtNIKXhBRF0AeUGY/HKxASBcreT/sprGPD21vxUQ8yX4tttHPWwr0gDiX4PqkMro8zW+zEXCVmrs
J3OcsRxdaAQjjbROTxbuCaY5WUCJ2BOSI5nocZZOhV1o7uoJOHpo0uMA9pkTMRDslSf4OTqPvrID
ARQ7ACSQgbbuDVJxp6JH4J8YbgH70AGTZCg1CSsC+jE/8KSiRz8erQS7kzsjcTZSZ58UVa1PvJLU
UFwfkUsXgswCsUnyl2OPn0zCh9CRKuo9LJiJLKaCpX2Qm32fSAT8MphNe2acvEfqX5GznTcTZfHs
aG2cp6mpi+zV6LU1Dnua4fEiMePCv3dTsWJNMyYajoOviP7bPUUl8OGecs92FcoMKO6RFJWadI2R
9jZin7YH22xN7UUETKgibSehbpSQPlRo4yYkmTGghBqQCFhd33LkYGcBIDdCwuoB/q7o5EpXJW7U
cLO9Uh827VDGSKLEnNIXrBqjBFkRXYWLbKRZCQsAV+g/O7CFSuHxZSFza7ljVB32k+zG8K5UWno4
mA20Mcl4kF831hqs7E47IMD/QW9ltucbiWazHffOa51k9dNtfsZwZcWomIqvb57RyDHuw2hcJ6s3
JSu+Axl2KCfgD7WkTTvDq7E/2xgN6i3dBIlAFCMeV5nX5chh2FHdNdXKxrRCWkVH+FHn71D2oX8W
Hv+xVllMCuCDOEmtpLU3WgZQFS7+PcSCLaHJjTclXjw6vDxcBWtDr/Mgeyqh1W/0fQDoJV0uRWWg
1NPpPW4L4oykRIeY00b2SmFVE6q/wi3sdSFqvUqNbKncL9CJ7QA+v0k/IpDBi3aMgCAoQ5L/rjlX
6HlY0lVosQPVsWfkIHr8VpmFFzfbg/M2e6vKqxIxnW1CnJtYAtQjMc90ZHPyxaknqiHYJpQ88XAA
xGaRtqQibQDFkvtgCFMHH5w5DjYeNbDS1ongjExo+P705CHX2/7ZN57qmU2Qyph1D3qVDk6eW3Yr
fZtRrH+mqSBU8lxjgjLphUkeziqt3iJ5LMlT0MLMSItWklZIWOSTEKAy8TQnLebAo4H4Kg+vn43Y
glBk3fo+6BmIvNoZrZV6aKuLylRVlLYlSbLIr2HFZ5xqHHUxK6FbI3L7+fPSvdrcWY74IY8MSD+p
F/PKuCHc5XuS86xVorWqX3OHKbHwnkzwHXyHQ7uAQmpTaV7rPVNqDwGY35a0NRy7ljvAv/niUV4a
u2vaaum4XTmBmFQP13kG9b4ae+BhvDnyPJiDW5/s17WNHfF7qEkfoUZpwSjH3RxRjvESomqEkviL
SV1RNtYXnEUpX7pXXjPXP06GKKuqM/CCrLY5txhm3P493sUpihi3VLhTnjkCu8tJi1KQh7xSzZvk
vwf+wcCagKVnt4PllJmcuSyaZtHboIN+WCT7U/tlLLCJxxiORVBUKh0mU6/mN40g8D6nKGB4Nj2t
X2KLDegh39PRA20bp77P2iqofFAdxLyWnlKs6FShtv8Tg9fA13s2kGvddFm4UoXf0Kk0uY9bnjR8
A3wfyUCd0ibFvTQNzZb8tW/PmYCLPc3ceH/WvsCne0vRFQwQmHc+mIMuJECFqBacQmw/OstKEdjb
kTTTCtOanKJUaQKjiNWWSFyMKMqQcA2tGuvEz8YX5xbn/CZm6BghRJh5cRrDShqo6lUUsap6xD15
R3PzJbVMFAjcLYe5yRFUweQ3zQji25N8CX2xcRiZUwaNoXo94eSOlGTQ48Bz3vf7XKJwUQKcmXPD
5bWwYakogd/v43csZ9byt0geaZsRfasQ0vvNnHT8XCqXCqSds8/05H3+btMbIEp+rppuIHJEGFTD
itxUvNP1fJmb7caM0rzpqrreyGU2tWcLnJOeuBB7RLvF0uAZ+n/mpcN+j458Kcw9lIlz6CRF8D2r
f7817QN8bXseYz608EnRQJfySNdGyjF/di3uU3FZdOE+MfYNBkmLvERiqzggNe/alE2IFjHD7o5U
aClBWq/V4NSblviw8RkqrCrseoPgc/f6gDFqGLozhjrI1uBy13A1rTMubd4sbYf6iJZ7K08skQvf
Tds4WbqEd1x0M5FKG7qZp2vNmsUa5M35c6Q7yBINpFHygUqaghSVASAovrTx0oVvStXZ0Jb0jqp3
E3MEAzJ5UsjzTK4z0Vz+F3VzJnQvNIYrGB/B/OvrqCXDf/dABgk29N3vbKo3YdQzPXzVQFbYrHNQ
bTlimvEDNd3fuhkRJxXIyxW9xZrXznrG9kDzmxEUkTe2W8Wjq3rrBtTBhfcRU1BM+HmofhQc8Q1e
ZxB/WWWK1KfEB945yg3gzicgBU1f3agSWInwTwOmrv3pGrblFfbNbuxqjeQqN3WQKBh8oID2/TH6
whulM+6J607dp6De9rUK+zf2DDAd0Pbym/Nv7Omc1lGNN0DPNCvkvaY5++tciDMlMGtF1uCjZvhE
fws4B/QC5+mJ4mN8Ko2KSZhxrcj3bC58+ogmxPuJe0krDwZPwlnY/lFgSXHDigXSlvDr3SKOj+Su
PEJvEM6CxVfvrM5aTDbEmMfZpWHZXd3Eq3ImoOqSdzldS991ylgiCEvRjjMnD5Tko94o1zRel3Rq
+vZMxF8cECKT+qIPAUzwxMgWQOkK3x3z0cR/6dXaNM43VdW6eqzRtgyDdvhOaNe9gmnxuOC2tQIO
vbafyeXA8iySaih4t6zkb0jA7nZLsLpnHm+onU1zDPuqgQW7jL09SHeHd7Qj6NwPcmseAQ/l46eb
L6nUsLUsmBSI2hbQQpXnvWzHQQWvSPDCAr4SBKozkgZFUJNalZcJWj2qRc3xJ2/gps2Zn8xX0M1X
PYC/jBukOvboGImCuyEnRCRc5inkSJAHiAWz2fwfL1Vp2TWgl9qpel/xs4vhW1pyAvrES0p8s64z
GKtmymNaVl+ac1GX1zwf/0ejYdJdyPXaP9mQHRiXm8KipIUcSNzNC995hG49AYxLMzsJ9ADXT1XX
PQG1YSWaHKF/sABUnNak03wBAs+Bd6wO2l3T8BTSWk9rAGn5raFHfSjHIGew8MJTRgf4ATrMrw6c
m6UzDeMykmFqhQo308JZOfCsHxdLmE8w8IWMuyiH7hBYs5gpqBZN5Zt+8A2Rly+UJD1PQ8hTk54b
ZoxGApaKoGDHnf7HuY8zBFhnBt+uce0jGqEOX4GkcHTTKiNqXUGOlNTDH/cZ80FicTv81fA0PuFk
SRvMwP0rH4psumNOU7ysyzTqUojyM2jQHSBj9CT+mMQZg9Co7TuKbR//KjlCLa3SpJWYq8QbfJDQ
e9mkA+x6sj9tnpu8zz8z/CbYIUUjVosB3bzQq8BcJwGTgeG97Ev4p2DTGcfRIALrnA1nUOvU8Vdb
lTs4H8l9s5XfM8U2al7QKrsWiTEapBa9rWzNGfDY9LA1vjvI73L54Oc18ye3Jb3KU88M6b+Zdydu
4zxka4vdLBkNJZ93IY9tyhurSDV9NL16dZCuwB1ZzH4YpbJYbvRyvSj5PYPD4KrZq2qVzz22cH8x
5j5c12ZyYHHP8ZPNRZYEOFNLe49YR9tb9wHOe//FwvWnRa+/l5JAihOHSNeK44+whAWQUxuj/F7Y
9qGdXMkS8Qiu1/d2K4rNZzwhNLMw0PoliM6Wcjc4WqWkISa68aP9vHI8EagcQ2m2uXf1ShRbc7OR
g+Ut5r6AMRYtDxPG3g5BN3+63I9IdwC+OyAbB2FyNWrpl2Csn7UkV7AQXJXJ9cjrBGciWz8zxl5e
7nEWXBcc5hbu2yvHNAjEvAz+nyJ19QTr4Q8hoQXgxBYlYUZMR6JxPFvcaMeZkdJ9U5au0mPq9hV9
fV8nsDOZf+V3y47cF1Fjvw8QKogUnhTdA3llPFe0Wxv18FHuYa5FeQzdos0LzTZNwhxahZfsFnr2
IJ1el+0pFVMH+aU/7t81Vli9k3Bl24nNpAYilRFm4HeUDWnofbiIaDsoLyzh1m1/ZNkoOy9Xjnex
N4jY2B9s+cz6MQQN0sUL6oqm2Wk1muoF76DBShBU5BHvMM/biH3Nec836Al+YIDH6DQ064F6+luI
QB1IDak2U+rnEDiSOWDs+MCVxL+5Oq19/31LQPKtmYqa5KA4XMbOaSyHJSBV2bwUzQmPG+vDeW+e
SR/sVsZ3RitkcgjX/azvu5abmAbWnQGPLFwSdh6bjAtlO6qtQF50/Cpb3qWbAkTAUO3WO6rEdryL
+txDgA91rU3LR1n8CKjXYw+yrCUkYmetjKixJwPl8+yNG6r+mZZFyj5RBuP+EUEa1UZFoZRx4u7h
EadnBR7XmFSl9P/3efnhuGPA4+bbgnGQqThHImVtZeH9CMhfoqKyE4q3y2Tv5nZk30vNI28OOpXF
3h2Lwi2RSJXdLDDiDgjBLkq9wfF6SSbDvzC9xCxodsLvzlFsGG7kgGmW76lhXyjxsAK+kU7T6uhN
P6CLVGWSf4VzOk6oDHYd0RdQ91cbhTcrdmIxbRpwBiv5u1k8O/fFqloeSJruqlm13Q/T+9J1iP46
QCKXeB5b3GxPT69WhYehb8YjryALIIygu3wO1V4lI32JFEPhPGA62i/XAfNUlXwhCNdY7EFZXiPf
ampw1giKPBwlRZ8ky+wmaKDp9p8GicE4Ro4685XHxU/6ccxhbsGzaVBMhgacKXTqypMq4KSKH+UQ
g6Hbo34L/C1O++sToVLkFXXBB0C/SspJLhO8ef4ksqhSPO7I4DXXKaw9P8Uc+5ncJ9tyw9vPKdV8
RSb5EIl/sHRn9IhQypJMS9rJ5KeZbsL++oCDb2g6idIkt8QxKwibnuOYayYClWkdVS/GaRrl1EeR
yUeerry7FThsophCEPBuvzMMFI5f8dBsv+2xqyWeZqp5D3mZOMVqlS3NOXOFUk8d8jI7s3oXKS8Q
kWIL510xe9nlWN4bB+uqNEHv6N9WWjLxqMwp111RdJS0+ijrZFGXyK6dB0o1Xt3Vy6YpiTaP2RsH
2pWQDu1rOUj0nSp7GVzDrAz1Eeyi5R56JI4UbTWnseq6L4KDriGsVFRLtt7Kw7U6ae4A3zYKXzuD
xjStL59M85ATQb/XGVjpV7J6i4WXUH/oehtLb2tml9e1HDHCKQRbjdxPP99Tt1ePjwOUsZoR/Zx1
bg5H70SKecEiBPDOuyyrIwdH3Fw3Zx3pwCkK4j25uz8UvoQtu2fzQv6/8qmCPep+hzx2XrekuV49
7LWopMP/LSN93b70OHmr4k+dTniXgVXAUkZ2S5ZprqKunF+BWyIoAbS0xzVScxUywRn2y6Le/l6h
qxsCP5pj/bnPbq5BcZ14D53xJx/JRTV5J/TeTPfwD2OgzxRXwduQ4Qy07Mn/Xvl8Gq/XubSiRsJY
QjCRT/XQy7Ujk/5X4SGVR3+tBa0O+lzcCsnm4PPqa525ulbVK45Y0Ix7Mj8rV+yUvTE0+CqcQCWp
Lgy79CtqCQdCcUy4CLGAKie5IIJYYdELPA9qI+U6CZogurNBBaLMrISZsSQvDElTq4xQCwWAUOV9
FsA+StDDAlXJapdASp2YWemK4aiokAUsq4K30u9kJaM8+JVNG/G9fJoh/T9fxohG5+JcErh7CiaR
v3zhK9wI/Z63tqcPluWjpVPmpQelxGWwxqMc1XR4VSDb8+0hcFyzTbwuvuaP1G1AiQULQONBKfqM
Hn0DAOKfhC4B1MHUNxyPOW2UWt2E4t2khFdcPNHK9egli5krs8CvBvUYFlAvEI4+F4Xqv+15i4wS
deNzMSoRIx977Oh3K8Y4ooSSIb3UF1cDDhWfHNWeelV8jRNvB9XyS8LaMzT7K8NayilEH38tk6AQ
7jqjYE+XO9iDap2jooQsT94ZhkJqa0+tOhS6r7dVhei/GhXLKr+h+h4IJRjjYwGA8hWfrhIfWXqx
d8EmmlrwqzzCwQTswzlwWv/BVptArGUCHawKK5Fgslc0J/ZG4ytxpi+EKbjLc0cAmtCcbQvVN4sl
2jpQ4rY85O7+epZs0wvgatM3H45FFUr3f2yMmqBN+OFn/zFQAAdxJMNHnUdMGtaPIlojHAHjqR1E
AEVCvTkhfxrRt0WB0DGpkmr6tQsfxFL819AapOQOo54Mgr8SfD6WEHe7h9YjZnOC68RUgo58Oxn9
+8gk9VANDArhyzlpJL8tQ+AGISws3gK1tqKitaSjhMjf1Dz8eq63fjdCOASO87hP7SIR6Sz8fwHc
JfdE64XazpxL/fqNDU6NW+rtGE9BvKHX3PtjLQJ7Wv3xggyAiUxWAX99kjybS6nqDzHnazD5Lo8i
aBsHiVSYtPYvVIxJR15794IZAVNvmPMc3ZbLhv3vEGzostyryCD5AazQo7UGvNTGWBM+eRHdUnSg
+mB70hvZuwz9zzZTtOaeslAeWR1qmfP5fSTnUSBBhIvYsKIK0R+igpiDtA2LpCAQVnfR4hQslm/3
Kul6h8WXFFEGXn7kZ08DyOE+JOyTFEeFdRGuo//vgO/sNrXjwTKYqUKVzolNKwgkhozeANEBvCrm
djZECKhTMqehe1FXii5WbpMZCv93pogkms058C2uKpSBK7DZRY60BKqW+jnna6I6l19IPD3h7dPr
w4oLc88PgMC6LbFdshuThzI5kSYWnHxhYbRc9fbu+XYb8LaTTgkakWMLMc0iZyCN0/1qiSbFrRqA
N/+pYHdE+r/+Lqhon9N+w+SOE5Hw1N9J1fksBT6pGLjlnOm2Y7m/Ia7OoAVrOf0kVXJposTj3nKP
ClIj9TnwvLTXQXwlr5DwHY3hYmZfoJlYxDWH8IMhuueV/v0UIZpZHdpwvL+oeEX+aCmvuSUx0pRm
ENnELySCA2DTwlhFTRyz1L9YZppQvCpDkcxVeHIRWUOFzwvaNV6sJL6ikb7YZW9yqFBgO6tTnGxZ
jEfXy5k3Gp1LEKhLozCv9LgNvZebxKCUZJp6wfP3a4vCvHbDtl/0IvZh3aPy5GixZA1gGtt6n00t
h3mf/U39Y4q314h7ukH8uCVjMUUbIGIKvqCuHgO8DipXdvmVWc3rJBEtjglWCodmmoQ/3fyBWscc
H8Inbs0lGKcQaOFj7VDXyI0X7dCvzNXwylPw+xT4Y1iL2BwKowhA0UzgA653MVk01GBp9QvDU+Gj
C4HwTKF+U7520aRICDkWWlKa/G8DjLwD0IV6KV3GI7DLnQAoD1ZTPX9urGRSeAmuK5Mr1S/WVSz2
GnWWISyDv1Ra3bNzTuXReqdpNIJU2c/w8gjPFi4trcjcugQ0ILeEA19iwk4iP/PIqQuxLYuP+8Ao
HduJ9Xjwl0q4sDTE/pJpaFP1z5cVdtO7HMoIMkee1tmE0a+npyaCnDar0HcAqQ4IXo2qTkioeFRe
WswqmaE+U2jgFdaj4qk/ys7peenOrVgbxVhb9kjlgp3XHbi2qI7XCqvCpiHSOgltCtdPeU7NjY40
Z3rOxtvvtm27FSybKrg0AspqWOzxg4q7vX+AkTWZ/BqXZaGkkCEjrGDuqkiBK6MBrZpjzwhgEnQY
RRjF6gdn5cRIG24p1AsEhI+CZuLgZ9wRjt/ysFinHLd8xI92HqPUElICNkJ9kd0GVPyv5W8nkwnL
jjEoNaQIau0KoYwegIo5ZYcle7XK1DQtuRcpJIKZbmrrqAKZwHcZYlG5Ts9gS5Wki0NSYDj+INr3
/EZ/2OP0qzc2NVPompquxYa3SItrcJYS6fdy1qxXp/+0GpQmmpwj3jZTWDySdf55kKserfBhRKXg
m6WqmdrDOuzPHMFn4F2Er6fSutUZR6EsuTRFYl0MtP4yNkF3On7xIeCOdOET8Q0QdPK4+zwKef1q
lhp9A+ymslUTIENVASV+hrfheaR2WMBrDAQ7xSRROMRuytih+z6K3MfR80LEwhh0DvAsVJTB7acc
sX/4kaXzV2ssWF6FnTgpWGPowpQaWkZne3moEtUdJpk13K1VfbYZr3SJg8QAzqP6VvBvaZ5DgkUe
1d8ufPEPU9HCnKctRTPw4KV7S3MbFESHl5rVT3+Trw7QHeFFd1CC7AE10cEABBEmKxodQcGqDdb6
IEw6d7ZjOn6kqytY94cHt+NeGIZZ1aKdtXpV+e8bipFPkA2p7nwY7BQ+us056McvjUoLKYpoL8PB
zOeNnxHhpcNPiPBrfiT3kE9n+jPfPpT7l1euVVuYCSHsoodlX2O7mJPu3Oj06zycsNQ/Mm3c7tVW
yFJWAE7JPlVhmNZOVu5YFUJ08czgimgh/WBEenaLFMB4ORbWTx9yvzrHATcnTxxEskVdMInbRlWt
rDhMnNbivtZZYajnDs5Tbx2s9peZ3jv6uX1NPBjHmaqpzciOyUm1x4Zslz5cSmdstE4zWYP1FvWo
4YAI4rS5SPtZGyf3BvWT8n9+KlKr07DsPc2Cs9Pn/btY/e0VB9cE4Ljr3iqajnDoWag1u1pV68UR
jKcr2OQvqQ8B83Y/YLqik6XrabS3cvma1PskQxYfcrqbKl7gvYFufL5/fR3dC1/PMzfShf6ePgpd
0XetU8bhfXzB3IAniWA9yyV0SLDny2fB5fQygKECtEio3+oFNiMojqSMa1JvhWEOg0xIUHpcuXHA
56ptb80UquoJf1GwxVoiQRk0ylGXgZSh862G6hmzaoDI6B2WF/kgm4xJhi1HBMBofrymm0wqX1+c
DJIHYPJbUodYH0v0Yht0lmWYJD+K5fjFFTiUOqXhuv9WRP9TNPrZ5XY+DbcplEm+aWwVjrlYKj9Y
XzpwReH/lbZcRhqBFBIJ0EZo0vwLkVMuMA1Pdh2uJ8Fg2Gi4Evyb1IZEO6u6Qu1z/y0Rp58Js+DY
SzRqx1SpMg9hzAB44V47my3Qh4fmjT9iZPxwRpvkvsZ/sUe68xvgAcEFTx849fMBIhvEtzUxnQA9
iWK9j/+7SE+UsnRPWW2B4kiEUqP3BxuYtE6Y0ElbACphv3lX3Jt7vuaimB+I6bMEL70mG4ctBTUL
puwnTJruYQBE8V7+FonauKJ/v4pW8QHwgsHXFWU2FjxH07eNBLt12WNoHr1xQc0HBq/UJghVqDFN
EVlLUyfhpPDFFaQz3ToEPihx22rbZz4FWNhKotToaYCUr1LOAr+q3EkX6UNw0b23BC/oGkkarpNO
aGsp/fgr3yaER0TA4i3JhAPfG6hUS68zYnQz3gciLfhhfOIGFrqpN9yOa4vCHieXN0zgDf8EGSF1
fRm6uZ9uhAlux4E5/0hOHeHSBEsK9TJS2WZt3X2I51ONPO703rndJZ0Ld4RGQxdg4oKq4mUb/Y9C
USspMpM3UO5CtT8gi5NdEU5mtGrzWQRtHBoodpK7p+nLtxyp6sYaCgDkb4k8aJSwqNGYFQYP2Q7z
oXOccNhUk3CUBI421dgqeCVmRSjVVajQJVO9R71Ufd+6HD8+BZPySq7L1poT3+TZpav7DGk8cwGc
uk5V+nVnx2nVYtibSR8vbnDYj7SeiHUX0h10QRp9z00QTWQAQyPUKORKeKOFo34gWFjI77aUcxKv
vSvKEfvLqv6JhCxMjmHWZkxE9gvriA1tc6Wpc167NyXe/KeHIkWvOj7oOaCNNO5qcXPLGY1jLpkw
Xcpu9h/ke/3qZ3n3Fs9KiTyaCCY6iiUTyb3NM3RtVXftr6J7UkyVf+q4L41WEjHZLuch2RVz0RF4
EH93ZHiOuZMVrd/Xm5I7Fy1sKhhMCps4tlSv4OG4SzkQFhscfa0asUggufLrFYVqTbqSXw52EuRw
rnA2iruKB7+yBQ5eaTRBzIzO4zRUXR7qZQrvdVREfgmXih6iUPthnBqwApHYRqr3M21ybNVkipX3
jtO1YkQ9jAuRPB43g5/5wLHDAFNDzMZsqBeAzlFI4AngSeAGGeHkd1hxKFDhbok1jpYig1Nx78CB
FcRiAxt0TtTzXKKjuMQ828zFGTBi3xsRMuIAdikU+ikFm3X922r4T0DLoRgHfA37OzkFWlzjtuhK
B//4GXpSC2+jiNm7EmH0iwIj+b/TOFpfRLQrasI0edXq9rHq035AUCH15h/jNoQD/nVDHOac+alk
MTgMPDsLXXz9e7WYG/OuFwZApVSY/o5Zg0hrZz9eT0rA5Z52d/feRV+AOq0DArvC0g62Ly+rK28h
rTWA/+9hQMRCWXQR9q7fwV6AJ6HNBpSE+Uh5SLI+Hg6uaiCjV/RA1qEG30GaBwRiDeB7ZVcAspSC
SzL3WQASHxayfSEWTaQPMDFZqbnt3rbtKZ+yF/MlWqs1NkrbzvbtsF7t9KWCuYVjbyB4LuekFPTS
U8CFWDw8UFuFkeiB4I3FDTtUkZFBXGyr4IpaA/wKOIqmWJH3GA9heWZyQ84Hnc1RWOgVJCpYnBxd
EGdqpKuBygzn6o6MUilYXD0UbWOxC7uCWhFOTcAoDOaT3uwnEvX+ZEDVkVxPoIaP9XpmBwdGE1ON
fdoL1Lo3VNBEfwJRjzyoS3cDmzE+HAPyRav9CVZ6sSRIzdSNhW/sQqJVJpj+rDqNLysiCDNqH5Tm
7ZVoYspFhKTX9CE1RDmF2sNLlSYN1SBnZau1hkXaHiIeS0oKNUdNWItrDgM3z6UQ676P/sosChSC
SGCvDzn9QGRTNF/HcxZRXpc9wpP40uwPvtvvtKpP4NVRSLnNMTkmKJYAHghSqSrizBTJBxjcdCWP
zabK1W/q66/FwZ0CRRBlLUlMMzySaqSC7MiaLN04YrTK7Eyh/QxdRVkrVNN4EFR7VxVLUMWtMLWv
cjSls9j2R2l4fAbl+VOTuIVptijbKCR5ZQv6xUYvFt3B73buVrfQ93zdvcdC0xfOAi/X+K6aBF6Q
COfr/NmrnY3QwFPkrC/cQMJlXezsWvNci+D1J9oKwCoTRYVAsEuAOcSrkz2dimbPHv6RyBAV6HfI
JX3YBYkqui5uo8lTEgrUv5xdOjlZvS7LaGKIc8Hd9a1pl4zgDFxb3jCxURPR6/uo2VVSRhUf2rpk
XqvqUMtfAbQjwmN0dvuT8atbefrvQ8bLfkJIPPceTvLKWT8EfLvCnqdok19izuZStWYXizkLLSni
vcmUBauhVQ16WSxFClcP5OCIGFpyw6/SbCHWEjEPLTdVVDjZv6dcfWobW/w5a519oFjidys7lpWv
QOpDZE0H3AhQIxYwTzy9ip+s6V4DBw7qqtv4vDG7ORJQa/8qBU/rnWoDi0ycHejBPm2o/IpLheql
Su6lb1Fg39BsRXdjgMY8GfqLdESYPCSZm0BbjYK20/34kNrgADSq+jm5MXDpukMCr5HlCoa4Q2qu
+subaVFot26hmTUY0f4E/4MxOhM8yIOngc+SuWhIDCJzdzW85194PjRQBD+A1dI8RaBPtIPVNp5R
IHPxmpQlLCRY8epgSVhMMToysB0sa+0umjsviI8wA/LWwOtIB1Yw0uX5sWgk6vRcTKG/B8UQh/RL
HSBM4qseNl6UdiXnxzl4KDM1qyPny3uOu5ZyPLW7PK6eulVkqNXYCrECp3y0tZZLEuWnTi1GH+KD
8iEOj6epx1cEi2Ey37VHkPQEwQm9H6AOJEyuRCerFt4ntjEiLTqEHg5JRCHAuSh4wBuFudq6AMd5
/ygYCAaueabReB4f8WDhS6pzhynPfooX3BejV5qnLffyUun28NJNuWlK7xIO36LmtxpCgJIe4Rn4
J5ID8fSxUilwUOr3/Pk+wSQ4JMiDX7im1yfyndRcGdg4QQmn83KZNV05yTfwODDaJhwIpeU464Ur
rnDHcjCBSkaglYfdADcjM+EuBJ6dnkUWU6qe3aJCJCAHpXuzVGLKnFpEc9caoRLmOFKocNJX/he8
dpur10zgMxZKYkA6MFjEjtxvfoHb/SgFxpVPOzmOiKMEIRZAoOUBKrxKzknoT+PsveCKTd9RDc4/
e9Rw3qf3xqAJn4uOzuP4xFqowVzCcRkfgToQWNo0Sre++9PwPZejUnu8f1aN1X/ioJypMKLmOBkP
ZDoyUd1jgc9Wv1eRqe3XV8wQGdN9xl778OQf5L6+pilvmLN9EU4VrBruSQKXjANhWvdvwALbFFFr
fkKkR9JqWM8GQGwUBboqisc6NuAXoGFEb6Smq/V1LD1N3fY44wupgX4sq5/ln4plOl+XY1bBs2kx
bGlKi0w35kbmFDO/t+8ukHVCnUmHWlk12naNXQ8GlxyaMF2arzEezlkixO2DV8DIw75UoCNEYA5P
ewXz6Olb0q/RK8DVeS4xUNAkik+9TKxcMm2R6BfFohG0TG+1J9F7Bls7LEK3gokWpwiSNdNX66KO
5PsLHG47A/obtl5j9+oa5Ghpbgh0l20+eOvvUqm20nDhylbGQN+tB8LxMbM7D5uXwpBf04ikCx+a
GqRQT4F6yeMWGMZvi8ZXrAyKMf61E4Ml60LuJonGHe++LuSEWZBB8dzsrNx6UpRLSwHmctRsQwK0
mDaplyYWSApInBuln/ioaww0Jsp5LHEK0rhHBXdCPnAoL6lb4Mm2twOSoonB6eoUnZ5Gy1CCYH4T
ONZt5ice+oGS0zzIUfbsmhoGBctRv9zav2G1PMtJXk8O5i9xv+guRiKgdYOCM2jRymFyqryts1HP
IbVtRGO4FyD8PkgjSDjdOEDRHOnailolmY+Zd8B2alOw4yI0K+LwrGqKipOw292BktP2MREQTZpt
IMmma/T5JLBzRLZGP0HLNMWboK9yE5Ry2F4JqBICKxOYoyrYgfafNEOHZ8WeqpWaMGWflPWJi2H5
5fQrKstqN/BwsB+o+qmnnIin26upWLdmWh7Kd9FQzX9h3Py/vQ0DFinMYK229EikqnMpEHckws9q
CglcLjjSRX3yD6VEVsE7i3i8fBe0SV1yPoyqtBnFziq0RtWKx+6iFbSbtI0yzzNKI9hlIq56rnYl
yJAd8D2c22BDqaAMq600Av/C1tEEdxymYpZkxnnJvAo3oa3ZzDEFfs8cyONOXUI9HNJB9qsuqvck
S5XwLLYSPGV/n/7Uxuh5NIUcy4RXLb0tcyDgUYBLuPsYT+mCPwmdOZobJrZsf/YwIFa3slCStlCf
jdT0vMPYbdpMlIPbBd1+2amLjmaclUEUtEBGj80E1dQsYr1BuUMHyYGm5QYC6ONH3scA7ZzBruQv
thLExdMb2YX1ZyTGKqK7CpgxWSxpr7hVt9FxcesRxd6Tt73Btlr36SSMudAfcCanj9WIm+Uz6x+F
QTlSZhCHWHnqr9N/aPw06P6Zl4sR86MIfrIWevBmd3xE1WL2y6ASv8bm7jdayg3aLDCi2A9/bAUw
42afByUg4ZqeYs27VqOvUIi6pmggoDg73flurqAsqfZUPIQs+HpFdGjkl9h26rPXKmmkkFGRpv8L
PDGhh/kO8swYJQNRWqEfbkK0CXO3GxwBvqfp+RZhocjsKcl9t8YopY0soHQu4FlirDFDhzBcQnld
Vkw3rDjjTMeZ+u7ba9kd8QlrFigzWppCDuw2hL/Nzw6sw3w4l7KfmQD4OZq9ztHwVHKaD4W6Pdt2
1bh68MheWvkRvS4Bu/acha3WuIw2GGwvx1XfbHhOyIdO0iWq1JZvntdbpifGWVQ2R5WlENKtjAMr
XyZtU4pdBDMm2yo/DJPnqB//moYAJ7TqZd76EnYuHknQdS2ZNS2u74Tb9OhvocPdwX0fKqGU1Cwf
Cl8z1WczuBI8V1R/Zv7oN9Xr8harcpOEdAAyLarCBHjF6sBudSE4gkju/+DTG2s/4munTr9aor7u
2R8JIdV0Avdqu/V6lcMgxV9nD9aUpiHi1v04/dQBuyC3AY/l9tmOc+mD08+TWuCmX/smTlV0ZpRW
wFa/0qTTfzPaYyqGqslkZ0WGlzFmw0N9+WdsJG1PkkpL7b1WOZpSlhXcOiI1LhGfwDiIk53sJl48
m56EJfL5UJ0wSgxU6gpM+GizvNDNDiPP7z4wq/HtvEPrHpv8RfNWLbOP98tCbjbl2egHr/vO1/Ak
+eSptNPx1Av//FA9KmafDBvicRXF5LQMmqF2sg6i69vP/H0hj5uDoDXXe/ZmT9YYizc2zIM8VoZu
YITbtlcidV1Zpy+puYX38HiFTBAspommJ/jWBed9UcuXVfhghf+GPkTsIibRji02ex6/f6vE5LvG
hgtbPJUpGIf56gYZ1Js1KT3652tKZlPW29IzuFOJcFz1ySdLyppwLhCk1wDu9CAlUS0iXE4pxush
Q3Pn3ad+KirvTcHLMlV9BlKYnQzm5MPclzG/6PsXHxzK+FcsYUhM9yc49cybexAu3IYvNMRI72CR
U+n58JApgBkT4FLx0LlMKVWlAcaSu7X35ovqfCxrdmaWXG143SU11Nw6UubxU7/LA9KoCbGJTuTF
SbR6L2622BxFoStvkpc/yPFkHIai7vuG8IYb5WJCsYKKvhbLptF1LixROm5b/TlVjDiY/UjmJh6R
qqKGyaM5VTBniQaiHx7Jfd4ewS4WW8sa8C3jjQ/ZBpm3FGxO0EOqYyH2xgbs+Z4RncwC7IT6ePEn
8F+BsiWB1zmKq4EYzHtMEjtYCdErAC24iD9Y7ckSfWrzC5f5TuUDuKG0uPUwpVQze+uEkLR5tNya
rqr9tubi7ke1ppirbwn9XrXQ4+3grO2kXsxpqVNv8gN1BbfpSztsC7Gktrlusb+/rsg/haN1hy1n
tmT2GiyRF8lk5QBSvjZxiOUjN51Nk3N89IKuXBYgKmvqUco8g22uP7ds3bKnpK9QbbwBVR/J51k4
ACnf59iTzy4IKZYwvrGVRzmRHqdwSgNaqJntG6XxIa7okGFGYwbk7KRA3puQZFH8bY4sdkrf2UuN
CYdbgndKlajA/IF+6Vrek4O/WqnIl1O+BgpeeuRq8zUvGomczYa2U8jCbpfnxsrjmT0/qYNeLLtI
BBmg+WXpkBP32LVkNZ2INsvdg8lY7FHadu3iRdbVLtPL/MdHV9kPnYopSGrFUXvbmVYAeHwX6oXE
rL3owlH0V92hOvAzHk8mRFsoXQzrj0tuyzA4mzgBzz6FAEvTXWSEQVOBuFSv/f6/TFKPFgbq8MB9
tTa9FlinKOOIJCo0bD3yhc1nfVEbcgK4JMbo24MPnNSCKGApfo/aZ41osycRqdMKfHMseVFLUskf
gOc6jVSmYCZY6N1cto9BbXCpWfInbWMlX4NSApalDzlbSM+UeU2+ezfByfLJ+BS0k/sqbKO74vUW
rbXRSh+o9SjQxnDL93O2zvH9waT+1qRTaeOMToPKBqDQ6a6seUWKVAD4pe4UwsAyEWpjwT3BZ5dO
rynacQx/R6+kd3rSb5PnkkOLQe8h8nCZyFFWySExG20Hk3//gYCXYdhdRuUgvc16nmmaKXrOqOpw
wl+uQskq4lkEqzIQE3wj4/7tkLHJM4CJ8/TsOOApk4Em2SSmJVzMJ+Q/9MIyxpDzSjNF87qd52Ce
cqz54tHkvSrpvrEtJ75Y79yQE1feKA+mpSsJWrtJ9N0N7kRdDTmtR+maNqk5F/CRWv1tirv4KAXN
hpZ6TkBBe3+WKbBUEcykdHtTk0wafhRSCDGALI6YX3QP7D5hXJWnL5rAcgd0var29SOlr/ZsHp7E
lYa5SHNyXx11pPrRr4hVHSbRwIgUZuTgNyPQTNnASQ3SJsJVVW646rkllUdymgJBy9a9yLvqqwK+
C4WH4xeGfglXUe7jihBsUWRItC8F2G8koj5Glc5nq/fMCulUfM/TLDG3PrifDgFUcPSR7a9Kxf9X
vThUaysWnIjjzzIThIiSlIGYPF6xscIboSVNyh+mm1cjIO/h0fQAyilqXxOeoJrbjN/XRsEPDH4c
ITXfVllf2fIjkguleCZUtQfSKnmHVGvo4iZ3zQAt7Ql0s8xtMKrM0jsw8/rvyK/mqAlhg9hBcOzK
QAJQVUmOphzzDynHJjp80qLsfRFacVG9ssDtZacHyt08AKN8hya7Z0uKuBDL7qaKudfu9PO1bFnW
Oin1x06WrplXsC3BsC4L4F362UzvN0qm0FAcW2EG2inHQz/bvzmXHyQnqO+SvqZfldpd7rVAEKpM
FJ630gop9hrQJTH+ePwWtvIyFtC1HvCJKL2JZr4H9cTrDXNvos77RDFUs8rUbYxP36kCkUBPwMmb
togFVF2xisI2lv2CNsdacV/1KltO/Uys0iEimAdMWgFhRCxH6dp0sKRCVwRkNNL9Z64cWka+FvNJ
mdPyy18gW6SKFd+tbSWp+MZQQX0ebBDhthiSNeNJvt3F8WsPRbMXXg7XG6mpTPZ2qgUuTZoZ9aqp
RBv+TODalOiQZl0txAin0oDCsr4kB527c4P2SIkKVegpRZNDJIHPSs+2S2tyJz5a06piat9KsSwH
XnKH9QfbSRBBa2JdLUvFPrb9KAiJeIlETIO/+olYfXxhMBFoE73HGDWd9bAV4z/6nW7hpijWJuCn
TvYqhB09JbbaOyW5KgPO7p8X3HzVOj55Ya0Rjpo6oUiwbE1iNFo9qREZs7mHuKeDMO4uG6Sd9tkg
ZzfNxxQjRIifPJT5tLY5B8RLfpTiv8qltY+BwAT2JaOITKrY9gPmlQOSM59T2H4NYeEfOpjIc/Qn
2deROSr2DJhVXCAASvfWVPuehuW54VWtAekPt6SCbhW+WUQVxRjrY+f1R9htRe8pp8ek0eM4OOXH
ERKbNr8I309OnhAawQAqcLm+UilcwDkIDdGM1fkewY9G0wRbgfbzicFkec0oa/bV1Ekr9ya4J8Pl
+wbDC0/6ZjkZ3p4DE8QMZcVVSf88CcTrYJqrHCnjSRQtRWNxm9QDaXWtEVW8Nl1us4qi5GHKyoMu
qbzQejGrdPYmmD5v/ioSUb4coBPTTCUcPvlyfRkxE+qca0JNUrjDuwS6bXqXdcLRMUEZhd7KdykQ
5pIRFYNQHNrniPhokMFyn+YRBBYf2c4yoCQrjOELaJKX/94BfY7IRAJ+NpAGCbdJ1r5ALGWw9yt9
ofzFSjNOeHw6mqrzqBSzhGqmS4yDZB36NkbcfNNOT8rB76J48BGsxKopOG91krgkkeZgJndbq1fA
gN+3KE6NeV1LNSZ1inDbfR6O67FihimXsbw8C0X47fh2DqxDIpzPqYN0BhZpUBOFCAbJJlB6If+A
HRLkoXGGX05wMPIrVjJE7X7DRB5N4gtZvpHYRIbz6ANhnwT2ABtLhmhluOZcZYdEl/zek6S9ciJa
bHrBtXE4AreKwuqoyEPaKTDzqbkfBhzZ4zkSfyvWnrz9alYmZ7a9bVt56y1Y22t4LmK1ytsdmt/P
OIYNJMBkh5d1NO7fPUnSw+EPJSkdwvmmjDJobr+5Av05pxx6ugF0cqNUtV+rUx8RQwYjBdfHPDUR
bErNfJLBHw1lo4NlChpUl+GVsIaGvh79qA2eRRI2LngvR9ub3StVziuKxBleacDSv+Kn6/Ev5wxr
+g4WoktWdrsneffzwnrvW+Xv/Fec5adqkAqfm8H6cfMBmIT/bVYVEknvaXsLUmC7Wfh7/qwZQnYQ
uPjNLjGouRfAFAoEyUssRachnIz4bYm4CTCleaeG0L6oRzLJmptSFouJQKuHoun46T+KkJvBKsYX
Vjrab96VWBCGpBWDZHAC64FJoyU7+rk0irmY3UD8ByePX4qwsm2YXc094qeA7cGQ7/aa80INavE9
XAalUuXEWTI+O9hZwy3ttRx/FHEztgVX5qxFzOLJEieithzmgEnBTUCjvHzfRU1L9O3arYccioZu
WBpSMnvrlsUaNCLOFmZnZWb7XwPKbJmpTlySpbJeiLXq5eJ9n6GrFYHCHTkV27+h5dPOyf+ad85r
dklwxvR/xyqGTTyZKEIYHPxZLLMD/328lrAB9N4A3wQgOQOfayWzAs75X0JDl4LfXR9J8n6kj4YI
3PuE8ex4bvkZtLBw8B/AuD3AeK6+dTQaDx09YhhyKBx8NhXnmG0NhBN3IMRn/Wbhm70RZXinCHe7
gr6He1bY8iqz5aIn7Xq1uFjl2y30Q7CmLVH3Y2zfavvy53WOQRWD6YJA/9S4Af/9gtKID8oIyhvD
jvq0E4jBoXg7iZRQmT8qlBzzOtSuk05lz+RV5tUX97X8i0V5k6877jolaeEgTOtNXo75o2zEyQDx
MSvoIY0wYY1/9q3js6VVtyad+MZp3l6k200RuHSfEPBPRWfBiMUw+8ciOiaMYfif73EQeoG2lDBf
TOYtatoeHnIe9O1jejG0ne7w/H8zphsSQRkr50mPYgYOX2ydNI/iwi5sF0P61itIPeXcW2earseW
TjYTqvqakKOxdGc7/I1AxZ4z8s3pKxyf1pwzQhM2ru5+0TZzeYfo60w8FLe5YmA5lqYNla+M2iw3
/TIUSTKND/CKox2YMJzhoRb840eXcJQ9Xz4GN100qgPLw3oCQB+2HIIHNhUbWrQ6FRJFP9DNxGmx
W2aUDvHizfjybVyGLeFqrnYopXCrnr9XAflbeeq2PXtC/gge+hu3oIYN+mt22e5siRv5igHsIShD
uyquktu7KRLLkrtHyfp1mJSmSZnBCV6dEDEDdaEd0cw1Xx5IFlHiWfZc0luc5mfvsHRXsUiupY9F
zWcpLYu5DVYea1qgB4+P5lhVpDpWc7NdAzkFWqxei4WGjHL7/Vb/fksilSZlMBIAV3VDelNeFVli
xZoBufKPOutzKWTPXJQ9HxfGYNGYt1c3vFN2CPj19/E9ER3oX7xVGtVoueSQn6BfuJFKX8HDvJA/
z7SY+JT3C/hR6GXSPkW7Su4GtdwYjg1T6BL6VdjO4sBDFaZWaQwQsm+WO7pNlHGBtvpVFJ2hFbg7
wVnaDrkizhw46jv6mL0RdMln5dzr9NoDmYE7jver/QV/BjMpxp/dulo2osD98ysZ/HZvd76kXnZc
tUEkMiFmWCu1p3i+rELbA5gWJJ4h8SXSyKKA5z97mnoEdWJ/fneQ3Mn8PEyxo33jNSL4BT6hXt7S
ZTOC1TbNpuwI4Y+3ovkaQgNzpdRpVuUDufMXp34pRTS93L0h6/rtYFi8Dd6bA+JqoDUViqo/9yfC
LQ1N4MW8LBcwoFnwmiuAYOpxd9le04/iSVSTLSr+Al3cVZEB9mNb3zfX1qruqXI4B5vuy6vVU/0+
HUJfdjjRLZdg9BZCA7W4uprmp3ELWfCUx7qDdImr9DcgGLBJiRSRvViTotFdbLjFdnjqN+KwwwM8
YMdJ9Ea/wqLJ0Zc/FelV5FSk21wnCVSacJGgkl9ZVyw2lLnahk/4T4vIPEZ0VKpD6BSbZYbWPXwy
2XU5eO/E4LuuHWMV3nzUJ1veAE6JSFd2K5jPb2LPmD9wLGw88Nttnc+38/6nh9A9fi450d+EwcZh
OOvhocG84vlDrz1pLncGeYKCa1SILFhf45VzAuLLWV1k5UJkcKv2bGt+xCAgdkKqxSd9GPEQaF/g
+zZMJ9JweRqMIFuuxibjn8i7Z917cgdaBQX1gvxYL98qB9cMtoCbRIgwX/oT2QEP4FV+7rwi0Bmn
V54uRHQAb7cG8c2rXijZT49oo/qecu/g1lC1hASZRnZNeHshP05f+Bt+VwH6Vb785ElNgJha+s2J
xCj1C4dXjBMXORpHujyeMrWPUWbZWGGQ0QVJ2VIBlSljVvQRCEXIPVLDux1JZbIEVsqWDOoi+FYl
oHBtUnL2x/5uKHIPo3S6uyNDpaKjXt+ujrxQsHJpS49uBBjBACWZ7ZbIN0hILzRRdd8l9+whe93C
iJa601yYK7p0TjlWnZL3IlL8r5OdRTe4NcjtYeyyksA0os1et69NibPFWNJF7sgFhC2l5kUYfjSn
VdpAdYWHo4DOOv+ku3710mMmzDq03OnsWJjbqj3aR/bk2zLrReQbJT2tpNhu9VwkP9BBLMCTb0I5
hMOkK0eM24xRDn1ABobOdnpQNb0myvXDe3vHY6wptPz+sqGBjwdYDDPWNPSKFh1xjhzDIp/jaQ3T
F+NLFDEOH3kcoDIS3KBtYO7LYYfzZj0TAp8dxHDUkKeVvf7YGlxe4uuc/xZLYX09OXORs0UAlDCu
GuYUaNdrMxJMCZV1PNlbbP47dnWPWM/QWXo0LhEJdAXUop4u9iwcxlemx6PT8Esbu17puEyR8T0/
n2jHUkxa2lsVdYKgNnX/O3Su3Ypxjba7Bw16tHGb4ISsqYokKv73OoYc0/8BDKrA04tn7MuHVnjv
dYf2FN+9Og3O7EljchtZubaCm2tc6ag2mVrJJlbOwK+Di474FavB2vp1rpcMl1Fl6TAMuiTbQBN7
KF0UFKP/gGNJ0CTBmqRG/a0ikT1B5BeUBQVJHK2BpXUPNs9GMCQk6yUQATq0wzGS1VoXOBU/nMdE
XDj1q0LQ5BIgHl0eI5TxPyzAyeyyn6s99UcaHwvBG9cD8xMKiW8hyPZDLM64HPSCglWnFueQxYpV
N5g4g3dR5otu/CDAzQwpbPcx7FDDgDwXcoV2L11IrNS/5a5fzCAb1UEWDIxrMbVYl9rLk/99VDfO
gzS3T/t55WW7Qv/+FGRCassf78Gi4djJaSacE0gGqMAKcfedxZsTb2llf8sHueFL2W2YoX+yyRtA
kJ+mNH8va/hTodgQ8lBk2nVe25tjVNxX+HF0YcCoTuQro9geOSiQc16xnoTBuSk2Q2Wv0cfXl12G
7UxqIBopPDmvOkg9oSVvzopQNS04ZaS/RqbGPq3MeRPx2BrE0S7bLrRHchlJ5CHFyHwekRFeFaZd
YshK0/VtLxv6SXsPTqri87DuiLD/g+b9OcafXIhV9P2iIkVJwPAOFwQlCsP5/AeqJ1koIxUBpVkv
Bw602xDYc2piIUuHjMVxVpjFogYLeD2uwPD9p52UFRlNkrZfZa1Ytt43xn+kgm5bu392mGYiCxFS
DYGi6o3hnrszXavr793YcRKEiKn7rPOfc3NuOQYra1BGHWzYvhXzZ186y8xrD+K2xqJbk2ke/TZZ
xvtG6fjRzmXr5SnghK1DRsSCPiwZurk0fLTgt7xzT0F4lu55Zj1GeFzADYI9BC4eUzF8GhdyswOd
B21IJMI0vonrD04/owtbOBYSoqS5Odcknv7mcShfi5n7qr2m3Yeyz+iJ1KSXqGG5JdeLlCJxzS99
ANn2ttoIi3oqYXY4+Sa0BhwNVHjpn58hT1LUKz36D66Q81sbUeyRBs+ZbWGqhZxyJAy5KG58YfM1
OB3TjdzeTt3qOshfVwpNXU+r0NdjVckn2XiW6mSAuYS2hwQgSB7D+5Cobg3XdyOPfALBtph2GGPq
1oT7G/UoNxmr+RivZ9Aa9AJv98ivVSMSl/klNgSEtjsOYLc8nn2HFpRCpzBQ+1mZKYrIZxr5hBbX
4iiWiGLOZ2EkngkFPnm7bT2zqVdoMIEamv1hx11VHFrhC3GMZr6hnZO4YXzgVuGxCkqiQxSJ2T6f
URwlG5K+pzR/qwjSw8LbpSXNejix1BAJaeIPiNWdqPxc2MVcuvwRIXBCLBJMew0+KOU3U4u8Q2Zo
1q5NMFH/fuGm4ufonA5NF33jNjChmEaKnOpr222FKZdTBdVXfnnXL/8sF/5FyzHugaBvPwSf+lw0
K5yNQOCl7uSbZklHv1eH73jPrKFQ69phTxVylLx6bQiuaRP39waoquAL9+shy/lIsiKLjY5qHFvn
sMkCQLIrrW1CWG3gk1nLRobsasXGun6Rk909CQfd7y2EJpq4RW5+x9yD6fZB5Q1huhlDCJyKFyTB
tcGIfiBNopWY9lLbSbTUiCgj2jxaYslG9+ORDpXY40PORkIT1Kv6H7vXfc9BW2uX+4EhLTWL8B4u
kNKjeUo8AlNGhm8OGMQIX5Bvmj0Vy1Y9s9wVL+GH9WySgK6z/04tVLw1+V1ekC898vsWT/4G9uyR
cHFT//EZPC9fqNuggulI+4MWhpvDKgyrBDwIExtXoQlXdLJeZmgJmXdewybqwhd7xjRbxuyFxy32
IbvXQ+L6kf9WJJBO0MuZQxBtAxyP+tTU5BO6Gr+P0g5gq2nyKyhvCSQbSNdLsQDrsq5HJhCqJ1WG
CrtH4py2TnRRExf8XSEWIkeZ6ZUn6bYo+5tpI41IK1JsO2/NtUNguBRaM0nCRJIvA7GUeZBucqgM
pgDA4Ypck4POYU0zOdcmddFMUr3XWh37tQdtME7fJuy5r96PQCDo/5gQUr4XnM3ZRgAb8I2aGI5C
q0VX/oTcFoITS9vkGsFCTBXfQJjxFOH9E5ybWa8s1KY0k30JhoxUWPOprMxCXguDnn+VGID/+gI3
gTqIr65Sciu8b9+i6E66IlUsh2p1vqFVb5SXjmozzUBhmvlg+/3L0546RW5C6ooETnNnY12Y86/S
ehgq+gsegIqbUMyQeKXRExNIavih8AtOiIllI41iYEr9HWaYsOxavrW0S26f1+MQL7bXCsiv1Hz9
rXioaoc0xQcGOrAblyUNFWFDHGBGA9Uo7GdTWGObIDNDiln1HLiUj6nRnT4MfsCZqkaK0DV69oMa
i3FHJ09wPwnf0STpGB2NuCs05cMSv9/LcGr2WKKBoAaD1Fb4oZC8rS7cD1UEYy5B4be4KMxCaxlK
lg2nxG9ZTJ71kh58slPnCPkQO1HuC5NFYZriP1JiBoSB7awPC3gs1Ot7DnWpZyDeATudOYPuqseC
xzMEwYvel8NdqZkQ27jSl8zUDe8xQKiPmIJam2SGxyumm/K2YGY3vqp/QaOiaRUafZONEKtMaPtD
RYOzlSNxV/0VhIbIBQl3sjqJDkRofPWxtPPrZtXO/hP4hma3i6CzOZsCr8evIPbO6smocxJY9aAI
5lKF33yauVmSBK1lOEDSlkh8cU1XWjNaRgVnVHWTAtFa9oBWT928N3xJwiZ49FBfOvVf68vbuFzK
+rsNr8u0dyI10Vi9j5vd3EW17w3v0hWThsEra+Wjg0PUQu/IhNFtPxMnEzA2EtZtjxSOpI2INMQ6
T6P2gQZE/qxqjk/DrJJ6RdFSBDePZqN6WROK6zR39Gii25PWFQx57Zy1nB5zXsKAMafp6f8s+yAw
BmprRnbVwNkGtmOX56SnUrGruJKCDMAE/vUWTArmkFPsamzUy2aAn/t6F0m4Sg1OpT2I7Wm/asVh
4PFSC7OhOCwTqBA4gM/TPdUxOD5W0XGltHX/wI8Bljp8W6hbZjKHFNALalw2Uw0W34bKZCPQTDo0
+mQDCcaQU7jpCeyAajoqBFZxeq4LPbGvaNYoS4+qQcWkBiq/nNkyiSq7H7C/RpMXf/zR9uGYz/Gj
NhXViZlIRew2tRZ6sfFd41hZFBvhP3gSwMwQkYTV9PZkHpraAoumVrwaPFZq+0ce7P/j5jumCXjr
4+/cd/lP8Uk3qQQ9th1exmfNYJzoxOKn1fnegKP9l5IeLppkRBZ/zR4C3CV6ZW+7VAUIwzh8dk5b
Ode4XeH2ockZnB+xgyuxRuh8ZuMqxzAwcdY3b1e3ffXnF0NB7Cb6jlFQtXqryF5G01ioWGIb+k27
cG8XpLZxdDTYvpbpuW1jKe2yzwGWO4oU9Tpfx8kXtrmR7LmhdbWuP+9nl7Ws9/oQTEoYd+jUMCog
K4TwururnO03qMFH0k5hmII9FnbNt1EOpr8ho4MWWlKt9TM7JPCjnhpd1bhpjmLAjhKtiZdbJVYS
OqqYU2JS+K/0DTDDuIHOd9BaCRNlw8FjoWo8qJuqscQ/uZp+jLNxKrPz3UPKyDdtyRWh/axCsWdc
KyfwKO610zVpZcJ16JPE5WE6sUkT2116+PDbZqH1GVrrBUjd3Fsxe7Lu4SZBMlbciCmwIkuc3io/
028UPuu82tx0FcaP9JxnMT4/r7LJdu2lWZ16VXQ8hDn5dvCBINVEmrUnhFgTqVGhIzxleZ5Lz5q2
E2qnzLs9ynSBiJw7CgXQYg3gdtVm+d8x9xjGTtEHGaMnZj6U3citFz8KxmDwrTYDedA56PjV4Bo+
J819U6c9IOgZmVDZQk0U85+1ylpoohJJalcBwWQPM1F2YdhbjS9c7VskO/ON755qZXU/HmPFD0Bp
305y79H20rnI7ZK0FGLO6mVP8ZngO1guHmP6GsrQU09uk5t5eXYit/68ei3dzLfF87BoAPa6qhBY
yHr0E+EzjG5Adqd56uR1+4Tdg5qHlsR14BnZM2qd+AJiJuBLssnBzrraksMf8olV2n5OZ6vzOGmG
hOBNyw633yXHudwosn9x+9eOOsRpuB2oGccqSSz3USCx5I6Ja9aSrHelBzgEYhPWdgvEOJpTeza+
Tr0OxNxtgKWClRii4N69PuwO1RoWi4HRHdvQy2dMz50uJR9dMXv1LJ9oTwVv4MH6covCGjpGlMJ4
MQJsNRxx5YSGyGJGDyWtU9GJ1+XfNFNRu8NXCLx5jHyBQid70nMZOGyKEfQhmL5TWRWzWCp/3+Vj
P4OaoKD3z1LMXVXd+FbwB2jpwXJlOFjwr5q0f1Kh1mAz+bRHayXbVPlnVRDK8+HB1HXtwRGig1Yb
iTn6b7pJ1SqkjojxNwCY19GU7XTdCxYr7A1IENjEwL4zybwBCDbwQzLfl9F6NrcBAZ+U3yA6kIqj
W6nCdT8ozjrNLuHv18FYO1uPIQ7BPHJ7zEw4uQvSre+pwmL3wXiFI87QW3IX2c7NEBn2IU+GrzRa
qQDZwePqGUJl7afbV6lGiY6sSPK+vAmwIBpnmVEc2NXDVy7JpEJ7iMUq4IxACROAu+zW5VqOYBK8
acB15rwDIjQWTbKYQnGm8lhOdYHxJB0qArdR9K4VAEKWhc3zUXEu3m8Um6/M31RfKaN5hfriHFQz
zOCb2erYpOj9gxfYa6J2rlgSfp04D3QCy/zos5rZneGNv8HJiC2FYGCyTLShW4jdOtFbldoNeezg
fTLcQyEp4hFCJ/JicWxfwFxAYLL793YSPkIc5ACPwFwRBkoTRsRlnDsGpLM1RRmblHkxJ3mDP0Co
Qa/DufpgngOWCnSTE4geo6A6bEI/4WE0Z7D+h0Qf91YW+r9Lq8UFs3b4IIz/wpgdQ8HbA8o8SEEl
1xGcdlnHde51hN4vT/2T4R4rj+r3H72VcHdMLvSIh468n0SaeK1ZXv10X0wVHgv8eRyCO0UBV86r
uu6GeETajwMwPHG36+/CG5EzMv6eS164lEPmQo0erL4QOgu3yTvMunNfO2ty/1S3bVkhJesbEutA
dXSJLy5kLfu5sNDpS8YvWqAo+5Pp6741mgENhmAingFTa73QtsH2Ixsc+we8BOBryLaNqJkbfavX
1p8txSTTVCnBW7ypKSM5WYRNGP33ibRzQCgKESUdG1S4TUL+mk8izPtIlnSUiJl3v/jihACBb/uq
zH35nxm3spD57OKv5Mkt2yZTusKsITzKsHjngEJy9Ay4AhikqKOjbJm9sU+Y7pnyuTt4B+THf28m
gSQePFuEwspVJr55cblFbP70I+rCPYoqNnZCMRSI5JawxdAgCm0mYVBt/IfmwNwPG/znsc4tZWCQ
PqUlaBMW5tt+17o0QLJpAjpjsKvshaWK2VIli3pSRq0/X/k+5gCb8Atri4vpT/1AIfRjuTvI0SyB
UBaH1B+HMBuLi1c/iXfQydkZNO5vJJ0pUo0lTVVag/JxPAbfYKQuxZdARFp3mqnjv36+2rLiRLRW
hbVGY1D1bF/hn2BECPYUy09IZbTnX3v6oy6L7giHj1gzF17q65a4XvoM+AMMVupPPIORx59QgCM/
s3GGcArw7PpEkSgYTqzim/Liy1wuAGe/abYapgJvTgS11DKwgXF3+gVbvFzz5qc88AsIn1NcBytm
EKlpLC2Anb1E17cqoN7z8Q7XSa7CdqU55q3pYrttfbQDlzDy+D/1b4ND5wyIff6pkXG65aIpI9vr
SAhhmPs66rqDDmmhFz4j2pflMcYC6yhpr4ya6Z6Ip6lDfySeQqaOp/e4dMOGB9WXseZYa9fXi2y3
hKs1F8ms4bAivacO99AzaX4p7oOr2k+8sCR5UmgczxeW1sRwdeQoWnYCvTKnZqxA7ckJG9xuOTce
v8ch/pBL5cuHzWcENUfSckckP66mPgRv4raFmte0q16mPCoJOGfiDe4R115q4BGwXAso3HAhgb6C
HccBFm9YQMsWeqBOjeMJOEwD4uJZhprGVbNKxvfxzyn+wdDUFsMaqK13m/2blIWoXK02/L6zdyU3
Luc4yfpwuZE8vXLKQsB9AVzFH8sw1XV2ui3axXq6kPMVAHaecj26qZHsb6s52Rbez1KbRmh5VroT
UEVL0MXfwXXw6/6ZYDVBriFuLczCywXoLrohTHo7EubZzddBJgAeJgZbLLt+db4hjcfq3Y1vJ39n
Xh2anN/mIXyykLqsLLPtKZGo2H8QhXce2IaK/9KI/haW89cqH42lBTCP3tqfPOrsqChoanZsMptQ
to01EzglY0XcJlb6u+MIUormioqpEYZwgDbhADeRHnoIuWRqdar4Q05nPGB0w6dKGSIpf6saXwBD
T8ouf7J53igDy+u6NlI3FD7V6+oqptOr6ChNM6cngZOWfsXzlv6/Ag+iJVVE4cszfgqIRBL018c1
LeELrScNBha36RNScsplFwZBJzQ5AePT4iwMc6BRPCuY9u3RmyjmDlsFOTacR5lK98YO19i5+QC5
uYcmA0HiQnQ9lwq5USuKpfdfWYmh/pLiytdwa4dRdpA6ySbqiq9sqta1KHVv45I2LBVPwJ5bQWTR
ymzfMtOL4fz3RtL1bz1QnMzQ9KubxByyIp3KNko0yKvTPlFJDjBNFmSSuTCGyLNfF/lePcitHHVI
a7415GUXK3igssW7hGPX1gtSGhzys2JY9ufrvtJL2K68msxkx7aYbI1o/hWew2ycMk5VKbROlSiz
/dxA1ULHl1OUOnv5+18C+7YpjXokZLl1kALl1/BORXKnqU+Fb6TPLy+6fqncIqRLqM2biFhchxRD
SWxWriIlBWw2u6BfzzFaHAIRATd3txheUKjk7QHEdgXnRTpZxZBKtQWpMzX27y0O2BHotP4xiz/r
euQ/+/bYbCUF1RzC0I7BMUfwS34bCBnP5mw+ZDcP59JyDn2dly31K16kfXxVOZOWOb395PfB++TD
YHLa2s+ky6m+vOSI0kuDxfxP/IGcQCSf/oq0MScKdpZxdBHy/4RcDduaRMWTBWEpOQ/qXdfB280z
cKoRQxMtwSWp5pzedCCrH4FWUBbf2Dsq4/oubuhW4pAhzJnCcIuPojiqhpSdr3pG8OBfnTLkL24V
Z5WFI+4TSK0C9rzvJ5vDGFoInTNdcPyilVkrHhb5MmBW2tENrb3529CMj5tF8vfNa6SZ5M41YiLM
wKIe5h73p3m7tjgn49snAULrap9u5ze11/vQEC2on2RwegheAmj2HZ3B12stezK8/huIQPoCaJkG
oWTrnzM1xVX32GsfYQ2x2J3dNSIdhOTZrb7Xwfor982/oi3eiMolGPk6X3APcnmBz9737PQPPWgP
g6kX23g5grz2qaxsWikTsftK0pGwLjHjnZi8Cmq/Jj2qn0MPSiPytna/QlWOXdoyWeRvjBbeJ5EK
GBpsfKi7ObYjYL8squ4c7sVhUnHV/caaBmjyk3EBuxYgTsATdTsSYXrvV3nk6DTKE85j+vbHXWTD
9w2YKKjObNiejffzBxkv8Xxk4IId+aeiGisuEeZ0ZZuLMt/3wGW0ivbPQtopZhoy/9iXwNTqp04Q
cSelB4L9E4XcsPp1JU9NRmNVJEd4WCfc/8eD8023Ru5qxn9Pl7wR3lKnirPoNlpETptVwSuK/j6d
BWM65EIa9LjfGWboB+HRUVcURwS7GWMhrOrbpTL3KAqw4YmnQ3Q6eHSeQuErzrZHmSJVqB3y3KhE
RqVyAgSARhXdM22oXKHff6bgHzp9jXMjunwQq2MmLVWMGlobppwATUfLq+n/32KxrGIlJj2NcmZS
ZMLyMbCLRn7hm3rIIshaS2qgb8qsv1+ew9TgLENAoNvXnSOxUsT/aK6hLppjCmdahT/AhX66q9tb
MdZEF6HCI/e+DMryxR9/U/W1rMdm1zdsWCGRhVygYU+PBI+yw+IW6YluM5MYKboKoNDnna9wa8lW
zBSKVO5OB/bePUoNnIibsypeuStdnvW3+i4RQW9PYggIlGEy70Lm/+UhnA9xTJweVez+AePFbcqO
Rsu4X5n2iBIKNl0+jNT8pszV0ZCAkYCTwbquW/iR6s4FscfvIboVwd3wlm+Lh/ukogolxa1SxL++
tKA7Ri3ItCYVFZ1oSmgyQ1/dkEdTKBv3ZvpCN80ZREqrEe2lGcbOonqByQDh/utwZL2FFs1EBlYt
V3UX+CYelfl3q7KKUXb1fWn2b2DUXKzg7gfo95mjuMuJ9ew9GPb+m/+i7FUWCsTtvPdA4qYSq23Q
JR7EsmNBVhh4N5jgm0CMPTfkJJ8jH2G3rzpho2u7ps8TZ8QuOqAUGYy2ERJNOtc+GLK/5ecvqRDi
vvwjNWZxoAPhR1ZXDfD/0RpdbynsWGm19cilwthSPcn92gtGLsz7lCsgimQ9OHUPaEvZzFOmUpqe
0HB3LVDgHzxDsM0NcHMhgjohIejQnrBgj/NaL0C3LXdxTTfjUWk+mijW7Tl5X74h0kqm7GForQv/
lSXavD7EYzJdmn24yQ8EhuYa1JJM3AN0eWyCweTMP1r3lrm3XmmBJnJgug1dbfOb58avpBA8mYJf
ZmDRHSNCFJlVfN2aGs63MJkPCS6bWAUdx3V6wyMci/3rGyOSEXIKsSzKOxEfpX2Rw9XnuJ9It1jy
MG5h1cIpbxDxlz1DUAw2D9Y8zNZkmn8IWF5SEElR225SkNmVcsdCmbHbm7cbPqDncHo9ccCXo889
uapKXbmfBYWehXOReWa2gnK/jgVNzVYuA6banah3IRi9WsorXqnzMwupLOB60QHASCguBJYPnZT7
9nE+93dF8PwRmcQ900AwM9r/cUmy/8eccZXwd7dJ25PS2CCVJGo5XGRSWv6UeLD35shoKPcHauhc
y41dppHVJADJgRcN3/ExKAFLXNVGHbm1z4uinVUsIaX3bpjKCY+LLkwfreATLXSC/6z9L+Mjhk6X
AGiMihmG/U64dzUMyIGq63Qng8/EZfsRi90SB1HHAC5u5NLWYvadsjxc2TVskGKlaBOrS2b595fg
XHIcNXZZnZTxZ8Kq1XEVGVh/UBqym6KwlM1Qnuppwiqc8a3Vnuy+F9ku2mSnLNxN52KZRrSDeSa2
aGI94RL6TikoIKV4yxKCTSeOFdHOILKUtRN5HEN/3cpQcrXKxRsJIjudtYd/BWAZU9W8hs3lX5qb
xvdkkqjsivfbIKl+NK6Po/YwrajwJ6zbVCwTwstQKTickAirOdeIiHIWQIhGy7SqW5s3Fxc6EtpU
QamIPety3gYcCxjfrs9EXubWHRogA2upuczME2T+1aAz21+x+fn+0YJc7n1JGpYdAvlh/acERlBv
2ZvzPHjnJjwQk4NuoO7fJuA9R+qXtXrM92YsMqmxeAq/w3ASO3yzIoW85SqCfEeDVF+9H3Pu7ZDe
V7jboktrzkJK0awC6ElTOJ4j2KamvJ6UcmWGdZMzKCG+kJUuwrAEQ6Fe/k5bLyZUZbbMC6QLG1P+
EuIE06QxpQqWMzkEsLiprzkjFbMEqD/6gDIJzps26mLNLGe93wGEu+JP8nYbE5axXtFyihy6jPPZ
/mm1YmatnSlEOURQx0Edlp6/s2R0ip/tN2aL/TmWSJeaWzDsSWyBgFfxT2jh9pkqrNBC8p3Tp/ti
V9/Ir1XQFkgqethUbCua/KmutK4pfuvZt3TGy7DISACIjuZqsua4WVFgtdHSF2kUCatnfZHP+Bfo
9gV8nZGkD6bPW4a2oZcs6IFjPUDRu46CqgrQGb12ZFROY9UuvqGEViuDeN3ompNBf5B6Q/JJA49U
pC7jceYtgCde0G7WZABhA/tH/rkO/NxcIxoDKogJZWgMoy6VQif7lxKod56ZHZZe0bHrVuKspGCY
UP/2or7LiLwDyiF/SIwCB7ftC4f/SekFZdTCvpLoSXbMuCPNuQnLgRrlgigJkFWDIF/o4BJHquVD
uCVRn5Ql8kLzmwAq3xCs68dRxQHCgPEMflMdwrW7aPPKxgvhQO3O3Pb7wTypzNYbvz0+D5FSIwkH
D0k5+Ue8egfQ7fQ5ooyTrhbkfpn6uHMjDCpGZLXhrGC7gsXCApM6ighXG0p5qTJZHryCmM7tSpH0
oTSUUBiSR+iYuu53mt0AVOJCmYjYDObQGik7DpmK8+8nSPiZvwgkru3LWl1evmJxm2pJPCZPOfJm
iQsJtK+ZmwW82euVVf8tbIIgaxhc9WzSidnQyUlR/hCgTidt3NNOCPDFDNxMEnJBnYwAlMs0DhsW
QFvC8FQtnW3pKAPkxSl5XOk/nN/rgXDpYvYTThCHCBeYO++JHG9PeWOxN4BHb9KkdmgpIYDNegPB
84gDp7y93lNG/25wkw0bofCJqMK27Qy2aI1ajwfbkNWtagXh50kGFuTUXqNVaP+jj1FnrWAU7+m4
qLcHtmwvRUbtSWnP48Pzc4farYZ5wLQWF8Wnva7iVoCeYjXAe7c+gXGt1tTrK+6TjTjQJklPfSf6
2G61zRLEJkSZ+iCtPpAazXdEqOaWil5eB8WZoKtjYVql64NVQmF2TUdGTxAuUoRJJZ5B7c/uzf9q
dz/CwhTEBoh0/B6OOLBz6qSe8XClRKwD8/cEfns0xxSfyyDRspnsblGkMQF/8pWu5Lln2ONUXNCW
wLaBHaOGQJogZZ9WYSCF0V70HKz6Hm35aL0BDfGW/56k3ZztlOWdw5a0nIeKueCfu7dAuSyb3MAT
2VLkfcgkNmDGEn6YxMWFumJ9nPpVGPmEEkKtimOGAaCT98CwmNqALcEifZBi1aCa1wSuSQV8rUA0
QqZL7jIEQQtkX4tjJQ1VyMvvTRruLVu5mozy/mmuZELiS8iso6ZTLoSX2eX+GkRV1k/47c/FM9mt
dW3SIaQolylJ1lKU0XZNNMC4Bi6znnCw1EifbnByAEbGhKf6A7Mrhb7EHUNX9Ho01xNuJihNCZfS
YWcmxKyJOoin8KRNlFgvHkr1mngV2fMx3xWlyrapHQbpcy5DNsYGtThhHI6OOJTy36a9pSn1Z88J
+E1QXgd7oLBKVuiJ4jq4xhaMAqkPyVVIqTS9EmNbyibmnuZklRnNOusMml4yNYZaKoZr7fIlmI9V
HK5IskS+WwacVvrELtCqJb1CZqzqKF4kVTMPxD+atmyiOmhlXpGqwMAXPH1gsUvkDCCds0GLrNsI
lTUTVZFwNdG9QnphwZuDWY8sgnP5cPLWWETmuJT6/JtJpViPwpF+JhP4yn6GxyHoVreaqnI68lVH
DKUxo3yARIoWDXS99iB2ECGGaPEgXzk7fNCwrmNsWWNgwxpHRYRab5QJ6Wg06WzjOB+rKqqCuag9
QuCKEEQQApnu5BHMHbfabVNay/dlgwuQUNXQFV9X08pe7HNXzZmQrotG5j3WdCQCwNcy/O28JN37
sqbEV7h6b5Ua+lAsp9OcWU0Pgw9Tckp3xfEzKybBw4Q75DV1aJhCKe/XXvxPzQOp0Sd6MDo52NOm
nLTtWbrvk51ctQXIzW/rpgbIG2OZjG2/Mq56W5DcbaRmBNIirTPo/zR2faiIvtVXiAO1WmcPsdBv
XL4hcRHUCuFRRti9Yvsskl2q5Z7VFoW/ZY/Wn9/cKWrYlVlNjVVVQjPmIC5rM1WC+AjBFWfcVsvN
6XkPqJCSuJG5HZ8xaEzO89KvvVfznIZM9/fW5Nc3fROQ4RZChXrwxyz8Ctx5Cv0WH66OjcqJBDc9
sOfiEKi7QXr7tdsDwCdPD/mcNi2UgaS2F7wHhEPdOI9Kg4JWAmb6TyYiYS3QxjhExHPz7cLxRU5C
yG+2lqr0ltbZrHMJv/oJ9iEy/J3Z8wWshydrnu7Gzq5AO2eyB/RkkqScq7efYPdqW7VitteJWvsq
FTS+EguVOTrqLijnNWNk4tipz0b7781fcdSeAMrWQSW237EZKdU2is5Ov+uRG0vqOrq1bAZNFb7V
145Vrg74DJ2NNFpgxB3lPu1qUlTgqd6V+cCP1uRpAEXMQBBm8U8Pp6v1xe/8RFdv9DljiWir/vz5
zzJnxkBRFNtHfXUabkqoo7eTxjCBngXEJBm5okAcwmJBvq6oxL8SMBO5TGgWbDFvhpdBiy9Ne+1Y
q81PaDQ8X9RPQv1/GdN5kBSNZzHp3/ECKVeck+NkXrDgPQFXcr7A8YJK9lxuwWzJ2dVxP/gtCwKU
54EilaRKZtfYfpK9b6/lbOqLEMF1aqzY3YsETinHM3BjTLlmcvQAu0ldBi6dGF/sljLgaJuK14F/
KZlPG42CPiS3dU52yU8KPjKajFRy/r31rH937p3Zf71xiNSr2eYt+P+Y3G2T8NntyLKI1QahR9aS
m2coEGGKoAfynVVXPGrbUDJga276W5Rn9QOPz4qUsbE/bswx4YPKbDynxxqoe3CIa4udmjReSza1
ErCvtB5PdpZ5mOEz/eKKy9czOJbaD5LBBGimIkCfYqvfUHRi++LPiQAHMcZzLie0awsodMHmF6N7
aaq/hFYFfo/uVSDivkannXessIeGqln+a299aVs67ExNdcn3NktiO4AIjktYmFiE+GNIYjTu/ySd
63ZVTqcr7+K1FJBjALebNPNiIbc4nzx91UoZAlg9m1PX4pmRfvg1cw/ML+Q8l/6p2UrmwgmU2lbp
E7WmXLSKaiqRN37vr1vaISljG2UzNqaWcSmNbOLndh1ztmG5fPQ5ErotkTbm9O2DapvrHJD/enTe
jNAZGuomSMYYJvBGc+j6fsE1uyjzfBPVJAXKJgUPeOF/E3OKD4YUClOCyeYWCJXLVcUMmMRFReop
h0pix7nm4din0JnbhSaDZgI9IlbW5y57JZjm+kj0PmeK3OFN9Iz9a5nxK5GFwbJT3+2D+cMtvKP4
d+fqiIKq+rJbK8qpIVB8vCap7oNqszINZh3aZKHEtgz+unRJsiPnj21sNTFDQAiJruI/3Kdlkliw
ELmDLy/4jtLSQQ2AMjBCOylkbUkGZLLAfAfMWPJ5vAHKjRvmyH3miUB3OYc0D5nCs0VTLtc4Aq8R
VkOscnYruRSQkr7qJXFouo3/8tJ8skMieRxb6SO1ovHoueLa0fq/KLvNRT/EXSOs9RYgtxJE20Di
ACvLFZl3x9tP4QyNZKDCc/Eb5+q4URH/v0CpCbx8Kw6YzvyS7nORBo9vfl0TSwi4Jg9OhciD6EZf
Zgs+32/9dE/nsiKEZ/aXut0bo/ENQ0QcJuKMt+4z+wZ4JIebVhy7H4NzVOboQndkbPtRtgpnU/Vt
tsNcRcdymymQrtJrLncNgehEIUYR/LmY2YLsMvs31YP9awCfdgcWhxqZRjldzEI6KnP63f6W7Yx4
FdqPZ+lBGYhoQ9h7yXttqnnQdAf99TKU39KjXv1LEldngVlZzJ2snnR99FIGjnLPIxWufzKXG5Il
9ZFnJ8bg7E0ruYRdpSzb869OG+P1R3PTpucItwZHwce7QNGqT+BDOqDni3ZddfgTgUCWC/GWeb3o
gJzTrJ72oDeWEgb4ZhQWWaAwDqb4mZILh93c8URckuL5+4KYs5q2pxhAXBmPL9JITd9B6qN+wwlB
6748bmkyWawxt+ehmGVfcxAbEaFoZK3HGD8AHnwFAxvrjziXmtJMF68mcctgNZZHroJWBRWhS43V
daEZl+tIBFax5aR3Pr1lxl3KY4NoxClfgo0VyWQw/eABPeqjJ3Lb09qXKY1R+RSFox4tDlsJzXle
oUBnzF2FwO599Ch86nB5ez5dn6I99E80FicaoM1FrmgVSKfmMNLe7Ks85XJEv4l7HtXhEFDKPoj7
rt8kih1rYmJ4LsQKXRZToCfDE/ij/Ku3D3bp3QwF4itG9bHTI4OTj/F1FIQBKlXjqTwCJVTCdq5H
2x0qjp5Yh3rzR6StNjehY7xEp9EQ3tTSbCIWlnXHF32V/f0K9AeXnhFpPz4OUzldPhFUhOMlKrpL
KiYVk90GE+RZ1e4bzRsYpyeenh7tE2Da7tXg9PKwi3dAH0D+RpGwcumP8q3A64vkbVoULKlmA7RR
XXg4MuXwrD6XmN6fUBfoWarbwNfidcava1FQ+GPYeX1H6aO70vF8R8facIkmIe+27kwQ42yrnJe9
aqjNXEUSR6L2SgYzgFIintQaIugKaN7gnNGMV6c4R6TLo/i4MYvLuNQGOeX0zRhrSW82fC8HXUTp
JGrYS4gat+Q5CAgTRCMkcFMEpDK0z4ctw6//p/OojwdM1Xnk/ulGLG0lOtPrlDDtADA/gfbHG5gG
xbg/TCTIqA8yjkePVu+J83en61rIZz7VkxIuw7goJ8l79ddAZMvJtsaWaE8Ckeb4lxkERzWJPKI5
Fg7Z4oGcoCuXt+RNByHfanBtb4BBk4QWkz1CAfnlpDBO2ZQfxeS0ujFyb1Ulwf/JEDqJamPOzSXF
KcRHiOsT05zoVCEFMqzYirvUQ3ueRlOzpa6dBsmiP6/4r67oije+UEdoRP1UVPfhV7oE62Z2d2vM
SCeJTgnW1bWN2nLAg4UMbWp+hnJO7cN8CGPT8Knxv+it52p/GyMMLtktjN+1/oRzqZqpk7LBXclD
BBy4ZMzbw872gOMIl/ICn8SOzOHgRu8HAVg4Q1xlawWno+YQ398XUHfnTFr8O2P24BQhGltBBmoH
2O6KUmeCCvgMRMhFRY8SEpZZkYa90c5HlLFJWxPztSLVnaCJCDpiU+8GE8iD5GPki9mRkPOUrqmK
9+5kyiZzeYENMGE3/LzCyBokcs3+ueZV0S3tAqsOcy1GRuwbFIM7mnY9/zuUUgl0sm2B7g1nEIvb
v5iWTa5A1qx+k/mGKb8QbRP6U8JoGpBfGjoNu0Iu2MnZp+MhU/K7rZUfesmeO7sbZij868LkmN78
D7cB6Zh8ciZksUQzzOtSLTDoiRWZ0K6HR3iAK76WMuyDSwuqjlMeD4Z+Ej0I6MQ/kjM4s3Xrx156
DMpjhqKIM9s4SfLOrU2phxYUl/jUHRJ0X1GQEIpSLtgiot96kd4YPXbkv5Xw8TXQDiJPBz3+5lc3
LyWtXi7yqUP/d9kZhKEb09FFJaVyLlLiH4auBvLTGLkV9d4CYWjkm/DhoecIDgMEAXtiMYEXIFtg
h3cssj7jXrkTIZhOCKGUsYk6v7ek35CHes0Wgb198uZAMCV9NRalnybIp57qRT+JNP/+1J2WHgMv
BL/raf72SiEqs4LdHUQNjMwIb05xbw6m/XRXrehd+01R9FgjsBCxN0GejAjAHZJMvCLsA3Fcaal1
skRQ/Mg1HPhCCo20gSW15QqlD4W0QbQRKJNocoCUJG1jr8tg4bUvMMEY1i9QdnpUBt0I8W5aCzbr
dLSII5ocBQpelwEdN/fD519GVfIxOFItkucv9UMD3L6aWT86BaJMAPfynHdzDE5UpABr6iCVjQPx
L+v9Xm0gK9FMW73QJgJzi1IEFcetsVzCyYx9jt1Q9bcudbWgqkIhDPJO6Mmdp3hnkgpr8f8dPI1W
nTAKtFmnEKIF9vzB2VHjSlumjoqzZ/O7x0UcIpQ8mXHjGLURg/9SZdROGAk3wJhs2qF4lc12Kf8/
HHnzQWDXf+c95k1n7BAOwNOJyudiAxY8eSq0xzzzB/sMpD5au63xrAteAz4ufQZIrnKWjO5rgsLH
z7CRboqUBaWlx5gEiOmvpXydyWMio6kC0HsCbL0mPeQCkd/Orf2cbk26hWcVudTPdQIo6RUKZcIR
XfCMV+/NFyplu/WyzWPZzwlQ5O3a2rXRJNLhOF4Yc3vjhOf+OvohlNrdAM6FXDA6+tNGd2YtO0U9
iW6bCBpb6c1dVFewNQ7qNfv9HzHWyd376akqUKU6CwEOQOMA5+DoZgZo/VohfD7hcwTkjFDrpDlS
XWpxcn2Hbnnds2N4qS+IQlYQ7e/C50WSBAQ+xdu2qXL4JbkxpmYZfFhQj98WgKpanG1NXlmk/0z+
+yWGV/Z+Niogde9pQzXSGU8MJEPDJaQGRhqtwRXnkAjZNp5BuAMjtij1NGD+ZYVEHUPUan+WJkFR
cdLJdLVn4M49Ac3ncWOR/wggS68gZwZREXtNUqfysUYOEuSA9w7KaVRrVuPLQaKAs4/pVmIOXcEc
e60pTnbbLl9KrVbklNO1vlcM5PrTKX+P0BuGy2KpUWVtA7xGIh1q0u+ydTVi+1IwdFhNrcixGhk/
IdV4FWPWvX6mMv6sksE6uJhW1r721UuFzzGUsCH2KbSGBSflvdRc8zjvRcSrW7HYBkub8pJW1dKf
/tdUEfxykjCz6w/s7I1JiqcRU7+caM9xgPbOmHAfx3M8AyDypaOcPHP4W0SXu6cHApvpucVw4HLi
rUPh2miGKCdqpitbFinWYURbvmttGXLNhYZCzy0GCSoaAu/o64vxgBmZ3GQfn8W+lhJbqqbeZCMz
b4jP9+EFQI2uWRv8G6HeB3TKN9zWGeU9mKFZeONy+YvFQ8icIMvROyZYQ5o2anyfWpoxPW+R4Rfv
v/AycrIgVlMHU4j96MZ+EoONVshlFm+LBCaTxiSD6JXsmYLn7ht3QF5VgfAULooBByE2Vvyo/QTQ
sHKuG9jn9xdu6eY8QugDm9Z8fXAh4jgbJG3mXSTj7f1pYElSmZHDhczuevEdD220JHcVxygSzfBK
0EK1pDK+Lab6ANUGmGFX60A/bYc/6rrgqcoYp8vQd+aQopXugXXomsnNd8wJvxbZaAv9ow0EYg3X
PwJdt/W1K1wRxI2WaCTrZ9DY8YtFcr0NXppNpZRByhp0B/L/XlpQ3CkX47RIwnulYfxvRy2mLxrs
J4NTVGBztT53yqSHa9VSAMYZVcJ8L2T5fuFkwSz6IlL42XnOITbxa2ivHDJOP2SDpOjCo0HbFABA
14TjLVEB7w8u5+rRKDvZrR/kPY/lwXxo4cR20xoE+Hcx3d1BDj0AG/DTVLg3tWx9bRKnX28IOI7I
AHIPnpIb1qMUA8EOm9hw+wuLa9qFQMGDMS8EphsgHYMKWTivTvoQXalTsg2GUcSPU6TXg2s9qaNL
u7x0Ke6JH3k+I+vKkXGazJPBsvxaGJHVJa22nr/sESDD8pC3sUJM94TArQ+pWGSbQ0Njjv1SXpG3
5SMgiwSbZacSRzVIwv8He1fTOeIJHMqNZ/ggnGv3167Z16oRPCNaEiRGnmZD4B6NIRBqPRlS/sXj
hI+I5YtfbNsExXsv3jTuWhhj1J0cu+LECkee5FwtK13rZYtT1YVFU7dUp4KGX2IM/BfAMck2QN4S
Mv1tfAmPcwQrigEvhhCJBydjLKTr064W44VumIg8Lo9Lk/Kb7ScAAdD+388rBhEjkS3A2WZSl/Hu
j15a5h4LIcXBGZ/xwGXCFnf9MrthX8ZiNqgoiAheWrWrzy44cLeAjAjQR4PtwdqmYAwwwYdEVjfK
9qaweitNezA8eRdHI5RIPatjClJ15Hk6j/kZC5Y+KImu9LwH6/lUpWO9bOY60G0Mp9MDXwcwnR5+
qJ3u11oqTRj+Qi0ARyPU3+FSbb7G6crakVMsoQvlXjcIU8otkDXQHmjfVzIk9FPV0dOChSEsiyI5
IZbVMG8U9y82zdmtu8VQ9QO6CcUwdB+JNjcfZTUM21NaUCoFbmaWxBJPiYoF2GUKX0jYh2Rd6dxR
ooPF7EU7X9ffyrW038fWwL023ZfIawcE+yW7YEWHhsh7YjJrj6ECXanXT6ZgIKypPx8nHaRDmlTo
M7VxyIZZlR3ZZD7Xpweu7TWgZF9nmjvdlhAPpLJtz/bVouKqBTBfHEEy+b0pkSvh7AD56c829NOP
K+drx+X1hX+cmpqmG3NdmbyD92touu6kqk6ZKF5uXgy2Zf17eP6RY/dfAFnPUdYd4IkbMLn0MLWC
DKoghXLIFSxIpjwVtDkC4Zq2Nd/R74S4kT00jkupKPVVQcMAkyOC5otQ+2e+nJs2IEIfIjs4CQ00
KL+S8QKMP2ztLFab0c96DqXTMYiETY5bno9YxfSPS3Fq5MVsGf+fBCdC1y1lDALCbFkPW6gR2AcY
BgG8SpVACopMSVUCADGi+JXJhzqYR2NlKrzBgTZXAqMFD1lxo3qUXI5T+rdxo5qqbhmhazuVC0z6
WpnQmMyv1Rau2vm/4WUGeUiHNPp4/cZsfSqCFo6Gl/SVP9UAdzgmS7PKy5u8WZnHZy3J6bi0kMKz
4HLyE/K+XDfXoSG0O3n5Ivi9tF8CX/4AHEoIp3Lxy0SZx6RM3OpvK2w0bcUX53YfasRwNs3VYhYx
ptN3YlTw9DHR/I0aTccJxw7o9NOA2os7j7aScskOQdXTFyYYiN/MlMuoz1J+WfbLRHVyhI/g5Whz
XHyKzyYWD0KKlScRSpsLduO8xDpsI0QZUKjkINse7Qn/MYNC/gTB3xTwGsddmKT9dHmIjOv2SSDY
97+I27HTQDPdvDmHhH3TmQq9OpYVs2L+KDUN6/BJs0Z+FotdwVoE7GRFzmN0dGhxFCEaDcdDorNt
QXvrqrO7OmlewxHG0w7uvQIDOwYYdM43DkjPs8W8g7QQoUfFubTFpq05SYalTs9ZBTbtBAzkFwpk
a6i7Arvz7jE44m6Y01hSPHyDFp0H1hJG4pImUdfNpNGu6lBfFZRhK+rzFSGFoy+6o5qrksYP8cIQ
ZQ1Tf56uBFg1ZR4pPwsI9HcvghNntoT1RhCIDyJwPZK7AJyFbtrr9Se/b2atb/raPgaCezeYiUAO
FRKzzZSQECNHLQuA7bvoR/rX1o5Kndh5eGt96bNER+B1ZO0MADRX1mAu9IThXTPODodnEJvvreFe
FrT72JcSFyffOgdIVmkcGtWE5A4AeuJop2eKX4iPDfuH2ajhz/2kUKBbBAyCcaBYwglCyxm9Xz7q
iFrhe4CpcaXRRojjIhOekE7sTVtf6v7n+4hv9Bcv7NBrn9OzcrMXq4xAHNSzjF4MROkORd58O/yc
xUHOMhewFMdNnvBMAEtjUxX2iUPiHgowB7MXkFREJwVpiMcuwacq5mUS4V0HYOTCUdWCECuiSxNQ
9BWrIORmEW0UUVneZduGmWEAz06mhWZ1xDAPA6eBFkLqWcylvmW7lexx6sOegngMOZYeVoUsv0wa
rWN62ORpV/Gu8OAi6g6VKpob1NiJD45dtWn+jbdOJg6Ulx0ShjmZibub4g0bHTCRU9EUcRQGlVQZ
Fa9lA7kYWILHwLswsB5h4L/ZUZhdPP8CY4zXGMQ28T5/zkPZHKVu62uqIXNl+y5OcgQkDKfwJT16
SO6FoHX7YsjEvqF3ZgDPDFsQJWZJ0rPHKj2FAbS8dCMivwD71hRkY02B8KS/bJkGgde5W6PnArtn
41JclEVO4vw4fNkk2zxtFcg4oYrD48iu9l7+8WRPEDJZPJ7AE3oJDUWdXFY/FSfvpWgwBN49+hWk
6ZkQTUUaRkcc5iq9FnsK27IBuZNPSzKnKJSmUtNzGwFlLGLN7L/P3FKnpFoEYLdnskkQfOiqPvwq
946fW+RRkutgnNY48c9g0phyniuIRH9mD0v9pK741UmHLbyZCPbxS3mOLQBn4hLPq8FBQDIF5f9o
OchXPUl2MPXZanPeeo6n/Tik33MXrChDJl75wc2tnlRgDd+Yj4O47oyyY5L7TJHas9HElOtuCce4
TduTIsMW9YnIuA0gGhZfhBlRgARfLg6SsAtzE8Gds7M5v9Inz1k/FOdaK8zwFYM2Jo2pg9KhVd05
UXWPTmMxDg6HScIKy6AvdI9slz1j6V+xNQLpaDWWWlEs763olVtLoCpzYUp2o2VfBQsGTCDpjE6z
eKFZ4v5NyYjkECPWxXTqiM8x75zU180FdNRWpe0PqR4WDBCp4tKtBTgFXKeHDXUJj5mvANGFGE1h
QrptdgqB5JbM6Qb2GH1dMUvLUGfsOhCNJHBxhDNPFple4sm7JBqDoAVXb7vSbaQ7l+sWmYmjjiXg
g7/4MB5UpQBPj8QrUUWjokK+RyEVTU2rB7XSJShwKBZigW/GZvc8WePLU27qfHAN5mZ3BbBMG8TU
yjIW9DnYugZq3HftrteUXEBJA5mCHkTPZM9t7HymqfARMG9TUfj/m7VkbVXKuaw9jr5Kr2/nRNiD
jHzWxlnXVbY2qSSJzB/uUwiEmpMCZ/p/Kj2wsZl9DE8GCdlMGPQqCJf93uE+pSlz09Yxt+UT88wK
WoT03uKdiMr/AT5Vk5FAOo5DaBIh3g64dkVTw0KCJuCuM2mZ1sJM9N2YxpWIJxbRpKEl95+TDiYm
t0Er2aQTXkpH2adrUuqyhV22S0ijpThIdnm+mU4Z8vVZmySDOs10k3OmboIC2GFJxsRP1rRNGCtU
H7lniywyr8MNC+/mesCYNfTe+xn4nBLEyNiEKvtKdAOCY1cidOEdTIuwzgYux6UJ7fpP6NTDMoEx
7vZJF7kNmscYtKACctjTK9bmzXV3Z3IV0nUbX8jEP0GhN3LR5knReZoorIKu52jZEfviCTbYc5RG
arI1OCHgQElz1h2Om7w4fcXl0bhFczmgQ6NXneygm14e8TysXG1pP1Ko6rFA7FuI4wQqizzwQSEV
r+Z7SLgOE+Y4egUTmWzdSvCL/uTfWdvyrJz50e0kT2If5x1PjqsCYoKxziaEDKMOOQiRc8vp3pe2
hzvHuQ1+l0CsnM+IhpKIK+w583dbRtqb9GIZ3BPDJtGC5domDi0bRU6/vlT5y7Vx0br/aO3G1Qvl
O8f2yBx2O1HFf1nn6JchnFc2qNeIyF0xvSL4v3kSH85ugUC3iGve8acz0oa7SMjt8ngD0MoU9ukV
X0G9D5FvST4m+V4DdERO51Qf8d1kixPVCm3k85D94e249cYgsAqK403STNp8+HmPxqYAZ6R87nzn
xa1ksWItxdGt885XPEBLX0AKsseoRww1xCaMt2VS9zq2hZwRce/dMofIoG5qnFcq6Y3vopOxlOUG
3rx00V/ul0rrlu0Qgx1bW1BqQGPObDDOU37jgKB1bDhlMR9ry4O7ZB54wG/bDAKts2gKZAPRkAFA
R9162AVsREklx9TrUi8FYD7AJhJ4A/clbdx3Q8Y4kAwWAIxbcYrwghT9GQVvONwAJcpH2OePBpGF
AxjpC9CaOumhlbS6ZddUjX3/POQzMDF1j2kZmaSFn690Pp9BO5ysEulzILqc5NyZyKVLzhQpFndy
fggxvd4h1XDUSf5qLMYmpHvVGgZ1ZofzqXyjBYu6Au1r21wpPqgL9b9xUFLGSeGwyEThkCuU6C9r
HbAfbjQbKeAD4FNXioNKwx2OgQ8e9QLupKkpNNO3VldM91u31LWSxJRz4G994jmNr+G7MbRchI6l
S9KbIrZ1l+8nVTzf2/UvSEAQomLH/RP60H0sZ6/eUvhfRJvYncHbm9LJWgSbwuOO1RW9xpLrwaYh
XGRwMBnkiH7AUQZI/hrWxKA4rPoH09u9E8lTCcGhzd+EtpgkrzG28eHDlS3RKK4G8SkU4jzkfE2r
H8c8tm/oDJEqrhUj/Ummojl+T128asvINWG/BWdezOyvn9YHLjST5OWYiMXSx2/9VQHOBea2WJ+8
Y/SgbMTh6XkYqUYP0ChJA6M0MZRibcMQYpFDBWIIOltkAgg1q6Ngd1V9aCwphcF1sALaOVDcbbf5
j2vOFxmmAFNNt2KHhF+JOiYt1ogcs3GKuWAGoyOvkOr9WWrQYTa2tC4rtPKDyT3PjHdy3Z5mzy+p
BsUhSbjr9SzaVoofv9m9zf/111agGPeiv1H+wJLxUeWsyQ61pFJICi2/J/tZjEStUns5BPAqkJji
NktVoLCqDDEdUcSvfV05in1/JrKiFo4icK1XE6De7YCMVGuW3lbcEaBShXpT+fEIRGFTgbJ0J+L0
ge2zpHwpC/LWGulaZhb1qU9iime/gO1y7g7xf6eHh4SIqacQ3bxoqpFCSjXyts+lgkYCOl9a752z
u0x63/sCPh0OzX+uOKcgtCGjRmRWwciY21TgLzawEJpOQ1zhz1oD0mJwjIEosEl4Lp0igMuPTb1I
VzXBTjbn48uujG+RCnuhZYtKs9d8gTUGY7xyfliHLZ2B+DbhJa6vZprQYAVBMDSm+Py5xR8MK73B
KQR774aW8cLWcg2qE4qhkR9xpQjhZnMFwJKVuVs0j1P+ONp3VH0atTtxR4KuykGC04mNULORzCQd
9QcqIxzQb2TqDrO6Ygo5uANlIhq1j/04DZuHBJssJkJ14gJAtixx0xXIkuUB/Jr/nz9oHndLLlpv
U/alayvgbvUU9iJQpP7Mo4pvDs0o56XQoke1DxqXbrhY4F52VHodtrAYj4wRl/SM+kCj44Tnb2s7
pJTUHbDZEDjukzM2AOgETsU1JaGaZtus39SRZWFVhjEkC7uG4sNwuCes3rt4w/0iW/zS/bZr0xI2
IoZNucCtgjtt6247HE0tDs88RpQh+pZcA5KW2sEeYBzHck/vpDtZju6dpQ/kS12+VUC1Nhs2FtSP
mJ2OfhEcn1V8U9wIxnVpMDQEMa78Ulqf3GrHThf325oTYv3U8uV7qFPDIxR57+/Qd6ASZpXJBy9C
+tAAojJovJyXQYoZQvP40agEHOmrLF/uevjkq6q3B7uC1mBjvkjOYnxk3khx7UAdrMZrmnPIJl42
3xqMaeHLtoUbTHDFxYsMG8oon0TFLbOCyo3WJdem1pnGqmwcKIsvffZwJUxZPd+YU8iDSGMOYgNi
cV51NZ3VcrkTnqwU2sZIV72bYcy4KHHxmT1sLeQmiCzX2csIqaHPce14rsgrWHhXH5hTbTIRiPCZ
/39j/AGK68j7TagOEqNCiANbHzPAbSfff1DEOcjbdZD2BtKVNhw16sacbV4pJq7OpdCmBo8lzgo6
g6+bpBCmsQoU0/swdpqWWHyL+DAulkb1kPPjQEr29ukyflHJMhufEtm4iCYPFIggThK9qVway84C
RJh8J99Bepx5/HkI83Y3ZT7/sEwRiU367tq34RFYL9wXuvHFAw7euiV9mYrSsUM1mAlPs46vNbo0
iOAsMAj90SguBlYWLWc0yw/zJV/sUjAVCz8C4K9E8nY4D6Z2fLwEIp30PzxI5Z6xdxrGXxguKGwi
E1QPFTnHgyw8LSZYiVFq9G6PUD+QYcrEqYy9a3j6R4DVzhOZIaT+kiXytqDpPS2QVmGuhu3yWlfX
O5r2nqu/DxDZliuIJoHmAZYi0gshN+UxHreNs77iJeEhuSZx28RikfD2nMSgIZXaj9xgBgglicUs
2duNdGAbzNdvTARs0Z4bjDjrULegLBIjztOc6aHKvS4IQ0SFCPuAb4kHf8VtNGpIxLnn58ek61TW
Ahp7F2aJyJ8PVQAI9CuBfWsf4o6c0VTlAbZEVM/KRhW6dppfHfDWPz9qINMqpU00omp38qybMSD5
YEU6EN99JjoXbfO85LKdmiRg6N27lAoif8QR7Zu9i1jR2umDPL0zNG6G6/hwOZwKtwXXsA7d5BIc
Eo+fgHJkboTXd5St4ZuNMyopjTWEP1s+q4LA8WyMM0IKXsZRX90YVYDsppPiY8nvdR8rdju4DZwu
kvoYzP3pgtA5BkSwCYpnZxumix+DN6b83xz4JuhGM2t835H20TP84GfMs4gPZxzyUdnv+dh/Q3Ph
DPrDwLKq5BrkHfHEFY0IYklHRroqaGOgvO5Tyx89tyknaz3TsnUx1i3XNx7pPhWv1DtMl1z/n9w1
A2TFu87/WXkx1ci/9hbYcipjzNNyCNtdHmeHnJZWiUTwAgLqV+5ORfXeQ5+fZlC1ppiH9Y5pVuQd
IW1hWxOXNAWRgFGuSpjvpdlC6hAIz83+5Hay+c2iQjFr1GpGqCQVTu02gdyP5h5S+Zplgvk9wAVo
SQRh29WqVbNuWBvv5OhuuK5SWJ79vpM6Ib5qgKVM3TOZztAxIvgaZ28EA5tt3lDDoWhtUbIen9Wx
CkXVos1u1RJGtCxUanqnUDnSyoWCQdBXht4LymZW5kuAhN09cy2rJpHkzJzAASvB9xLFtcSPJPpB
6DOPMZLPyje1/pFsR+t2Q70bFGthFSPhyZ1m+/txXxap7xL5Km5HOw8pkj9ykLb3G+82kH5ys7pZ
xAftY2/XSv1+OiWHS9VbkXDMk0ZwMKHmtUpy1YG6/8/QZD/IZX694I3u7w72Ge13dLrfnE/rBRbm
JviR2jXJiDNiLQus2QbFGfUiKo8ooAE/5IRq8+AVPImC/sxrAHAuVoOfbHwx9Hu4jEpawFE3lRBw
dXQOr+W2q9zAl6FQHsLwDiFmQt4IY7SpYgVAj3cez7H0JSEkpZAGb4VgC9zD8e0Hiez47j7QBQBx
Ad6SL9qcE8nnICCf4bo2+EcdRqrHC/za7pk3zgzXofgBNFlAc0DP3+qxiNs3N3UA6sLmqwEIO9i/
8Hpgt1t/ZJ5dxnumRBFi4+nD7cKsPmp3jRk1o3Z0gCrSkoUMAZxdasGFNf1mLpTeTeEDwOFaMZbz
mq0yBGTR/lJ5V1Wk6vFzswQ/kNXDCsfNBKYSUT7VDc2953unHuohFM4EU/LUpdinMpTHic/dwFs7
hQaLQwlG+VZWti421Ch3pUcBhDv9Yoa7ZCvd7JUGvuApGtDglE6RWyQdLflSz4XsrBEBhYduJfVD
6IJy1EM/o87uj0no8b7eUc6tPytOiSub/a4dAh+6/462KiZ/4r8n72Ri0G/qQXWuXSAyiVH/cWNJ
vDo0YKmqHFHVM2ucwY5pavUEDuSIQSVop3lo9OKIK7INywT7ATCiHqSU9nHGljAdr3cO2nQYAAkZ
Pa/qh7xFd4vdA9jIKczg0CY2HomaaQcNQXsPmG4gG+z3UcG/iNWzGrajka2uxcbHRTD+xvkrzM/b
HkpN2mprUPQ/x/zMHPuGWyNLm+2yBkHnPw2RkTiYGQLNQQMl7SYWnhb7/iEMYdstvW22Xsf+Dsl0
+u3PjkgJkgmCm6ck9sLazTsEUNNO1Il2aatuyDgoo53FPEm3HkqMfmbSrGL/iAZ4Tcwm4eZIbrex
FoNvT+TMRK2zeNagcD8rczY1PYZ6v3SarhW1zJOtzUT87AxQNIFTuMrnSA2ndArlaDt4pCJJTl2h
wnDRToJwb9TkxntnReCABG7drgpzesN+m3bZ3UZKdkjLNgDzDO371r6OSO7pCQ6G+LOkgRr8WhBg
IAyQLxUTH6riG49ER7cq4Zu1cQMpFZ5A/LUq9ye7fHjAh5EINfHW843IHgTD7PQl0cf7HRwJFORg
lspywOKtaayZnjMXHjDx5tq/qK92i8LkICtUvslu7768xqL3hYyOq5brMM1kYYhgINicDhLn3nEN
GRWsZHKHAXE7sqYnvvBXzrWLR/2eaIoj9ewopsflmQat0N8UNRfYpsx1HxwPpbY5lZkxF1zRPGgW
4yN+6dwJ1pNXj/6O4O/0oM1gdjt4lwpfYigzePdnlY9C3y9GXfj9X37zcZ77UgVA3yNJILZqU5fo
VpQ7GsL507oBd283or0J4pEopfS3eS2kpjXVTUzRUOj7uEZhuisxiIsuu6GlAhU0eq1E8mfM0/nZ
pNxhsA4cQSur9Lmh7U7YKpdy8A/HROGuXuUcB0qO/LwOZrxjeGaCOeZIqFKvpl6bEgx7pcfSbJYk
zwmy0qVSUjTOC1QwsUIEoKAT2Z/FDpJ9SrSB/YjBVxysR135cVeKSbmkHKwVZ1ezInJNVdoOKDn4
xOyoXbQh6nxJsvElAMPOLhUcfYjXx3ZdPjLhhpz4tB5HPlu1wH32Rt/5F1dItbJQ8eeY2dxMSSIt
PpAK5k7/DkyjwI7wtpevf/ms8oZWnZ8GHWcg8+6tDUmbYvBcynxFj1+1GNWRjfDZwiWAkEaEubk6
nr8vfnysg5uTUByY5/kDOyFICMMH/PqydeyNTaXtcO/7KAOnhRqJLyh75o+dDRbUaBx0OlJmootx
bOc1+HtvNd/z/I0jLXEd+G94UvhX/CeIPjV/dWx7PwYrYVB4FZS98RnWpzPnRHlAC3uyTEmPE0AR
swygkjJTsjCqKrOfQK1gWV/sP+a+fHLmOzN+9+2MrER8UswsHec67d4UJ8fJ6McU48MxJvRb4Yzx
tq8Ykksk/9hVTszdUI/gqnpvL5YtaZOfkz7kamxS/WBts8ECVxIS08hGNZxN7yR0fU7iOOAZJXy+
C8A5sI778uP/sMl/c42v/FZaW8yunXAe8a47yFOuQjmKFuKq9K0dQoyOVe/kfBJcH0Uile6ZpRDH
8yNF2/ZZJuoNncUU6G7X6tcsAqBe3JkbzE4RC22/24eKUvF84/ckIR+5xFdM6c+eZgyJkc/TDFdh
h5TxpdCDMS/aZ7zWpbk5CTjmyNsRzDsv52vcWGmmcwTUitFgS/zlI9djZDQwxMEqDVQ3mrgkUAU+
F4faD3Qal2x8wBPq7jjc7lhWIznlJ+kWBH12oFTuNx0wbIbHfEEkiRzJVtsfHbzqJiivgquJGX2b
Y56l/KalnKi/Nm01vUfC4eZTq88FbpxvNoH1KLOj2FsdjruWgfAMg3N3VhySk3mmPtAE4QsClEtj
yo8Q2zOepfaIwLQ1hmV/jj0EH4NbOQ/Oxe4jenHrDpVQpmp2417J9aOWG3yuZ6VeKLohcjNQonIx
IKUEj0MBJJhUx5r7OsO7lBm1FkPcdp7daAB68a+8huwdB64uSH5xy3iqxHRmalLiZPMh/BSUGZKc
XSg8OlU/JBAxOdGUZJd3MRrLCpjT7JNKL2QKtyrJ7SlBy0qRPQ0SUjevGfTnAedYOkEg/HBEzMKy
yTnXlt5mn3cBbDEDn7YSnpbgG8xZxfROkzuToCP7QeI03uFKM8aGCit+jn5ZdBwWxbwC+d41DrfD
SVCiT1Exs6hYF8iz4zGkRQ3TNZdIllY4mp6XMGIxGlSoxYeK56aK+UpMy2bsFb09acfDwU+JR70B
gSSbxhnUuV3fxS1rDcJc5cY2HaYQa8zI4zjS3vnr6tRGw2W3M4Vr02k0gq3wwC13nnVHyofhObn0
jNDpbFtgP5cYTW24pBa0BE/Yq8hHW27hIUH99LUJpeiBf7KQxOt0HYxLt/lsAjaZYH6eLKcyEg+/
sq5ov4RmxmISWfVrqChFBBJbgzcvOscmJpZMLsBK54xZn0ggUplkUVuLfETGr71hee3ZIxX2BSEM
1NzxxuYBATGz/O3WANQTF9cl7vwALGTqzPsTSb1ym/2G2eAxgtUfl/yOmp4C+eMXF0OAUvkHZ/LX
29+Aaxl7hxKnBJI7CCKuuDNliKYWpgvUX8kFf74jJtSEyR891+Ke+86HsOjtkFDD6lFX0jHM6HNG
bwbrxud9hCEfseefD/8Rhng0m5HwL/lhLxj/18RmkxgBYAIiO04r++vz8vsCh07wF1fIQ2t5T5wd
rrHzMreJ87HDLMrrN8z6BMcivkup0BobB/vV1xeKeLZBW70I6Sd0jS1HJgR2szAj983tJKIwW17P
CRu331NUB8PiOkHOeuTnaMeXGU+f9FA1Id3wM/NrJX8sf47YkpzMvWy7kbwCHqv7OTRTwJXb7Rxe
DS1hL4FtphBu5/9f8smPUsXf6oBoXQzeu9jYC3wFC07Fss1ovu/OjW02xybrNU14Io73dnhH057Z
7s0vMBOC9QKw5k2PKTxzoF9mYZNhJMiI2+EHH3KSm2rQs7BeEuixjqV6c9CYzxIvYpmf8V8ZP3iu
ftv7rIQ7WdHyRK85smPzZFEwUdqeKaitD6vPbKk2cctpLTAymu3BMDZfTfhy+b4rp4jhPbt1TYnT
2iUW5wXgUURiUTKWVsD7aHuZJ2XetOofV13OwPmm/AKDSlEzWomLpp/Zv4caND0cRLbyC4wThKwB
Azrkp9TGXOfQseEmpAF1ICxxn8iaEdD5WY3roVnFQpxdnnx/G8pOBLWzbpsov1vDhFDL930FStq7
uTxU9Yl6s8rxBkUDzWzHFtGOs/Aw69uZ65wGgzd1mzCLrViKDmF2Y34NrspWntBTklGVQbBfT/60
gnlIhywDvRdkdX+AOYjMnOgi1xWb2Cd3MK2lKOPAxjcIW3nt8M247enW1DJ663cJzxdQq9W9lNzz
wXxSWbEKFiQGNvTJHSZNEAb8ExdSbKyr7sEbDtqPJ9jXYM3x1PO1VuGlxcwRGvXmCeUZ/4/clB7O
0mW6gohtrT2wehuObshw9SSnAS95jFit28pSHZoHsf+5VnFwAnRyabHmknHE0ajd1TSYcx+TLNCv
QjHeqHdUwRT6Miqzzd8rz4ngRCA8IQ+Zf+CH9UgxWKQgCPHNBqBZZfaEcNK31BtFY4lQn/XZdRFH
5noMrFZLnuPlyBtDqjX5/ZQSD6Ga6mcTxv6acNd1oo2acJq6PmexFdoFWy6UkZhGcufPc0vbNLG/
GktyMcMwgeNZGvu4LqsS5wnKCM3lA5hokhYaSHFwzLwwVL+XnAmOIpkqiSRlNrDd0JgZoPIsTJ3O
qntRZ5FbnaDyQw2t+lO6UmualWX1VG60YS9hQ7ephibasxQAUgWFkQ1haIj6oeMXlYmdMh3l9PDy
m+V6sI/ZEqQe+4Z7pI+klxwE7J5ywOhq1s/g3JTbWrDrXZji8JKrM2/P/qIWZg3o+7Qt0w6JuSsV
Bt2ZOVlLT4efSb1AFzRIDpJeGFMu5rwuuxLTq7QzGYglCfBwEJYGW0060p/jRR7ZCDXoFmFAk3NW
6iJhrEvz0gH1hYsYgB+AAmO37LPwze6iM8kxux4MW6smMhSoPi6S48j5wUQveTH6+nt5VV+07xz1
lgpDNeFJ48kyw6R1R41IelO3XQJKd96Mb4QPf5/Fg4POvI/uw82sIpaQOKeS3duZ6Nmj3N7EFXCq
v1U6kgt5/5lYZGTr9ETUshQFajHpkGAgpaheT2LIM/gN67TPCLpQXRcMWyFUR3bqaSecFW/PCzJ2
tfkE8RF32Rw9iDYafM9wAkPCn6+2mR2zjEX1zkVK4oFE0A4w1mk5iZgU9DeKcUpzYwXqO0xA+Fig
ALY+D3FjvYtwpL5OgpiZq+xqHER5emQYbAV1jBP22c5WZT+6TvrVj+wqqYWkGQ8cz+ngCsa1VQDf
qCpaw9+HQjxsPCp4VaDZqup+P9lDdjo/ja2EZ/4XKah+KNAyb8f2ElNPSLwbUrF8Kg4Kl3dVVk96
he6P94gmW32ha5FJikEzT+s/Sm0/aZFhQIl+YQwkYLd9xKBp74udoiNh8g/qQEEuQN2PcKXSVsrX
ri1A2pm/x7HEzpMLVOIcNZWvNkf1E+VIhen50MGCziRdw5NAqMLta4sKp1C5EbvA2Ypr8QIbGNNq
7lHtNTlvEIYiiKEVMXXnLSYRCOmQQstUJWSgQgdF1BoFrOTUdmqYWW7jx+8jj45dvmTnkoYk99r+
HHR7tm/nvXqEY6oubzA94iMoU9wSE0Sfzrc4v0oyZd6tFoIokyzhAyTxTZudqmrQN0PjDEksYKPH
+t7nJwJfYokfUpP7cjrdWk2TYXcMJDpOZifxN2pRnHjqZA7N5jlUYvpdTeMVU1SK4kMy6vP+G0Yc
7Au0LCU4PGIon5T45rNHAYsxrqAObyOfb0qD+0QRGjP2Vys/FotnSGaed4GLVVnZrmV5U+iCyqpT
XguNjheqalAPdojYE+SBWiWKCQ8GSIYcwWlhoTIHkwnfO5gbyOZd8tkBSWyz8QBC9I879pFvx5V8
xaytu/dscssLwtRafo2BU5SyPq1R1NgGu3vrxrcFawVvMYhLrrLz0jYWd9wkvaH2r2Slaqhoh6zI
FXofSyNQqmbCMr194YTTnf3mgK4As72oLdbLGEF2H1SupXbwqiWs5ahFXl/rzFftxdiA0AQ4VI62
eyJ5ngwlip2XQs7B4anYj2t2r46icl/bk/yEXF8VyZmvR1xWIaLHILjtwOwa4/3AeI8e2eAsPCme
2BP9CsJGzN4OuVNT7zAj6a/rHtejzX1afExKbKSMz9D54ynygb81e+NYU4Nz6Xaa6RXL9HpewSMZ
rY2JbP5FTmQZyxm+B8UcoJbYrEgrXeh9Ask8R2HDi+a4T0h4tcYbZ+4kKCQVQp/rAHEMpDr+xPYf
/I5D38yJYylVj5+EPswxlCrQ9pVJnKnLAvZbtFERcAHFdVKNJCCoRCcbrAUczBhjWuF1QImC6D7X
FMeaQsrZPuyhqTV+3IWjicH5HcpGlKhDYfduDWkjpAtaebKSAIfQ35sficpkxJSgiC/a4raQBIa1
GNF920Tp22uptpgcsbmahHDLalw8tk6uSjLVn/ZJHoKcttLPb4n1B5lG1c5k1gqqo+98o6rvgeYX
SCmeZkxXtoXy18W6mresvRfg4HFpKmb8S9vC2/3//MqVbUZOAdSxYduc0NrsmbW8qvaFnVvYvsNG
/zui/EzwxoeUvabFkp9bMaw9v+A/gA03hNLlN/+k1DCZHN7GEcNzF9Kq809gLH8khfvwzdR3Q3nq
7fZToqg43DfwDx7zWNyfRqb8vSKofEEICOBK3kiLa3fW+xmcV8GZJf6y3ShZhlm/6LSBFlD24a/S
NIjUvZcihw8jPcY26k6s0rqcne9D1VwpEXvRjdBkHyzH9m+7RyEDcRmJsVZSHfsKnwjZf/+Xmzff
PbeOGSQiGVL2V7ETZB/bzf9wLWdDOkfIDgiXNfbJpAXuiCMzzKYvSkbyTZJld2G/eFA3M7z7FmR8
NLTjnWKsAOYdS4JbCDCv4xvBIA0ay95Rcno0ICkdTFvBn0h2Lu10BK3/P6dCyGg+vCW5n3+nVeAi
ImlSNiXdcj6DOsHjAL/dQTC1rObKmDIMUAboxT5NaTYsXHcQaEXyE66HOHMvSLVeKScILRbHVo1R
ptVfj0JRO/YLrPUavNTZrvFFIkH4jQRc4Rl2sdQKJ9v5mvWNIZVU0+y1Q7N2KdlQ7Et5AWdJJRcX
glcsNEfdgq8Ufh6tyEZ0aSzkq5C7XxBGKU56y8opgN/mC3hwK8Nn7v0tlmUWW+z+S57HhEUhsXrz
m+lPXj4xQSMpj/bLhPp8xPchVTNjcTC33Wxz1EmWwJwBgB0geXhicvIkBqDiP53r+CUeVebRRnoN
v0XUjSG1Q+BbxE3HaPGT/asTopfBqfZBWrVAHL+/7kCOQtbGKcU5bKRNkLU48MqhhoU1Drw7jhxA
crKbq8TQ9MBBX5tNW5BwC480RCe9PaeFDxFgzEZP8/pel8kTVZ6hdzyf36T8pLenKhNoQtikxn24
bBq67PcAanR/txQoAxinMDGwb3N2KOQaH9VnjqwtOSVTUkiPo9S2BJR4AjQjaw9DtOD5rsmxgYVM
SNkI86rOpfW+W8yle1ggORQK3EJifKZlIXqDL7AYPaadKiAA2lhSnJx8A7kB08CrY6ayomF52irP
5X1Nqo9BhbFyKHTJx8PsTyOjl1LBo0ai0t1visSpVddhN287eWCsWtbAOUsWsHvvCo+Su0fd4CR3
uN0uMKHUm/1L/MK7DgJOm9VmVUSMlrdd+op58ofz2IGa/ohZBGckntn/9xdILxjQyfpw5/5JiXdW
dWc1cfE09kUA1S353dcSUXxY/xuiWnkx9hFsj8pifULfVdrgIMVoQ5hdybDacshut8KsUAqmVk4S
C7hEwhA13pkTZ6tcTrBn0ZD9yIzTIhMf1TOheEnvtmAPmbqzP8uZczZ2OdbZtPB4Ya5J2x++Fkxi
OofAe0tl96WkUUmc6z4hguPcNJm2usIS/v2XgukKvcvPs5cpVV9Y+6KU7bpEfbq5UIGxtzukzV/r
DyHV5Dr13rmyEedYi9APhyGIvaUvZTKYX527eGCrA5rBXDvbZdF/3AZhA4//IcEzKSrfHwPLKpHU
TX/yHp2oYmlbwrNiaru1qzUnfl9s2H6qUANRwAANxQJsHOr7mCy5jMMVTr0AYUGB92uMO2p8jQTB
0skMu02tFAOOS4h4hEJpR60GH4c8XxPdTaaGEl+DyQVtJy75F32SQwW2oellWAxhYJdQ6crmz9Dl
v42bywTR0JpvtNNaszkp7ucIQSDFboHuCFIwuzMbCcz8fps0M/tuiX8FscNRX/PJqUg0fmGm8CpX
0BjtYdVetTe+AFcviGVFqHeG7dlck0bFCeliyO6dZN/PjhyHUEl1bL2JlhQxk/vgv6ttSkuszrhJ
Rn6p8ZQaypanFKRmWKRranqjYEQNYdc86ri/TYgCRR3MYDLO1RXdyWkaIyU8vDGjeeIS/Zyowoa5
vR5Wkf9YMa6CiWdUGQ4mjFkp2dxpPhKliJ+F4l6ZcrHE3UA9q4anzAGFoqTf3sSgWCj+OSuy9wCH
mlJm5UiBtF+g82+WIDJWFocWfHkb67/gs6WYd4X3QVYROHWJFCB+mxMT/t3gZ5OQwg0T0rJ+cHe1
U8G0QpdSJodz2ldFkipIvrM5VBv3PDTv3PpfKvk9UuQKKwbdt9S8evp7SgSDFC4+4CsYHryW8tLu
x/s3rsoRnvv7iZ2DVR/i05eKwGpzoLlbUZW9ryHCckcK6B0TB+5PUouGNA3xTuGsWBU9hJFhSLCa
CsoFy5jqNTuY/tijH4Z5mZ2haQjwfG443rUCcI/nZu1taKsJxcJyd+Ul4e3woicd52alU7rQTZ5j
Vjtp1bClkmznSx1FMXL9Q5FXogryNWgwMJIiQ5nOiq93nl4mo3V+GZLbzbCbvyADAdtDSzB8G55S
g7lHFAaXse2tV9HlP5cY+ii4QY5PWUWeKfZ1tbzE/1PlzAw/AQIS1loYvqcINzbAPoq906OLu1d1
dZgr/9kBIHwfjmvjF7J9ZmO0kWJXn+KjoA+X5b8e+XYO8uaWofcPjYxxsr9Kf9eFFLdvSjvRtAjI
lFFgWL0mC6jSUFPSeeM/1Vf44S/pMlgNf0H4F/I54H/LWYNXnoR9ofvNDW4xTOW4YmPPA5xzRzFR
beIiFWWAze82CNgEEUhywNQnYufjZA4nOCf5xTBh7fyzE5dBoMw2OlGUhZNmX7QURW+rb3V/lnmx
LITAMRsuwMpo1MNsFTJlCXV1FjurO5/YB0oF68vy5A8K2PhO8xee9vJm4PkXa5iWUQ+La129CiLj
cr+bTu8jmHOS4fUVoxw5V5WwVRlUblJOKik3k9TmnIj1Z1pwQFfDTkCFFV0h9O34vmZUm3pE7T20
g2PFwrzCvu2XbGjRJWgpQPu+QMfxT83NHkxPz9FhoOwUlgWM6Irv//NfMXzBN9k+p8Sgj0Zn6+Gm
Fm6hBW0/qqH6owpA9/lo+ISXUs66Pbu9bYg6cmbeAirOpNmXxZvxuT8GXyKmfdpbcZXDZL8igI2T
Ruf4XBShpE965AhzEEC3sYHhDj0DPXsUA1pRZW2pybglqbuDg0SyuZDZPY+Gcc2N2kFdYxI7lMiy
+DF6DvVhwT0uQl+Y1LDgIwmPKxs0LfNIb/TEWpHtKfdIRooxhmjySkZN4nrGkLxsYmLhV2WqMod0
gAx7vVtKKGSsZanhWAoE1RQSbSo+igHuQ9CWvlbg5IqTGaTp3HC9j688CDfLTMyTmGFQbMZo/Uf5
89xm+hjTqPfHK6XmInrG45D9EK4gCcdz0RUn+48u7cH7+Q+yYz1ZVXhJxSKiG8rngarn3uDcVf1C
Qg2V/+fsf3aEgdXJO7AEdCOJfDryXJyKFx72N/KI7TyIu3FxDr58PdHbXxxyfW1wbZfcUYh9fn2N
ZNeAzd79px8chxYQ6J3nw37OIdv8QOEX7s+CT6M+ZVJ5N9Hy9JnND8gID1yWofaP3rd3Hloumz5D
qRMnijLq6FY9FJUrECUJXQNvVAkVUWsc2pLl9pX8Rf1TxO2vg4F1ZGuXqtd/ySyOO1Xgwt+yAD3S
YI+HpBRpN8Q7UhrbhtsUwAXM2RYCsg0ZAHe/BBxuDd5vo5wazi9rtFVqevqHjtPHco2F7l9WhObm
7P5Uk4w6iOvPhUy9NJPo9x60/pa+OsEpg+aOpSmZYcLTbuBbigopdyNilw1erIZbQT0o2jB+UiIT
8+aRua51Mc2peBrTsaBdI5LTElOpEoM1qgcc935hJqbKTYS1QIowBmp65ItNPsVW6CNCwdaREHTA
eQI7j6bVmxhCvA6XLafPkBx5tEQAmZ+i2Ibn4VoGzxySqDjSVZLj0K3SPlNWh8HZHA3lKNhbMU6P
W0QviTOLaAUbApvfvnJyL5N0BbyCCoT469wmax5d9Kg7fYyM2LZY3pXVfCqwnvRz1Q67SFUaG+ah
gps2CGyqvQHTzh/KITM5j6zVVeOcvBmfhC6bLMjDJNf0F6fnpjkwskl4IX4R8/RLU0RmuvHreg8O
y8LU4J01GxfXF0NX8zbswpvC2dGhpf/BRl4++MPW8VtZ2xTfo77lwf3ntW3kB5YMNLCRF7sb4/a6
YJ8srS7KjmhfaXEOpxo0zEiiDHiRbaYk4iBURDUkT6MWp58SSYlysBjbnI1od/9Ayem8mhWeusih
o9EwICpB8pCcBYLK4L7xiP9RW8M2BIR2W4wjnwo+MMkEufb0bVU/B7HTb+7W/+vkDHHQ/WDZvo2I
pfg0b3ZY0LXa8APEe31bMCx45H+JeKvsrSXIihiPXXq/5dNKlh/nqmz2t+dbLrqvusmD7wup1ofy
gEZFeUsCZK5zK0nzOX9VFZUiuKOxMBsLY4XUEhYQE+EpEgYxTUaB01RGCb1J6g5NDS3uyVO0T7rJ
rO0w1Sq6yGUTsAyOZYFsW1VI8YXUk/B/RC6jRUVLwhtxz05tIMcQ7Z73R04J7O2etwMESR1awr0N
2KL5gWv4t2pzHpHYuBkIIEDvQEJSmrqVIbuBlm7a/WVDpW9FStuRRqQcSWjOvVJN+Gcq14k78oBl
0lhVNPZAvFfr1pWWxC7I6jYKVvEbHGAQw0Fd4B04iiDTt7ml4lCLhmKrcm7s25c+VJro3nyD85px
oquL1CcZ1dJnI0+Q22e1tM6WoYKPMdtUaC0fcR0bSHlmR4NLkdynUyFtoWbnhUW3BIytI53oVHw5
zOASUXUjKkyjYEGktZZj2MCt+itrxlA5tlKqqQuBEhUnVEVDJx/IHwAvKQkX7xsGA7g4rCAB/u7U
5aeYsHYv4wL0mrKKwqqG3ltjhPmdUFDo9ejCM4APlFRvPFZJ2nISfDVcy1Ho7TbY5HtJ8jUUlS3z
crGh4Qn7/imTVbnYyY1qM/MCRCqsB6WTaWfCa6UGuE6TBA0+Cfj+jA+mPEity/UNvpMd6DIZq66P
MmZHHpWGBzcgD/3RqCqY25JZdhS/CyLIvlUfto/So0mrthI5Yigavy3AsE8UFAodALqkHv5V0cER
YkS/YWhUtfe8nNIJ3L3Z56/aQoCJ/7Iza+2HJ3BhY0KTNMiTjH2UccfYD9lmD02YVWDYtW3sqwdZ
059IvGw0RxPmtEPjY0/mwgOwrLok5EdWEcHZOdu+JW99Udc7B31AvuS6IF9j0klzKKi3C4jI31d2
+n7GaarkEjc6ftIL2t5FpxpCEgVZg/5urHfE9CSCcI+/I5vbrNd69YUjX9sPhT5QhBx5g+S4Gycc
zEEugvwr4BEDs00N+H9ShgbVK/GRe4tzWz0ezlzkbGObXroV7Af0daZJMt0JeKMLRJo0YyZ6KkuQ
8d+YI8wSVu9TmN0MqqJjOYriyjgwJbubiwEJDrq/kTdmDNn06o55r3AzljOguOUqmsqDGizKQZUu
IhdEXv0HavTgiq7R7ffdsrowYITnSerpMONwm0U7oKCC7eD3UyeQOCeU201hoC+heO20GTZAIQVt
SmXAeppGZjnB85EZqqF1Y0IkOWQk8XLmcT6KwbGF2UlkZrJuOEZRzlmXuy86jLbBSSxkJgwkXDDg
quAwLo04kqFZr+93Nn3HljQ31YzaYZKKbTD8o82r63gDz071PJuNJSabxR1Q9qLIKjsjzmc763Fm
fS/7kKuhR0fa9kgxp5EsLdIaJ8Vm49B3C/Dr+89C6rHFq6vW5xrcsMMgBdo00j4lQ91t1ckugUWR
e7VNCKRXcqSETdHTAOLq2w/iq4iyYuHEyUJ0+JKEsC0lTR+6leAebnEvPUquf4mFEG5Hdvfrd5RK
Nd4i5AxfIqXEdGxQH0yZ2RuGMvTyWbISJ0J4EAG9+sGVhUqhRqA08wesQMZrLFv+3HrrhJIUFuPX
UurjqBYupu+0pF2orWtZf9ntXsIQrbanTDi+0jVDi1gPEZYDGP5xP+XNcyZ21mGXRCwRkJUB2lfQ
B7m45xLJRp+uv6T+IDExmlJ8WOL8BWSbtZLakac7QxvsHcYC/SSx+G0MrmITqPgwbY7QYA66dKy0
Z6bZFQ2op8Mbel9tob4k9EQWaytSMUf90SgDGz2lWpdmGcwHbPKpKw3reU/By9+v51F0I5V3ER8t
H46/rUfDL69pks9mAxHaJbQ+bbKiRXweqTP6VALKpSMWmHiM18yGDvkKBdilY4efc5wEgQy/V0fC
wucZ6iljPwCllSmYUcszJO8NH6iCjEM9cqVPUBG6vRYwKwkvSs7WUjpXz8JKQliEL7aFQXgerfQ4
JvpzgeTDn7/53VH+1SeAyag9rgjpNdhMapLjBaFlUBbVXf20GcWNfcNkR883llhFHKB4YD6rD3Kc
3tSxpDOwkSzS+RKgbMQvnk0xe7e/eW/9I3lhicYPJQSToTsWOyrTpyGGDcWrtqxxRNtt8eWxq79j
DygLGAME+a2fqQO2Eb6OQ+MyeWzpaC+74qx3SEj2XVsyPw3OEQ2dq133LhNlu90mAcq15pEXqYT+
yGGOGF1f6mCOINoL6Rvli1f4NkiOwpY05DtQiykNfHrJolUtwiOmibo5OEeKI26fw53KnpB1goQU
kq3ZNOTjYKdTqWFE9dqwCMG4UxznRrSqjD1VIxfUxSKg5rWUpop8p5DdV9nhGFsiipw+GLPShQFR
OGEM/OtjCFoLDUmMZgUtebp5YMgyxP9H0Uu1vjGwZXZcZTBk7BVDuFmiQYLwxF9LqsSBJh/0mMJM
OUMLtnNDES26MMQLFa7qrOYJkdPale8YrBP9NAjxDuZbUklkY9Z18jfgB6aHIJtpSIXFMrOZNYpp
HgqXg2jwFvOG9K+Aje7cFVSRNj1sPx7u4eNOMsuLry6mLzhGkcavGShbK1RWB3cSKpVUTFtT1TxW
G0uopC8eqRam4XwpkD1wlinIRlDkxbMpzcH1EB9O4DsogBLq+jG4Pgku8jeuV7mKYTIH5lll7tWv
/jhhlWIMU54eV4YoatsRkHe2SMSNVsn3+G8PvZDwovjAvi7FPGTeI+WDJ8wmH9hJWzmJvglyC7PW
SLYhLqYwYqUDL+o1MNIRVRR8JQ9j4mkHbAhf2twTMoZzcooM2K9pmEmuzV1OPeS3cRE0zfq6rbg7
K5c09smGHOeh+aXYhTsYANdYw6Jh0NfB2smD6/SMKqNmhwy96Mkv3jtgzhWiWukyqX/t8nYSve2H
d7tRv2PYiulAEHpZIxwMsLpRJMgegBb/YwQ9gfzOBYQ1ttFmBer8FjX4T3IglGRG+Z7vHhJmUqTr
vNZibx47Jmrnr130YhLmFM/oxGvDF4XXZnxqpt5kV7ruVrSU6pim89ybwulWMresY8Wez+B5FLwZ
TRmb9F0pLYEUdatO6M17ongLnAn+50ySesiVYyPOJ6WIB1JcN33LuB69o37EMG69RAbOph6jCld9
/bQTaLdTtfODIENX9wI9zTihzuQH/Gz07FSvwgiksUz2flSMftwSoP3zBCTxNJCuCDihlMIPxxk7
K2wr5JTVBA6Bq9xUL99bBUtXaxIPU7DsKZA2B5lTv1T+RQx6v0B8J3GWicVDfkICvqS9491qLyQK
kzBWEBQC6UXnmofcCYlPRZX2dCKj5vk8H7XHObXUVddB2UnDwLXoPUcjdX8T4jqo3vw/9PsWWmfE
ANBFVNPCVDa9q67yl1Cfw+4L/1863nvNexTpCXjKBDZO+bcIN8l2hl3bOWW5U9SOpPIPGC2cqkzB
xiFQfhu47SlV+l/ilPHSaR5MWq8XjjekxHYexntD74w6A9GZ0xHbM8AxfSx5pmCFgUY44WJWP7bP
Nyr+uUBXeuswfiQhXczy8HfZk4zSC9DY8Y8rxWjttJpz/zl5y69MNidXDO2pdxy5BYAQOL9dvnj1
+3Itpamn9R5A20iPW62QYjpfY74htLVK6Wr4056c+fg1f32IpxE76nOc7b0mCNXeUUXtJYtpF4py
az5UooRdwItT9TWp5ExIlGzGWjepIPYJpQZIYEOVpcefuzmaS4CIgpkTTNhCQO3EerLkNZm/iluM
22EAbDT/hdCFJg36Z4NUxLbFChCm5NOmV7BQodD+ujSLfZRe3OKQuls+Cv+Rkoxr5rZ4hGxbtGgR
M94xvp5hP7oOVLxOjuEbizBI+3pbdhc7PXlpA0kcOTaUkSG9FqYVri9duphHO2XJWSRk7AaLcHb3
VsJYa99uI1YcUTa/zTv5HtUfNwPitviMzVBGbGYWrYdozQmZr+EvmNCpnwihZyLFIvYb+GH08wvP
LX89EqhzqtwIgxQcCIHXwsP9keaMztQWRRfSKu0Zdx1t/Lr610XSaUWks7pTigCIcr5FFPsB+Q5e
tZtUm/4Y6UwEF50zqVxvKFYwtJ1hdX9Ccj8IamByPRMDtCRxQT3v3VcRMo/VMM6zEoHfR1CQVQ/m
ujmGrQb228A4rnQfys5MD2zAOBpOv5LJ7lWlfLaeul7iizjrClfKiZ1f0zIqfDtKnbxLhXrZPJy/
9vl5no6/2O8I3ko5c0P49+HDfhEoLL6no1IBzPamBzyUBaaWLszmyieynGtdwXDR23XZhfidxYt+
awOrifGhPLaTz32fx2aZ23EBcfUGOd80FAnj26ZVbojvNhTBVo0fgmlVBhxxoXo1zLPRBuAG3Gdd
MjYJ5hzzjbkQy+ukeWqFow2oqbeZodm7i4pu15/CkX4lqlEwBawTpWFL9nRx2tLuhNmgwBA5qiVm
iQ7CnDZBVSirHhY5vbWEgmvOv8a60vCV5uY9EoeDAmJqZlYYaCSNy73+brA3P0aVywM1CYLk0nAS
KOwARizobFm+jq2i/FQktB4PRR8L4DlH86iioe8ktt323146H61nWDblUlmYvG3UMIIM3CFOyjMg
bgUTNFsPAEDMHkp9eWYFmMyxXglEefBXO5RfTwzJHqmudr90SPq9PM1QTWH/Owu/uG5QGJu3W9Uy
6H+ZVAOp8z9tbGrPvjl89Ql+mxwRIUIj7e/pDVDMrS06NKo5KeMsVFfL0/QGM5uL02fO0EQOLOkC
6cTv2G829ItCFt/CFwlBk0vapZCo3DqEalX2zAjsjg5zYWJMf1hPkkxSRlrh+LQwn2V1g6FvBPvQ
PsGLh6emGOw4dtk1PDzpD8VX9/lNh4vcsK+c6wTeqyBzk7Xib//t1hBBVPbiq6v2LfTb+rN7nReX
UdW84sxDHtz6ebw88yep0dBIxz7uV2yTLeps6Hi0Z/q5e6EKpth1PwdbtdGmccrCgTU8kAaILune
Mmpz3fH/STCGJbvlEY/TuEq94f8lQLJaudvVsyHHLNo/0TFpbegm9S1Pu6RFYpGw/6pM4o9S9XDl
aRKwDS09jA76sgoJHVM3TwNmiMq3c9pnd4MKHuz4R6pX5GV+gQ1WkVrgCkbTUf9D27HFc35me8du
BKj1zmxApFxKxb8DXCwKKWmWmQUOXb0Yn8gVpe0t9BuHrO02euOgLRyl2Lrx1qxhA1mWM83TMk9E
tren3XOzNAc5FOxiVDU6iSgkOAwfYdZ9N/mppEXbgNKfrCL71SXW5D++C9myLUzueGwSnSLXzio3
Qca/bNBEh4Zr0iLNHaexAzNEonAbk1VSdi8EeEcqjbooR4Ab8osfNxmCBT9Wa6j0xz+N4p7GMLTC
ulB6oAKIP0+hb6uYZD1/sGUr+awDi/IRJ5teBYc43kTKj5ojk7AyGpvN1AlwNWwFmjjfG76e46Bg
Te/o6N56Lw7XZGuBC6/CKNXThUTK4nb7fJPWOdlcjKGUgRV5NIcTyS87/05zWccvvue4cXF1IlJ0
tUUVTKZFZnBQMuhDEw2DXLf/AchdQLnL+LumTxsG4EsE37YfBcdSml8QNtVii0qgA3Da1F8Nbxuc
o4H9aJdUzCkp71EqFjE9QCj/17RlcqD3LI1j7SrkqblVfZ//B93vYN9DB3ofpmKa9S1M6bsopzVe
u42YeAeGPwA9ER81P4DhqXoAkivTb7lHMRlSdZ3PMdpOqKDhnlwWm7tIUgdpiGvZ0HO+rA1AAPl7
Ng0yTa1WEt++yu9TuOQ2CErmLBKCruJ960I6Cv9SqhJ5nc2FmGzRKmq66d+fkgIPyiYEnrZp60ki
RRYimALMwNSO0bg64lsq8nNovLEfUpDbM99IVYlxy74VnIqXvnF3Zf8MPoV3wlYcvyQDKc5CWWY1
RhUdlzXBlUd1qkqIu98UUB0ZKBzy70c/Xa5Eu/Tfqy+SdEB+yZMmBJqHZ4EPCp5SLTrOljtoZOzq
Qk43rWbWWOmsFSeC7fiEx/F2A6MxyWCDXBtp5+dBsxI6kuw7/1W8YPzkG4fpvBQeWUf4oEvXAQTi
np26LNZ2nYpnS7VzOhp9/rlmKjio6uWwItYyByPukTDSgu9ju+17LFUY4jpzhj/usCJKnY8tKW9c
kEnWal99zWrW3A8wH7k0AwAwUdGVINs68LxYLH1uOXyAWFQPthK5LkmAHGFshFZ2cZziHBCik8Ga
UpMlVK719oRFkaXVMYcHsssxZbPeM4jArEc6T5MRPWaHSVjXpduhzLNvb5P+HBSSLNA2EwXj/WDe
X3+z80BWwwCFpEBRQyG9Dc4VJQI7UNgCIStCy+rzElzfbMFvN8xIUZUF8HOJRK59l/d8Neg5n9Y4
ATUoeRKXX/vdbbQ2u9tsMHKUKae1LGkt0qeMFQfxzGWSrItNezoPypGGQv/dVKTJ4cm5eElmRS/8
Q4oZzEFeBhUlCb+sb67oLOWNpYjocqJlVBnb1wYMdaW9g1u6FnhiomyXizNDN8Q15K+K2ww2OdFg
6JYQCWeDh6n0Q3HAIXb+2WzAB+/i160tBHfE1FyAefHyZudgE6mdjeQ3bOtaULDx4hFpCWrcjmkl
jLG5B4HbJdpn9r9zmyEI07QHreOUQbUbIO0XpiE7gqs0FNx8c5AbYIgj1Dn8UWFjKd+XcqRddYZD
XYrq7wzVTEeToqJwl62mb/vAIMUXhHUWbYhUBRS85aROJu2+MvE6mP2CdRt/3B05C/NLfwu3mXDl
IcQzwBhPfWfaigOngpnjBUSfM9IhcZiTxb+Jrvc5luhoz1yfgZot74Sns5BcWP1Qq2wXIHjxE7Ag
RHdDci4ojD/hVCmtVWaApWhcfmSxEcj8sPO99dGFhG9CDD5jM3JUKmpVlD5M4iCDLKtzcpW8w48e
BF+8dPTFkLpKN0jsSA07pMFQXBcAjQqUSJmcTVAbRW/EL5XfG/ZiLBiRYNBK2CedSxzSqhiyXk39
b4BsLruFhKM66mrFLzyz04ZFPEMmO5FerU6ZrlG9qJSxxMuc6KTwiGHBcxWWTjiwmnE7E94WlnBq
a3LH6+BA86lIRD08sXLJUvXe/efeQ51fKV+uwFftZTdhYJmdsXH2WjZPkh0pz9HgkeZ23BuRq8mF
LEPWyNofnenqtV5v13AKfg9TDoRhtHt2dBQ9ubU4JwRBAkmfhovuTBn4VknIfglGXc5JDkxheeaf
06A55jxItwS8VdFSFt0fVYDXzyZvkY9YwwrGVQVYE1C8wPBgLsfkkXeujrmBjvMWWd7GtGkpmISW
9cJ/1beTL6VqaNf39hXCo9QZcQYUAm9b2JKVLero79wicdBct5TXn4vl47XNQFMHQheKYHym4o6G
HRVQNGGqV5MRjbLCXPTjY8q+8zmeEHS5Of7/CS7bA+LJwVzkRniWoV3Sk51AhVdEmqcXHDbanv9W
H8QzJDsD2S6weGXhPYNfBRtpLKOjAAd2yoMYNOGwYQpqnFcaQvJm6pke4gCz15FMTiqrfjRRwRYy
g9+1bkNxfmwpP2gjOkvf5I9wAHYhtezX28VzEmF+FEz6n6H3BRx62YKtGIyuj/vvrInzmOiOxgEx
OIZ653SXl6E0V72JjayWlPoAR8JBzeHxcwh73yxOPCFWuT5F81AtPcIB364yQMbKueo4xGHhvgi4
EEJo1QyeAqFgG/6duiTzK+7EUI4DPYE17prKcbHyOWbN8kkkOD52YRvbqtkJ216d7U13T74php3n
vqAcbMiUc9j6jbG7hmjlVrHZVX3SA/Fn2/E9tJ8uVlMj2L2RvISBm1iqYu/HcCKaZbvA4iZor0Wq
ft6tYiGc1Bi7mD855xGGmdCC/OXvgEFz/soTAWOIBSPwPjEo+a4YvLP5Er93f+A+aOhSOQBeo1IP
bIiHERGlJcmLslo26pI9mMz4kNQ/hevpk8uMtJOVEnDo6VQJQz7pXqYbUjDmpThIiXrPqZaKs59o
N5H8i5URJd0s4QDboBppuN2oVSj3kZkTbE9AfXJ6ihTKKf4N4Tq85ncfBCzG4SgZbq5adhB2yBhe
pBfCIIKl3LqSv7Ocl59mz1YUGg1I8pBsMrjuNDX5/FhHpXT6LuQ3lkf99yJZINNeVgrZam+/EDWV
LOlDfIFIrXvDQUZ0kAlobXsWh3yWzEERmtvRcMrqodPHb2FiatceMdV1ELrKJnc8T5Zbnw+i3dt3
g4ak6KDzYH8NMNwUShs3fjrjVO1h4guXMvzSC7onHARLKU4e4a0bfRyJ63wENlBB68C7JUzKwHgH
+O9nDH1kIWgjACXwJtFbZRDTC2IdYmRZWa6WfSk+4daUdeQO19SO6R+2o7bnbFHB33e6k/x/rBpV
hOyL8DBUUjTsE1DzcjZcxsN0ZKibQwu4G4w0X6fUi52oHpsJUTccydwBl7zxNpOy/XLVhLjiVRli
kZJ7lIXGgapOeeyV9IUyzfEfkKvFrzYPkC2x8j7K73+5QxsqZFx+p4BKqDnKc+Mas3SKwitvLqNh
l2Hg5ysBZGtFyuPtTGnUJIMNUsb8LDwN2C/HiSzDOnt9wkT/zPyirxFgfoyA9OqmsraFPF0gbVQV
ytzVIT000BVwR3HP5jj1VmWaGDw/ver31NeojVR54eXPboyP6PbsvjWhsdzYtJzlmmf7/E/Qr9jq
XaSm4cevr+Ogs+rXUa8Yho+De/MDS3GJmGsyvDIrt3qOBHypW7MVYzagQ80QGfjbiCOlIVUP0gz3
CC4EySnnhEOxC9xW4fNk1CEkidvez7RYCP8UeWUCE18kK+t2QwZAUcr7IkYa7TyOwGtfl823LRXd
e3YkinA7+36RZ0wQiRGp3HmqQtBT7NfpI8y5Hmo8jq2kFms1Pul1ddpPAkyFM2O2IyiYKjXt6d9d
MIenpl67hlOCznkwgFm4ltTvn6i8vHDJn2sYDMb2Z6PXxcpM61jvTqh5w+rTOhilVa8u1yIsk0u0
knTt5nZY+MTCLdynafHPgsTfZ2w16waPbyDUSRNlP+DHbqXxfdmReSFK2k7oe9ShYc8GC2+cyJVE
BCaXt2gcgwZjxs2kwqb3TFfrhk0OjOOqxUd3umeYC13dTuzUw8a3utVyBANoP9vwn4+aPy5UZ7zU
ujIMaEESAYUVu06NVPmTLU+8eOM3lFKVQMZQcBlH2cB0SarGRap/ekj1P3S7KNRqWHGUfwjj0oTw
PL2rIt5U+Gn15Q0JSoY8fojfLmsWr87wh6XAgx9GicmiYzU1isbEpdOcw8R6s9jm1XLQFaQz0p6b
NFogT8kgBkFdVDmrje0As6Q9HsTtamfrJowoMyhaaNM4m//n2KtoJx04Va3A6hWuqpyZuXz3gn05
nb+OTj2FfmQpFAB/FCVMN6SD9lD6Q84F6T53nBWmE2CJ8QcM9Wf9LQB45XcadDMl4CYpnogX3LaK
2NZrGrhJUqwftuKdPUBolO/zm7+Vh7K49PAazx7WllBfgt0LZkyfPe19AIDiRoNmtVjyU67R1wmH
jObmxAecnJXxMoUzXD3K65yS1/XdfhaF5HkZae52pFC3IpKoXJKXk9N1WteFCLZrLtkBO6UA41EV
PvqP9KBYWRamqmqzrHcZ5csycNmhfUOcPCRqXGAWMyPlbMHn4LdmXX4yzKIB4ewfb2k8Qi4A9f/G
Svz7CCXyncuDnULvnag3qNv/bhcik1n76RcCWioYjywW6b0An3riXLX3ZSh4fTrs6Fe5dsaSKXsM
Ou47Z44upobpqWXIGPzGI8zvGfOeZYIR2PBMX5QD6VHTVv3ugz5ggyHwC2s6KOmO+917qIaMLnLy
KpWKpaPXIcTw/iASAoWu4HWwRKQl3TSxWIqMr0vA/COmRV/WwNSuVp0oBppDEp7kbjTOzWna163X
vhKy9Zgb1NC37jXcwZzxwx4wbZ5uKYT5TTqjp4CGmnm74QfyCG54fMBA9iKNdj4JFl2Z1WP8zHwH
WkzJYArUP+I19bpualTg6dBd77jGCCkTtmh/OkUz/7ileCpYFCKD01hGJU2OvnIBwei3llNWo4Ae
VtWqULe932Geb+pw3gk/KmqKOMfDUzsXPIW6U73HJtgf8/Zo4rqJTXPgu8ZuT9t2UPReES9Mt8Su
CdCnDKsaqXs3Q+XZqsbxZjO3x/QMLdfuQo50+jbG6aMHlUSHWwVT/ImKG25SvmpgoIJ/4j+p6QUD
hgJpzuzXeZySpO3ebEeDAGGV6EuR6PwVR1SrWcZiQx1TjA3q58yV2HgJAJuSN5Co1VYH0//0ea+4
6YgsYBZyf71uLNcqkkqtjSMiJW0UqcJg9iekybAXTES4Ae5MpGrbQwHve8Q1SZoJPK4WuH2K5dlx
ebbfL2k+WG/J5MKwh5oQLGMXGMJd8vWI/VvMd20jLTqkbwc29LWpIREoMd/ah6ohOlKHb0qlHUwe
pzUEYqiXSvR2ZenQuyyuV2LR/FOLSzb5d6NBLBMyQOTiYA8H4rqz99ImH/qS4vltAz4tMATgWGxo
nA/OCpNeyVaCa+tSmev9rT8npQcxrbcpnFZsqBWgKWwhVxG4gnLMVIyPDZTK19BwjusHQh6GY1Kv
xhQLLdb2IHyFfa2Ov6obub8yAlWcJKh4IbkTRP71MsqYKjPmuVW4K3fvBxomjH4PgDrkyWAdvA0d
CJbckC0tCunzQIL2p8JACa6xhP833+9gwndOh400s5KyXcETmTgcskXkIM/MR0H167ImcgIzqxgi
1qDHSVITleoOg0f8aQpY5WhxxtflCJMPPuBgTV6+FQcyHTqIK278Gwj+z5XwCRGb5llwtkRV0LP9
ikTW30JwreX+nNJhqUuVLR+oXg8Z5fnu2BASKht/mrECEI6SwBq4YmlRXbJZROGQapBzlVz+8ZXM
9QrZ3d2CNvIRdz9C0SYYMVGDDSDygXXf78psWycbZuAYxDshKpwqdCFcTrdupXEhRSDNN19WTmRB
o0H/dH+lvwN/vS/qkWKVEfm0cSoLOkD6PO5pYbtpKrYwvDYDaG7MMOS/5agtJoUM7/wXApP2LyzC
DyJbVQn0KPhdWLMi6Rz0FEf0UKUd+0aRiSnsnFmr+RquVbZIVOv63r1y2mr1CLQ2e/+sq29+YSoU
0q15Y1O52BOsKqEQoPR0dxm4vfNQeakw2XzUvUCr9WlJ2JKEEI7RIsQ0rSMl1MeTHmpn2I4i2yB/
uBkcV6f7dapDPSWUcuSZd2Mf+sPNr6QL8euDrtEZ6TvDjBHfkIHcK8VAxPy03vz87l9FXUQv8ITt
OKmLtAD6L1yVwQkInMILmP+ipYg0xTI3l4OEBfdwPZmPE2PhQRPKV7Idt5d6BhUIc+zO9/O2nndf
xz5m6fryFbCMgVF4dFZdzcbNvDLXKyN9TTcofGUCFrvGVLAdoF80YK9+1zWLhbEe+0KtLv4dSP0q
MoPMzmcGUdFMoirHqxS0H+/TVRQV/NzGBlZALW+qlVzSxW2zsbiEDawj+tf4p4t/SSbAAJhAQQwN
uPkrBllykMM6550wXgzSG1ckWCBpoMdmcWO/kwVGdJ2epO1m0H9Q23im02VEhJ/7Sh3w3gd++4aJ
sCdwMunUcmHytPv5yF5RDsIEcO432N1pOt/GXj9UmAglLdnTgmssg6oA/HnSOj+468efccEjmiUP
kxE6tNNczkCOS2EdYYHX7dpDBQ6imkLSTjjbgZWUmcrvUCOv2yTBSIstL+Mt0rhNyecgnv9tQZwH
/0BGGVZDyIWC4dbhJ83cFk3Y985ByGNKW8ax+XVGEgu16QLFdJ+zks4ycOd+pJqvj21b43qCJNlG
yu8E2/446K3uYOWPvTSkXYeyKUlGwa7zvB9BIM9yvkaiIfXWRcczNZLcXRGZhAfAEixp9s6Nrp2v
6szE71n26MGXAIHelM10LMqHab9c7eMP1aJ/8QL7KDy30UPZF9AVbrY1xrsfVkIfQtoEv+Vbo1UW
U3E3QRjs/5dW+YJHvY4BEpdUWIIAvRQpc6A27PTbjqdUZCPO46kGdKTpa7EM6uSiw6lT2UbpnzC5
NJmKX/jhF5G754nl6Tcky59+RDaaEOulecsMR7lpegETbHV8lGHuk4s6xTPE5EL8z6OByBPAmFcM
yQIhF9eklAfmSIsWGHUfhFLL8uacjdS1mpP6aezVrY3eVcVkN4IN/6ys9omyCNZSjVNLAiPZVBi+
exu2zK7I0rIuwmCiUOzDSYmJTdPI9HaTw0LxcNrJs+Fb32MTWtPs1c8pFMZBCRYnkguJQhgZVmeL
aVzjjIKMgwgU611087rNBy6W9RdL0dn55gIOiQ0iTUHSyLWytF+FV1aSlRM3HPjKrcFoeNjNyTmo
dJ7jt58cSL4smsomIKQVVEeB/j+6wtzZv1fhywx6HBKYJLCjm4PHwcZeWSMEXjcPBOiLhwXnHuMb
8fQdSdUEIddElyhdvYFN9wloZp7kmJv8Bf4HAnWOmI7NfCT12zvSjPfCH9y0ZA/dFBk9lxNI9aNo
y1DwdUJ9dIczu0RvfekZBFsVKmZVvIxxx84Qg31HROHeFajG7AuM13/HxrB0fAPsQRH5xHbEEJPB
G+6beWtTFHsQrW1qetTxvL8XP2GcMR7P7wWplHgH9ydNN1IzMgStNyTqCOIagc1Sh2PMK3iZt6V2
M4HxhQyBqBtJIpz5c2gBpdlS3EmgGgku6x2svtVvLJ9zpXjEiYPkW8ms49fhb+5g+78puGiWkA8g
6LjQo8Vy1DK4tEONLLz/nNjEP5K0coM5iWg5eRuhbXd3FlmewXOXUbAalld4W4UigUlrl5XytN08
9fH0JoBcg0pxyuUhj7iXc4UtAE2rJdIsnweGRSJtjT5DjE8e+GBSuTV8IIVUqjvgLytb+v4h2yc4
s1E9wH1lJqKOeteB3SZBOFj1TJ8ww6VFCJ028f2Xij2jL/FEOdHcfeyUUfkYOq3YUGTyJBk4s2LR
4+ZOG+J8V1fLNBiJmAbKu/0EF10BJX8U8YIZtmjRqEt47fKt357UMr6UI97j6cQinaOAeJKvAx/j
xJPG0krne3rCY7C+I462wvg/6H46ojbnFElHSQ+keTsxeDZvlEIiQ6E64PiRjPRrj2iXhIydAsAs
x7Y4RQyJaQ3it9HfKm1TWN78php4wsxNf7skpNn7KYrTJXMh0WEBqCdPtqRswxDrrbDrbiKHd6aZ
Gwcrip3+Zn5BzBoSgxF6f6NhoX6F4F77Drj3BjoEKX19/AxaXFkvisWAWR+esQtn5YrZ1fs31CuZ
UIgpxqDGnRMQEyZh1kewhac+QDzi6bo7Hko455eulnkf02EO7RdXK/4CzUmgIzMrqJRKkNjI/hDj
pKeJvFwjxVIx2OpUZ91j2mHVLwNZGMrLWz/wwsGe4G9xg7QmGuJYGc5KarEE88JvrxbSRHmobyW/
f8qR55WLKIrxkwk44se1b46TomY//3VhQ1dcX8ymNAN33ZkNGtfLrIDDBC4MjilK5cvhmwesXUvB
TYHMa4QYmyI3fGtJ1PsIqjAlaEMMTaJq0PbwsNlbRorU8j9D66mMXtiZBbWWr27tIyi8gU8t31J6
H+6txoyejezjWKaCE+5FfyohS4tekRSGcZPQcxN7qNK9e/0szRC1yVZF+oqFbPWyiYmoCzC3aps1
cdk2micHK2rH9tnEhkI1Q2ar+UzeVXqYagUSbusTo1OBU2yYs1YHPheDDE0VklOtwJTwMhCKA4JS
/J6+n5qRhcBc1UeGPCwo3vbqylECfANV+tC0sfbk3Mj23zPMMwuinS3ixZpUgz4YlTLIVeZBtuP+
hOsXWlHlkZfQL8dXAnl4eX9wsAqxSePL8wnwvuM4N3umotvmK8iKzeW0W7zkRyDwIjnnkTBp/aPV
yXbn1Oj4jr0h1Jm7jDJAq+YB10JOpeyCWRoCNZoNw5eIcJZO5fTUG8vvm3XG7W/UsGXTQDu6IjW4
FugEqkQI9tLsxI+5eHleL75eeXSVDH871ukU054dvB2qZlRXVhFjVN+f68swG/HvbSp7lqL3iGbi
NmuvNv88ZJP++y+076GeUI8zuZ5ZZRwW64Lnq2i9+6/hxp4536ZlQtVpQwlKaZHz/WCzl4YjG6WM
uI2IPkrlZZX7g+1SaoF9bliHneSCPFQEgSAp5ovHtj+xWZQYc0w2Pe5WgAmDIiAPKYT6eGWYfenc
Welgi7tJdjZZs4CoJqbH+HJR00m0J8xtGjMOR6l6gmiF854oCHXwZbHkusreW7VOHN5PbDrmUb2u
3++A3VSwNjwaHG8HYFYq65HYhd9E+BTfgeOTGMzE2IPBfa445KLdw/OwNhQqxT75H+US4kL1XBl4
Qix3vD7TwviImgzPGoWtBL35P+pdaykXHyvbb+eFShSoyT7IEgEaKvjfBHBjiKHOBVjKhbnrDWpT
EVIXRdFGncXH361pkuor77BcQEXXWFwGz67lKE5sk+fOr3d6Sf2y33CAe8Jt4F2x1uMkUK8u7MQE
yaWyhdwb9hPlOoPTpfScEJSKnADHn2C96ZQes50O9Qy8vaCqMp18Q8y5L88NbClNHNnkN9fMfQPI
3oIaRg8SKXdZDjtmSvQ5HsInpMUYR75uHCzxbqxXPrkapUXb0SM/KI8OctJqZT881xb1fPYIsSly
DdyluGKwPYxuhH760AqFFJXJrBpKowH+u1pJjc/39QEyToxL9/PXH9GG18cOrUlbCkF7CcYHww6E
GWl7xTbj8KjMvEwFRDsLTqsQxweS5/QGgJhUACBb6FCdsqvQIsTztDrd1HqMQtfKEqw+zk0nzSmH
+eKndsbqi+Rja0ZxH2DBAH/nefrODhkYraD2Zt0D0wWs3rhSfuXOJD0D/1id+zrtM33wZcQlj+TW
rXPLL0TwV00lDYx2k1APOd9otJ4hAvbgkfCHfmg01MHQ0cAxvTjqu6MdspB892kHtzfqQIZkUAO3
kTV6OglcQcXGAkNDqYbdd4Pap4lQFGRrFiAL2ssgY4A0rRFk0pZahE/FRvynVaVWkhPjoFMA7BlL
vB0ShPb7Umyu2Vzt68OWgnew6zSeCia04RVst9oMJsv7d0QtNKy62VTJxHdhk7DQC7VqYNB7QMtI
dRCDVRifRQnfWDz9Yza07sovPPD0C36j/geahIR8S7Znq9IDIKFvKcbpH74zNZlqWuysUHVegzYA
j+djaZvfs7QTRdwcpK6wQ3Olv24iM3havoR9xBQs1dRlhojnTa8cOH8RbjCe6zl+LbzDq1ClwaMl
rg/NboW4PP3KzDMKU+Vj2SirbRfcjGqfejuft5sE07IJdkuh2qM1y4U4SaBkG0JoRIOoEm/z36H6
9hs8gOY9CRUYkTb13bf82+3/b257Nc3KMi/GKIA76oGtUjrB39v0NlDzEOttak1XMWntmHr57WAA
M2CFwkXDX6hvPley44y0IL+H9rV97U6LaVVaqdomkPOyqLxByMAdbQUieUe0Lb61g0AOGMBhDGGy
crDXi6kbINbVVbHXGypWBbGTBA+5qpzep0hGRhQMeNldIbAlVT8BXLeVXtMvXv9V8ssBxIKvSG6r
SwKdQm0YrHPQkd7Ew+7rGnVRV3S2p+Ia1PWJNKSG+1BbFjUjkjzfrtJXF0epBDzlPaRclrP9MB4Q
nlkyHBklyV1vNkYzxPCkvruk2p0ZAw/sPBHT0kbwsaGtdl7UXDn4QOkiNF00DVLkrOD9l5x1+iNa
dB1T4+9uSP1c/cr4ngKnLsyDRsRjc/OMfHXyhDNKYnRkOTQm4mGdmmMXhXotK5/XBo0Zik4StmvK
r7s1sfXnHTtHHAn779hktOb1pVPSqBIXv489/P/cI9uxWEtMD+N9yCJsCcafxsD/gs8Ths1oLT6U
gbZ5Dt/hCCbkGQXCCkrNJEEd5LLAlPRX95uLXPrxj/veJoLGlOZvzPES6Om9YuRhCoF+hFmWxg8t
pazITGzNC2ftMceFMMHsNqFN0nuKvAto0LOR8ItPnn0bD+VfQnXPQmqHE5j+oZX8oV5VhTVD2frl
HjylwyzObAzU2axu/G9ft5Af50hB1+cAnyPzssmIvt0zTPn5zlLcLs+g3KaZEaRO/jxIfy7Hsms0
ykIIu4uUEbqS4ZlxVx5KPbDJ7+ibyJzEgDJk2/ywyRHolyNgs+1fxqA46CbkRqfSO3czIRuiIP4Q
IkS1kne79VH4KHD/x6pPValrO2kGKRhYyjatQhkffHN3zAixc26ceq5zIZ+me1Af2hm9cyPZhgDx
d5yG9Fy15FMNTPSNrz+3WCPFjf5RO20xHbDxQtoTTMhtxWRxGg+/IRVwkM2sHmaWb9+proN9Cike
OQO98TryOWWTLW/pql0qpUPZAQ1kFfhQbvXWpTU2s2XaWEroqFxx0sMbQAPU3BGc+kI2apPcAgHh
f8qNXD78vfd7VOnd6UhHrBxK8PcMmG3fOEclVD93sMG3O8C8MmQ3p6io2zGSbhAa8ShAirrvJi1C
EMQma2Vl0yiNEMDOoXDPypt9QioAEuCIqnZVx22OTLbv+qvQutLSZfMmB1yxnqgUOV5j6TvWAvS1
umS/V9NblJhgnQmj6jfCQOw2ojC5xUdy2FurrN8FQq9lFwef7fze5ZzHLPW0aaK0iVuz/qgxeKb5
2URmNRxVXV9uKAdRtjky9vON2KNZU/P0jRCHsPdx3dGryDJjv3lIjmaN0BpeOB9vrwYc3pSjH4MM
PK90/7MB9/4ePTusillgjFW29co5hAvwBgq2Jxh/cS7Z3XyT8u0gG1eaoPBDq8uityncCyAVUj/h
Bu3VtKwrcLF5NPiSmjh/B4Urc9shpt+y5H/CG3/jrLqgK9nZ1kUw7fvozzw3kE2Dt9AhZUyIf6Pu
abP6aBRqydI9pMLTdmY3gAeecfLL3ID6YGiPa0nKvnZZgRv0UOr3urTKueDS7Sc1KPNB+Ejkzb42
UpXTolY2mK0lCxSRX5DYpgDuHMWPt1KKpEaNCzkLwMJRvmtbWZUqNEu2T/OLnNlxnn5Sri3xq3vS
nlfTpM9dCMrxNEdo+4yGm7GIf1tHTJJhGM72xfxY/kJ136HXIDkamTfvx3HZvzVD3A4w1GbV8tYE
517mN+uYGkzJYdyNV3W96hLI8YSCfeLFGPXXA1EIGpp4H3p83r95XB4I66CWZt83okBV/7rTvL/+
03QC1UG7mJwyRwaXs+tgtT34+vZzpNIWfA0ZxthZtvJAd/zHr7LQDROwoyYQH6AzpD8zZj49gfhL
0t0ub/ifhUgocuRovKoxnIF8almzMoBCmY8hpE1KIok1YxNZRoZzpHGOMJAUWef92G0geL1xrfTG
d+eZ+dC4eszBeFpTEJ3QgpjIDcScA1zM313qQisYS0zWaKTksr9ZL/kkyIPqqiyN/JKwvO5xOFfm
KP6H98rCag+sk79K3jXf3/RF+OpQnf8SvrW2CgYU5Dyjl3XLHa2DKTaRZuFikLJFSqoh4o7tQfBT
IuZ2uYdGpFBabw5w5ITeRy9twhjrdGyDcs0iwRGgfPtu0U/C7lPqUBZOU32WmYF31DBdPhlQsXlU
tVOGe7RDKuOXDr+kT226jZWyTN2SCPzwOwmwXkbrVZ/t+Ey25miO/HlbWdK6qYdOstUedNCbjkol
1AbZNdPXvdyVmE9B3roNPl/Tjbbky/dD58CUR5OdZ6zs8595L0ArbDa0jSLWH4GDx69/aZoLfu3L
S3b2LAG5Wpbz5clcgOmDnxF9keJSiXr8Dzc9bljCKJjCyZEVkOLo5HqLEJiuDn/xfh/zMQ2yj72E
QUhLN+00lpv2uYfzbzjdxrlH5M6OZpnFobQHJ51zFFaU8mf2pTgFTs4p6Tm++YX7uivx/PlSMT6f
/iGG2WyslYp+L7Lv7lHQGQP9t1rO21awPv63ErJKnNHL9oVh50QSyhVJJr5uYcBkVijndWUAffK7
GMnG7bgAgv1eJMUx/rkBZQIQLk9wYBdnRqlT6Urx9EwB+Hp1Wjr+ZB3J9n5OcaQrQdJ0o+ABWx/W
8n3mWdJCvuJ9v7143YvQoJDiezlxbpNB7hxzHQsj3IIUqhBjUWly/s3s4ybJaQIz+g5fxbeDFzDK
FXgbz9gmqAjm5yaF5CMYWyVaLqsZ4nQ6QO9jkIAILRdfTF6oDjjaeRNoO8XND5aD0LFxyQ0r/2P3
KCGQT6yC369c/FZG/i9Ka7eOGG9tmgCTpBhHehO7Gqny5SJIADqwC+1jTPhGnwo9nNJp+LrT81Ra
oGvAN/9927zI9kMdMEUWbmvLYBiAepPhm49ROPoKy6z2ggxuj+FWRw0xhx37eHiLVYecU0WCD/Sh
HSSFSnGoER598EOgXUqv1nxofVNxknJh2PbwWYpKiIqSQpvLRw4AJ76csdGF1Jef5ZaA2S60NWt/
CnpokECAD0LPTQ5+td787XejFY4wwVhJ51IQzICtV1yiS3sgXG25dcLasteymx4V0J/2nt2BD9rN
HDX0uRr0rK6Bb+qNb5JhfmjgO47CyluHERX28aWQMxBoEtQom25rTygmKsO8u5bdl6qS+TIxEmNf
3a1N/iHLG/fUZ5+rkyDYblPUsa152fTLplfdPbb4g8vRJvPXQr49IqnomVtLi7gmbtE5jbuYQAZe
WDv3frn8sYRUWEpb9gMCraBUYhVyT0qaDUbF3DgpKv9FnATNXxruBcpjtZZ0FN8xW5kiKv+PFi9A
epZyeAkoCMxSjVeQCTIaZ6qrywDFsOcBmX26Cl5fTkhcNieI8UPkjP2ej5n3hqE/ajP3AzLTtqX5
4SnZgbBaJdxP9ANKWODenrAPdfxkYanf1i1rQD5bSsPHrnTcLvGBGKfOW0/lxf+4f5NvkT49tJps
KX6EhTRI23COOtGo/KI1yhokMSymISDa31AI4guBWus71JLQ3dhLwsYORCcEtQBSu+XiY+7BGkKj
39wB6/7uUUvule6brQxxfLsNagRUR6Epagw14HHJid1FIpFvYCrRcNd+TpwcprKY3bKz4NxUlCr6
zWY2FJpqf+IcaDE0c/YOHsw2xlVrOQDH8flZH5FbsP2BTilUOXvZ9dyU/4whTKVqLCwtFFSnsxPp
jfHpKtOGTuKbqrRmoTk46flabpoqEcckHs3iUraI1N2JAo3m0Q3qAaKdL/sEGxtNEdJT96dnUmfL
DCQq7Thhl7DAFaNQXLlWtIj+L0IjrL+BgiwsZCHFDanSlz+MO2JvtBkqx0pg3D+6BcW7USaykfM+
NgVAwgpWHT5vii42fOOuP/Slg5bATb4PVitACekNKH5Snr9/pt0qkLGT96l4e1UcZfE93FtzXOYT
kGooeB1ajh1AjJIMlqBiXgHfrs1b2gxbL2S7bYniamxBWURSbhho39MkSVCGmvcaJrkij3XxQfWV
AkDbzcvVTHoe4Rrp/XYRkP2mibxbYv/Gjx625PSwb5qpLYIEKNbWCgGkcAqtlsesH13rmX5egYhD
gE1wZXNsRDTy2niqKvbUz0Y8sjpCnmwlyPW3Ogvby26/BOC5NiVk339AP94vpaMZYM3ZCSywFnR7
ClD0HSqDCq5a6MBKM6orALW5BDsYxF2Zjn+FjYKYbyD5ctwo0KDVpCSB8cMqcrRPmy5OQqfQ3CzF
nfPUYk5wYKyOHjzLrD4Gn1prXvvnbLHukBVTe/OtayYQU2oPDcwUzWBQWFv5LlxLxlVmLuC718cd
oQAsVc/v6suzm81kQ1alvW0xLM3wXecTyjO4GJICiXFKIgaDs+mBtOQqIteY3RVIr/KjJmXMq2i9
/OdDHE584XWXbpV6/DYbeSCqJg5D/UCK+2ThovhOq3Cyep5/JcwMmh3zUmQqvzEMFlRTWdiPf55w
HGxVV4Wcm2VVTKtCFadMF9NuzO3+Pzv0Iya7XlOnMfUHjp08u5qN+awWnhQVFGS5VuCqvW6wY5Qj
rc7tTbcoUcBRthInA95gAe4mO2uETTGIAxAFMavpu+0GCEOzujsSXuNB4dElSNxvR1jbFi/YoIk3
MULoNoICOH12dmIb/0ywCqLF9pD/vUuaMohvYIDKPvTzGIWIkQv5G79TwEdGHd0P0l8yyZNBa+Zf
9UIr3WwzSSvViXV79OSxkftqb8TCSVUqRKC+WMOycss+WYVxqFgbPlsoFkb6hZawmz56VO53Nj3N
967w8r1nB/apbQueXRj9hMJvVAyHLZv3beLsWgdJicLPlJFvwpVOQ6FhOo1fGHzOaMmZk7Pnvyyx
fDllnvcWDMGSn0CNY0IzXNBWSBhgWXCEyiuegrIgL95gO0Jv/9oJMCUpBfCqPp+2X+IP3M/gUC2q
Xy2hb5sFahdVnWuP+uyOo9Fhag2nFMYp3e9eBz8gNNxHpApZQtOonqgYYwP6/VH5Pau0LvVoezXf
F9/oCw2CGHisHA9YzF6CEuwREggeePQB6Zt0kpG5LuBlu7zUGI2YG7wsmpaocAuDXIeFnIwOeTbs
REjaqeWq+HbFF172AwKLtVJzazkK5bZSUp1iKe0WpImd0NA1p8oPZyRu/nZPr4EeNhiUssCW+s21
kQHIotZIWqDOmkDgua7uwSgWlkyNn1+E/OZ1GTN35Zpc1NeuIzQJMOSLkGpFNYmvzm6IacmBe/2t
bXtuz2Z0OjXLVYlgSH9l1QsY8W09e/Azkcp21L+lopRzSPj65quyHs0arDvVVBg/RU6pPNn8PpoN
xP/GEEgiiyYJsisM5BYZlDnV0seuvaH0NzOT/GAKk8i3/rZ2QyHi8I6zN02IafkPvQ4MTe9c5Brt
nPHn0nKriHg7qvDhgJzBdiKW/WWJiovNYR8hi9Nno5GgzRISjur0rHOhF5MO7UtIe09Y+4QOl0qF
yqY7z2ad+6RQJdZ3AC+mS6uzZEAgV2ACuoTt2VUKsVvrB9O4d0cXVGhSEopDiYSYjCJ8quUMd3jW
KeyGM9tPIAJelGzx4CAIn1a6Hw6jtdM5Qq8a+5MyTlYvTDkR07uWNatEWkB/2x6/18VfHge5X0++
uljCzCOR+4Q4JAZBFS4EzZELpiiOeBeXD7yjS1LESPphY3UICaa3l5TwG8OTndvpxynwo6PW+eET
r3oUpszYCx2TPoZ6I2eNUUGiy5FNasGWGzzn8V5v+Mk9FIX3P7/Ci3axj6fjpCfBPSQ9GB52R2eh
bbQ0NBdlp37L7tabq3F0XgTmI6NFi0HoKsO7jo3McqVZfHB3+k5iepFmfydUGtuxqc1Z5B2qGtiy
TpxZetyV5EIuefMUCNVF+HpCVkdzRHJybsFzJnpovTSnlpUAwXsXQIha8x+BWOrIdPzuqUm5/zNK
oiEIahVSA1vS3MPYoR6B+4tljUYRZL+LfAwTBTJha4gIgf9ioSTWpmDYZ3+qLYjxkgImQCEvBer5
M4BljEzacLeZ/M1sfGW+8FtXsPsCQyYpcAuyaNKYaELwHm/2F0qDKQuWlqa258+4Hdr2CS8Ix9Ba
72KBXOP/V5Oxab7vYEZxvZ34PM9anxl86Viw+dRoI9RG1h9+NAf/TttMgfOgamNijwUW7gfPkE4w
vu9qrxS3GzxNuto/QO6vRsfN/dZagTqM+bKRQJ+fTMEmskaAQQMU+KqAEHyv+KR+3GNHQpaYKqIt
LzSIHE2KAhQDSRYC9YC/el78XeB72zEDbm0qpX6xXxRux5cy3cMH/Ik0ctqVBDHS0R0BTNEhd+St
TIcc3LTlibdLPYEH70KQ/ibQR5RGIj2xfQlp3QHCgUy7m9FcGSkJkWWBgnhJC/cYB45wZTHbyoaK
h3MEHZTwJc810v+Xn4SXsb9tZWYpV0Pq6Np9d7o3mzNvgHmp5ormiYnohS+XUNjtw3ALxu18af/a
Kzye5MtKYCWkaURn7+hS+vj05ieF5Q1pKg9C9pO7fsSG3xQ1rfCX74bfvoP29RKMfmjzw/sIXlyi
g4q9K6AA1erPb4xOjpZxLuCRV6e18JBdC8JWtBj1bL38NQ6eekIOkrVVHToxSudvSvuM1kj3AkIA
uDz8+iGwuHDxusOthF8uBzomYPirPbz5RuOIzyCqUbzYdo+ibqDTnNWZt8fmsquuaWDPpCuO/2T1
9ASRWSnz7MFZ8iMARHTIhrqLIfcWaQa5OwLpAHoVvWz9SM4K/nUOKPnmOld2QknNCS1kN+EBc8yt
boDnDRkZ32x1ixaFRfuyhJyluDiebHZA37n1psdk3qWKbQGZDKx0H1K5reHKqK3qYoK66BljbEba
xFKbGrAEKbWZtjcbuAVltnkgyCn4vK9DEvBxJJeqIQUWGI7VAy/8RRo58TpptUwUM0j2PoXFnVwc
gQAXGIsH/fDgHEkIUng+Cz2HIhNvbGWP2gZOt+YAcYxeHMG7+K4HynrRgNTWZUOIEIdURcM1ZpfA
3wDRueprrfScy7bP8saExwPCl5JsiGwOvApl6SYknOwpKuqmbGq3pHegnMcO7IlrAHb2AuFWM9RQ
VrZaccxCKTvbvdiMjXwvznRvyAh2HDAhPogpJ+kpEHljb3wC/S/gtgwoGoLlPXmWqLHgb0hXZSY6
zwNkt6q52XV417HBu1LuZH+ny7BzmIc2MHXXJnSiL2tANiYqgKiSbsCVI/30ljj5TnBqsOJ1ZY3Q
etzd9t7YJqgYj3krmUN7gHfrG2VsWzDuIgblcYoG+5c7es+gc26E4E1eoQQg8VzH2DbRL+YlhAzB
7UpNKYr7CWpFfIctb+8kNmtjZVJCAeLmWlb3SyICzruD6dvXvtTbSy1aQpMVcPXWKPTSqkEaJ3WE
ZPwlR69e248/2irGI0nYOjc81PmYM64qWB65TvLbjy+kQE+5qu7JPWqztnjR1Gaas3kzYNPCbT0o
xAkfeXq0wP8oTfX/ofk/t5mXFpTFAQ1Lw/SvkgoyqGAwBiULGCP+ojB5Kwe+OsqS1OmrwkzfgpgQ
qn4Xy2PXd0rFGDIDYgklm3rRpRjd/XkEPtE4lUKl4turj4JCec+tQKm4MwOBcfujosS4FrPan+1I
07QKN2GJ4PC7KN3OMNl+dxXYSeeTGZbV2lU/rHbcO0wn5sgM/sN3JA1r8jFUVbr1icsWL3WitpxW
miRqgyjfRfe8c0afTIfOQ8NnK84t94sVMGJasz7/073cpxVMQtTqY9UTNvdzjYEJA8W+k749VHiL
QHjfhx4OJMuDGg/xxlnH9m/SPqQ06t1xy7wWUvJYFckpt+XUa3r3XvZjH/s6hLjyXTktLmtyvtq+
F6mQMLsHreqHV8w0iul/wuyBX0FFZAxabt6pQoTUl/89FHtEHUezqtKeQ50PAZqCkdhzopeJ2mUs
ke8fAXWCebzDpBPfP5nBClNFIrWIXLgTfSspWvdwKDejc4oWQpRT+abruDp1aCiiLRK9Ndg/hnpl
REtVqUABTyl11cPM/6zvYRIsnlRs66uLyuFcTaxdQOcXH9bKgH4U45wMm+0g9Gp39jyteusyzjba
9bfUUv9lg+/Wxe5UAgzsnN+lwLCF9OZi+Tf1DE7SJ3USMqfj4jAyQ24ZnH6pZzB9n9Z3T8E391xx
4mOJYfUM3/vvF/stkhKrTV94wv16OvtX6s2DUGDWyfLUYZq7TWEB8GKY1JW4BeZbj7HxHGfTmWRz
S6raCxmfdOVyZGivOzYYOPqMo63qipKIK5GjnWPCLrt7e2UVExMGmlMArj9/Mq6rwWgzrKYwC1D9
R4IozoCdky8+7cWtbk9LUMI2M1+Tl4ggCMRASNboMyA5ycYvk8bxjt3fUFma1vfqcrlCtsWw9r7J
GKE84IONt8dxta5HNmx9XlJkFqAjkXhcQD/k/TLm8Rw8v52hoitcBYj4J4Qa0/rZZoG/kM/spoSx
M8OKp0yuur7BldQyxp4ljejppb3m2Hrbo5P0uZFuVJBuT7sziu9/R0kcY0Kn0T86B0KdqM9izW8R
B+K7yE1E7Z3W8DGWiJWspl0+c6Fss7J/neTDV1z0+6jN+vNCg6KLlhakS6UDjR9nr55kryxCIaAd
8jPjY1/VrEqVZOEmuwyFZ6pT7kfftDeRei4I6ZYDO802GJzP1+yyx3ng2eUDgRLHiGDb9susPbuY
NajO16MmXDCIWkFw/214hBhozVbMQ149UZOHxIH9R1v6Y+tRAXrLLVsk9hxfNPuIUMekHikAEWRl
nTC/HuV4Zz93qMPUnE8trUv56yezCik3rBq6OqxnqRppJxWSOAXzz4DtGIVBgAd4q4OKD8TGDORr
cjp6DtCmzG94QyYyLVWwQWVncXbUrlBbuIeOgD0G8ekA47uEPWRwp/pMjJI4PvxWS10jxVzebH+9
68N+NvS1k2vCFXbgh7xpKojMP/Sz+gn/8SqXonn+56cYEUJa8Tob+vrvvc3fvmQqejWzUbkImsQf
W0e/KOf18nE12Q58QjpWnRyv/RZbNDVOoMMb81rgQPW+AO2F3I2GbzOXD9o/NYfI2z9UNc5fBX2P
Uk4wGIdyl/M8hj8UEEDJHFhk0GPKqmq9DszDF8F4zkE+y6CNVGRd9oEMqbRI+Qwubo8kwVwiQJXo
QzU9ldMXkVXGQBlsT08dm4dqPDaZCwnAu7fvQ59FYUuLGP6N8prkB7mA0T+RxwevdXltmLc2UWQc
6zLrLcA+lyxc6YVWALnJGzpuX97dlCYjxGjDk8NwrbGkT/FE7xau1W1IGck0B249IVG23pGmsYG1
JVhUMSvWb+h2c2fIuGO6SQ0AEPIc8qY2ZnNlkasuaHQMAquOeZCkh0g8ypfrkXb4bTdrSRUBz6W+
NNhgkoqGKAXdeME8/4d5Qp4tC/1bohcb2BGzgawv6xcMNgW//50NqWRIUZ+ML/9MfnVxVPszjIb6
ulNCq+aOhkURe2cwuATEwDFEDNFdavzrpNxzRds2tvyl48TvlIeZ6xG93v/T3xTrSnBWati4gBhg
H6KmtOt5QPBKnQG9tOF756rr4TXY4NxAh/Xim+kxzkPEGN3+PB1JWfUNxsFgzb/bRfXIdHYKiNRL
E8fiCB4+i+Gb6WZwiJ3dGX1CMaSKEPcG91S5uFy63VgLBWMe79ZIE0+DJWjUg9N6D73dKtcNMQ9s
Yqx4Q6G9QUCR3EFH9AyqFP0w4w2Il8A4VuSQOaUyFruGe7/cvvFM42WLCvaFKCDLl6zNc8BtXcNi
y2tqGd/OxQcTPeJCfSeMD3BbHLiE+ARdKwd4ZWTjLfcW6azaJO7fQVKI0jOpTzlqbwJc6FoLes4S
0sDXMXUhAq0bQmJIMratEffRxK9LxIwLKW6tXwWsg+wDrXgCeztzPOjDbOmm/XPKHU9QUohO4n3x
lTMvRipaVfolFwx50We51lVEdhzU6WOVHk3xL96CoclajMUONZULQ2QeTLvhrB4nSQzri9qzH2Mn
W+ug/aLWVLlDqNG2gAF6hyc+iN3bHoFH4B3jWXRUAlP6FU1LAeopdUaZlvgRMLgW5KPZ9oxdvAqe
fhBcquwlWBb2iJDWbGnsGlR+sV+jcoBWelRYu1h/WhufWVvlZ4Gx6Oa9JV9HFy87dvaOa6XQuMx0
I6ehGH3xDZYQWyqqPWeNt7bjVE2zwJhDAWazWIPPjhdnMWAT6B+kDJrpZqCsBLsh5zc301C3zHJu
xZ8q6HIb9/hX/Xb2f4UdIu2hgqNXVqZe5foReG8m7w9ObuuXmzMt9Pq8yP9jErS/zIsDesbY1Hzn
JALcxJTcJeTaxYucivaTjAER1ISrWxQD73bw8UnHe2vy9BrhCp96NGJbsCCNjGbNMLPnBrG3FzpO
XXa0IMY36Rphtp5pcQcVPXJe45tsmPkesU0/eUL4eUGMkUf26bup5r7uy2dTPcD76/GOLTLjVDO4
GXs0pVBYKiJ69WVw5EWAbi/pJQFkRzb8ULYQk07TJosPG7ddfxo/8MQ0hbuZTCcaaVtdQ9TI3mzl
VObEOUgDuIxiR8kSvlKCEaxIqHXJM0xnNFi0J3/et+6dNMexQkLYJRg9J0VvWHOPGdQ49Xtq+oaY
LnMjuU5O9KD1gcSEQ4P4AIvqVNliIzqFW1GWl/8J3CtK5KEV+qapcq1EW2z0IXD2r1R+WXXbI87S
qXS5+NHUs3y/3u0YFw0OxlhWGE54x3osRzOyg7ymq3aRY9WLPLcQ5kSjax/F3cSLjtAQ+2lshnR7
oGa2zWoul+lXEzHIUmslG937eyuvJfyuwnvQ6oRIOqjeW/pG1HYDmEyFTiVer0KwHCnoma5+vtDg
oSRqSGMPhHIldOsMyvXpDrtXt35h0HYVOE7Oxfm03ndYN0M84LHCtcRJIr3PUViuIWYCxuBG6ecG
7DxJ97aKUF+NU3SHotAJYLs7mQMTZkDFpmmNJQmK6QcWnD9wdbLNt21saEWgP+kcSl1xYWfIk+lq
yJ4Uy1G2+wwCxlJqSJezV60L8rqqcuYt9p+gPCYFOokXqXv1IQRdTFyvAHSUt+zlQOmMV3JRcDdC
YVO9qsyN8o0qYZUuJcHqphozl4IqI/bBmWmcse3YhC7W93gebklquIDSOy5TEmP0tvp9JSTUtcI4
jrmOLigWrqsvFNA4dC47jywoO6hABu1yaj9zalC75/1/LaP4WHjtk8rJXhbhdri7wLwo36vie3sz
0G9PkzrT8n1K9hrMdTPI+ePd9B3H5fI/mDbDeRtfvspJ10xPzmeHTzDLkBfPJEQnouujRA0f+y4A
PBK6kslVzV5tpJL+bbVk+LKMrlhy3Y73GTUoNp7YVNTEtRPinHkdKMXS4GKpdpg32pyi1Z3o8H3z
E57/vy5rOR+1SoWHB3OEnjrUlrymFogFEyYDLMb0VcpnNQ8EF9NNL8DsEWWqhU7c4FCXACkpHaoK
VrvIqGwL7iZlEx/4+CWWfX47yY+7cne2ahaVIPIz5bXdGYEvYAapUZHXU4XZQILGe7gWY+Zb22p0
otJuidte8ZFZ1Zp5LBGWifTscUluKfE9+gx2qkKMNQULeWn0DharCJ3CBoS+cK8n5/I59FzBxsQv
tWMa3eyloAOKFiIHu9QlM+vI7H/zEQuvj/WOwtxS35VmPj31C38RpUP3BtDYjP0p8lR2j28TYMyX
UedCZXMeOHhtyy6NdI4+KFTwnojo2uJlXLlD4iBkkYDyKx3kvqp+noK1MQ+jo1zxGF2wH7wdXvE6
GtwVofA1U+TJGCRqmmkaoQil66GX979qILNpTNLgt33kgramBY5L61ZFW9DnX8uN3xV5WX/+ptr6
e/xDO2VdSETIlaMBF9WDAYJZRxsbkIUZr4IBDDXYG5ZMCNz8iDj+0ygnHFc4wDSvJ76HgZp9s479
ImsH9ZMTV2RxCyBriMA5+qV+lSK9QxfEu3Zcg50UqOE3Rt9CT0T8psDeccHUxgGf1nAR4C+XdLSN
46R/2mBYAF2MNnmwD218nSVRfYxsltaGbS+k/a1D5AtZJY5/zN9V/DuM06NjpDWuZbsbpgd8Li1k
isO9RS/2xej99Idt/jqFX/HWlk9pe788QVf0MBuz9dXE2EjasJFoAU6hxngw4qr6qW4DnURkIrKS
ODjo0lAdWOClPVZeD25ueaqe22l1HC/TNtZjC6p09qGY/hxGX54JQkijc+xGNH1731tg5EuxMbAm
glBfP3NN2BXmMiNUhwklYGrexRU/zTqJGy/wJSnnuGFlu8tGcBS0S+iWY9+7FIuaydrlFGuMQX/W
f1ijyBTAhNE/c7n8xoM8w2YypYdAwuUo5+aEu4t/Hl9FydJCQRcw4x+2LeKtcF/jPAQtQp4aukpN
7Dv2Glxfgfy87yLFFFub0VJ2LZdMQwqW7YwSU0XUYPnlbZdLUxfeGml51uxpNysl9B8E1Ope196o
y/yxqLyu98XIFwJx+h1VEjx7pwuCV+jES3FG73PwmDeU6cBAWHToGGtv0EKPALykXVUs4Can4c0n
3MNKx2ASZXaEibdHvQUfR+AqETslGpV31xB0/ADRqVQOE0ZXrqu1XyzRdRAvqoSa+dMMlvKKCzlk
4DhGzWSM7F3Aa3z+5YLsLJiizS3WPBNLQySJHfA7Q+pZ1PhoD53nnXtFsjkjflIuD9uvZ6VgjB59
y4mJuHstqQ4XRlkQr915vXoYHEz0id4L/s9Xa+DE326y1wTV+5vlFukCX8X2BV7w8LCx7giMoaz5
HvBClY7TvdxJ9/srChV+qyBKsuVIVK7tjR8sdficZ4goUR0eUTQ/HpBRKEL/Xbz7PzeyXYmg0cHK
+1TXElWUr5yRmdT7S6IkDvK4nz0uL5RoilzUG4vjVA0HNEW8cipS074+60Q03/YTqplxZkYsVeSK
ho9RVKTp5s58TSeC/FAPcFdhwKC290hSFlsfvioj3kPShNMkQ9PSTPbVaEqA5kb+mdrlNB7Z4+pn
V1R3YJ762nL5U5jCMW8GGB6fLZNl+ZGqWRg4eHt/Ebmv0bfWYhuQklBeprYnDuTsSZBvKzqO1p4D
kMEhhzTmlWWBfyNtaT7LoRYdRFUTcV33b1aIFP/tmuVmH2kdQMpJ/xvm4ZlDurb8OrswCC2Nvlbt
nTDLQ0a7IhnlHt2SAq32dYOpROrQrWpEsF3+dHZzsDF13M9hWuKi9DPMuB8dOWW6t/2OR4FvkhtK
0jZvXqKU2XSKfCNGmxZu4FYs99eNxqRtiRju80xe5kxs1p3N5EKcNt4STQRUFGrqwT0UKrZvGZJR
Rccys8siZqq4aHni7mxoGt5PHXQAoNKpJvQD0SWnYlGLdPTq5GKP7OiSy55Xfj62/nXLuhY0stUw
fGdXRqYw/J4BkpaX2p2OcR/hElQZVEMi6PV5JfMiJmyUkKcpP6U1jHqHC0TDn+zNJQDI2hpmG6pl
J5aTmAMVc1syR++KUpst5VR+bI+5ePKjo8rXbcJe0YDYqhkilJjYOL1t6F4NiIzsOSnLx8tpbRC3
U6zG0j8ZtdnvIk1+jssUj6+JFeOtk1y0VC5SfjwC3w5FBngluDyzjtPpbrAI66A1fRmqiA+W84/V
7eiya4a0+GB6CtM1LLogcuAtKMTG13qs66CGCwtVLRcW6ZMqw12GsH5DQaD6J8/+ecr32UgTXX8t
bOP4XzndR35da3mijDa9r2KK3NEXVxP9aeqsp6it5kPra/DtQtLCVSpNfHlfD6koew7zFod84O5c
CqY9PoGGGxyJaN+RGqMFDpflG01KiMNI8qNnsR4WFWnauKYxJcGbNqF7P5X/LuPmdMDPOjbF+p70
XRboHm1/NJRDSg0rVQEP9MhVgpvAQ1+dlRk+ll3S8n9/l2mcXRzpLbuQjx/5f67CPAneImUEq8cn
5O9RC3KnEQfXafQEfNNsa/STjSgJI3P6V0/V/iSK0bVTkIPvvPcCIZ+2PH7ervbN/NTIMp+ZtP0M
pYMxgEy9CFK/KKXMqLOFq3YYemqRdaME0UrJhunNeRoMoaNd1Qt2Syu9PNFdtbl/2kEAPQ3JE0o0
Y5eqvrGLqAFtKc9HFM/0mf+Yj99yOwYXykiF85VoPf6JCj2fu6qgvlNtU+5VUu4sf8x8A6jB+LzT
J8DUC6Q29LrTxUeQUoWaNrRlUZfNXe22LIAlm0YiDf/uyeDsMjNeLVHd8YNe2pU6nQEQM0QILF9c
IuqoFHCXTjRCf2gXeJ6eYV1mzKmyFPcEWw1w3g49pVvtu3Ma3mrsHm8usNLZG+Xl6ZRtr03ngZx/
AaXrClctEOlC20Irn9LM2FY9AZGpjrmFuz3ajjVQPCNJu+sYV98iF71zyEc+FaLwXmxC8t0PVPuz
nY9uqez9jIwS/oy6IMa0nWc5Mm7+ze3zqiZEDDXnjSW6e9Whn7A6EpS35WJsiccQxFNdcoYIrsPk
u8LxcQojTAjKtct5h2R+SKDPXUu2eKmCt7i9O4itZD3VL5n2G75hIUV6X0EeD3IsMRhSKMMp2R+5
FPOS71+cwq+WnhtETc1UP3x9zuoTr48Zi5rMeADvHlgymDyRMN8JD3b3RW0IVPQd6riO1UXBmIJt
rLu4yJK2H00RHdZEvTK66E7vngSFeHCaWuS6VGXuIzhHImFkOC6vdhJlt2MqFz3zIz9LJ7GxcenV
iPbDOkgqZOu8FFbHtb+BkDxbTCm55YLSH81M3NFdiZ9vbDQRPAzyfL66ZGbEaRValFdMMCre3uOg
HZ4Qykfa7kdWIBWtcD4hYwjHq5UC6yKYHUMHYaVMVxzQPtC7vhe7JNXQFEkUMQ4sbsHHwlZGLKN3
ZoR0jz2kjhE8ygS35my9xRvRT5qamlH740RnWsevqbtWsbNMLjmDgsPOYztkPsucOtDGc67/NZqr
aXUpCIhtZ4Lt0ofzdJ9mEL1y7gQK+zTMsH5fyFPdUedrgQ154g+Jg/84hkwc6htM7IZR3x9FUYAZ
NRdiCeGiRg+7bUlr0XUpqSryx2yGVMZyakQNDeR1WWiMoV0gwNdVLS1JAY5SjcvvDGI+22sxw5vz
swKQV9PkY0W1PKootoCJ3GyIlu4si8/ct0D4SRpNQR0mdHaJ/XoMbK3R2/ArnxrfGyqYKuQsIV/d
EJpNHnIPZ947llpxU+XBCSsWlY4kksAIxrMzEBxAxuoKNZajiy8Xg6uRYIrnzAlXMvS3PW2jYBze
3QdpMnPNXGhfhtOIKMCOm1GKmlBH+SIz0nvI8djOEMY2WD0f8Jho1GPSKjHMw0OeKI1gPIfqaWWj
mefNWNHUdLsmAMFIHs960AF6b+3Ql9euDsHsQj66zosBWirbh5VLv3nVzq3oKgz4/Jw03q9BWpOn
ydI1w2vdCqXBOJWYfbvMg5adoOWzlpdnoltROfhmvHppwrROR9Qc6B/VJhNYNfVNoPfWmMFhMTKI
yB3BBzzBq+iTxsD7tABjWzT21KKAF5qgy0AH7nbceTg8OzVLg27OLnA5oiQDIs12upzhHYmCbXIn
d1AQ9nvhek1v7eF9iNiJHN/pq/voD2oAAfvr9ZTR/zJbj4BJ5L3cR8GaJZ2bIs/bcst0ltuZ0Wfv
wDzIhR8Rew7X1t/Dm3i/IpPnQEWMwtfpedj53PQGzSyFrxhitZBWEfyT3PAZMLEmNpiJhfj1Otc4
zVtUKChnDGl0XD/u9BG9X7t8ESAHzHdKYeys6XpsgLrDKd00KykWezxQO3jEGDMNR6RsHMOc1Fog
3ISW/DLA7NvGF4HouIpOzgpK70dq0Gc9Gznsofv1ftjfwGOvCUlyzMYOlfVcnIgL0INgbVLOJ9s9
WN5AYcTB+jA307fGjMkmV6ItbaQ48pvbNLF7/bOOOmUXaIXgdamw6aJgV8LbT1XnE712xudbazWz
J0yetN5HDqIs5mN34Lx4TWgMJlY/p6qlL+z+NDB1XRVaMpDu3cWk/jfavYTsLyyKjnIhvg6D/YMs
NNroAcpPpKYKMa7VPnCC8CIDmjPLPJL5g91ZypS2hsUV1MshQeWmtfFRApFvJzCMT/qBIukqUxw1
1h8PxS1fyw40j/BgyYNRuNXEx4OFrOz5TTiT3WXbIm5Bz7BWCmBMvr68aLdvFA5QdTnDoz0tJHHL
dmFyIy3h3snpqAXY9fQHvgw26YpKdFyNGEAB4sK2NkgrZ5J2NasElM+AE2N4DFH7xlhw7LsVyrKN
7G+u9ZMd97OZxZ2vj+M0FC7nKymzf2HmmmEXrqhQV2JpNrKMQsN50CxtFpJylYLvF3n1RI+VG8VD
31zz+Juhc2KmRr+hzKmTjrOQ3BcWeFprWmc1QvyhpwsV+AinTQjJxyjvaeSNLvKo+TsJKBKvWNv1
yOUrvK0Oru1I0FwldWdtOmOmR6/5MYl5azxYCTW/z7+ra41JRl4Io1kitvblY8IBAG8smPhhREHJ
EPhbt0WOKLsHnc8pQCP55cTg5GlcyHUp1MiWsiEBNzXr+54cks2JTOZLC/nicjvXxM/V31inO4YX
QsegAsaRQU+iU/ECpXEmBeAJ3AFqKdf7m7Iz2SDww2y5gm5mhVmi3TJBY/c88c5Bmdp3GMiqCX1K
nHHzfjIIaazIZtaqyQiZsZ+BP3iy33ypYYkEQ6axcvIMUiJk/aKyTJTe1NWshRgsOOPidofir+Ns
ySOwNRdZSD9KYSXskXasu/RcUUjGT8wzhbK2jBB6mXbz1h2w3zH+Xu8k1Ru/3yqAO4Mr6g653u0S
aIg3noKf8ZDI4MN1JsAUkudwQrYxp1z0dAhKKxFBsrQ+13/3mMwv9vvi7h2bUiMlJQvD0uOcJBF6
yIzUS7nNLlKqeL94szn3P2EsyO/FYjAXJSPjohp3HRad6tZzNGoI0JVLA59X/qw2myXIEz+eqwU8
YYDg4NynMQ4GlCHIvdBHUAViM2YtufxB1OeQ8XOCkq2OM1On0xkkJIu+JnO8DRoK3gp1ceERyyFP
a90WxXTkECuYZvXEBJze6+WCpc2bxcPQS/k4iufzbo0KY2g0KU2mAtOvjTpx9MLVRFb0iPalf63w
MPs1yLfXeXF1pNwwAcuEGM2fxFAkpzwO8ro6D6EyqSIOuv6PBQ6k2jfKNDcTZIvxS7rHYO70m2Vz
9zmiggxfGk1CSsrfj8r8oWy/jDGoGQyyK6IUaAjUiJZxnpwY5ELNr5IhrLtPD1zYS1OgESpX5DfJ
rGqtogGCCZnBEkoOsPvQbxSCRJNF+iI1UJqBb9Kiy0xM2rP7xtyNIS8XP9eTiWEfvg2eRbdmIWsA
KxKEwIoTUJhvLuNFVIH2fcf7b1kpsSouk5w/uIhWNiUkv/39aOCMa6l3uAB1wHgg0aaCLSRyGwXW
t5AMn80JnZnsD08KXLNoSC4S81L/br92Y+Cj9sa8LW5UNsmduWLcn5e+LPJV06u9221vNPC54zOP
E26MaoiiOCS1PP3a00Je2oblXjuYryE0OARsWoYkYEVgMAj3I9QDU3nPH6+FO86hNkbDoFlO1V6N
Llh9D8+fRF+lEKgWpDKC9qebBQCPzo5ioVEWNkdbO2P0b0KS9/tm0GQzBkPA/mbvgxs0QZIBnSlu
Xwd1VucP4htraX5SLYcbVfbMk6qFvOWZINDxzpZyqN7S9+3nP0BRtVLxznX1BWi5tWTx8BCcW5Om
N+gIz+WTBumUTEAK/wNqwgQl5EkHKttIxyGWKL1A/vNQeNslZCzFrT/8j2JdjaseTN9wUJnY7E87
BQVwqxJzFlTfprxQa+Q26Jj6U7REtG6bgFGCNyMqLcIiCeYnCqYagwmDzm48yEdzCutOOdbTECud
Kki7zK2Y9G7HEdfP0rPVK5YxtkpS3LJKCcxxwUtDGMTOeNn0W9UJk85CLy62AiPabNN3gWaxWHy+
vjQFIWoMDt77UeV34hadpPI3cTa1p7rPhxJChYpoYT47jZRnPmoMvSnrpzr1CZidJMDWaFMrQRxl
LT3W4JYqHxkAf6k/uUt/n9bwWHm/SOO0YP4x8pxUfRqe0EhNMJ5lsw/msU/+kMXIYho+fjr2AENO
MCS9ngPg2vomrQDzM/w0XThTp/9ddbedH9ystuiXPgEZFjxil1zhwceZGzMhj1ZFqkvwbGS91VO6
kC+4UDYWmX/74HRSPQye0IfhWUEuUa/J2XDUQZEQSDl2xgPXug41wB7PfUl8Wv7+JjWHp+fja/7n
m0gdvtSP+myAKOIaxjgoMwfnHvbo6ISs3q63me8Y1tSokkmpTIYnBuM/ejImkDRg1KUcexgrrPc/
D9cnkRMxcmGjOgeJ3xm3Awv//X5LdXLEwMAL09i2QCjIbMyt9o1vUrVA9FI1i65TJUH9SZa1fn9j
F6qTdUsgecQgneM7wt0+xIUUjkdMqPDu8g4qUN7Cawg0YuV8eCJ3ZMZ5nVve8MJDGFYVwd7VkGvg
f5nuaY1lA5316UcW92lPX5Kc5NVfd34kmUK5y1JjeM+JJrCIJUDAfTMcoAlp0atuizCDzxG4fpjg
o8r+fYH0lZKN6LR7doeU83OG69xqyTN7UEoQH7AGBDmqiL3FxKmaSFp4GCTi5Bbcea2MJ2LSXkhW
VJsiyXJV7ImA8MEjZWxYeaCovZs5CJpSMOwrrN0X8ytleymLdV8n3RBjesOohAVhB+92Q1TB1c9z
EQeey/U3PUQOBYr0QoFlCU1Zrx2myba68ItdNGNuffXjnopX7yG2+zzfhA44XUqoBOHIqsTquq+b
+mJLBn9Qm/ypqbRBu0he4j0azsGgvyA3fWibxAooaEg/aThcPW/5WrzCW1kHvHV6An7E7ig+Uj5H
Y7jj6c3Oho4hKlrqiQtD7MV3G5pK57+ZvLSg25hQnkKn1iiJViqWrrjtONeArDeeDxKB7QQvk5KC
btZYz2RH6YtlXmY4hcp7pbsN4Ien6yB3rES/k1N0QLoqZmu5jhzA4Setid5CdMh4C147YMFpkQYo
bmKD3uKDakEm4wuTt/ZJYLdhEPrRWDlfkTUvBrLAHsyNoVg5Eu0omWs7sSEQGf0IKgzusbuPFzgW
u/LjkeqXcQJM8+pL2LPX0xdOEDtIvIASx6YzP0+a8eu9UeoTZuCCaxFzYq9st659kAR3wVBzfqCY
gfqkcHC9KgFn7NJ8kcfJYqX2Zkd5SsCC9LtTS4Uv+qffm5WiTFgSYDjm1Pp9vlcaKF+sJ/Jvmp5a
Ay9miSFIEOCAozH85krKB8JWkM9s/fXrKPj8CBMVZxxUjQJVJXurHrzcv0mv+fhqQNa0LB7za109
Umpmrfa9LZzPEfp/mhq6h9/5d+MBJRR+XCkpXb0AH/I4JZgTJ8ipj0geEr7OYwCi8VPhwoYK03n1
FRkZF1xmTD6b1qmvnnQeP2IxA4B4L1/B2s6o16A9nBCKQBsCGcO9wWxoYZiIYBeQOKbECTSrZAvY
A3/yrd200qnoZl0uKJ/8QDbIU1YNQjxCD1nOqe7Fqj1niPURZf+dkZBozsQhmEKe2EidNA8k3wTL
y9acnN4Ya1er7O34HEpF1HgHk+qi1JYvKB2VFndpM3JPTZAarXB8HQDwBNDjKeVRzFdwCxHCGDwJ
IXo4mf1q6c3lVpExQNteQ/E3f+LE011b/x29Lsi5Wt/GWNEhvaPEhIcc0d1ZHh+gC9AjAsWKrUTe
BfXnioct1rSqKsc6UqkurM/IVrRUdZO4m4wYgAI5itvF3eZt993iPMcwzLXMLdThFpvahCLGqwu8
8j6qSmPZCeLFOQLY0W32lf2G2bHcDwB+PGxe/WIaPo827BEx9nHJJHIJj7cT36OCoxyAfkg7J0uf
Ur0WwPdgqxTIcU0DiJA5Mr3lMzj0Gdvb1U1uHwJ10oxPc7jnts87hl+T4NYAPXSNZ+jqMXWVkI4H
vNlyameJ2YKY5J3bIHHiMIIip553uD/TbGwWr3+XjEypI1qUdkq+1MHXjd6OHvO7dSG0tu+dTzJ1
4NLS9P6ObNMrSANfGKvja+n9SHss61v1PFKdn6K4XAvuHdAvX4Zl4U40UcUHMkXe8afzAbdlHYRW
NG0P/Z9o4rUn2ikCmhMnA8brlwFBh3Uw/iyVYCl1NVf0qwOvLF0tkmVYabXQf02ysScIu+TpK4XY
A/muWryR6sdPa9EMm6KPutwgCvC++a1bQN5NNM5Sc9NT4UiRtT1sfIl2KFKhI+5KpNPclx9597Tx
hFI9lyL6JaLoOp29D1nM/FcdV0aZ9T2X2lDUctE0uIbQbcoFwRcfdCgFh0yGZjVo5i8R8kPDV4jx
/L2vgpD1R77kHd+EYHpHkqDCoOKj3p/BF1svUV4XyTCwWlgKqvTt4zfvWTcLpPy3KwDdVVh3ZbeL
IiqSCIfjcMrY11xRGR1MoHzLsAwIi/1+SfX5a0qxrRh1+59vaJDYq3WMNIth970+KMCuc4wrqdHw
b/3lCmC9FVdHMFk/DEWNGRgx1QUKWdIpKvURG7u2W/BJmJmzbA9NsJkLH7XQLiQ/Q5dECgxfjO/N
enAyl0M+TAMEpsTB8uL0e5MQ8jv/ONWHlzYhg79ZKFiR2ohfafW04OXJ5/1n/K/Rbr/An1Xfyu12
VoFWKn6EB6ZdZfsNqGZq9V6pl52lKOL+8Ke5gcSnu12IvXEZHHK6qBe2kr841bzZlAyCzpxoXVqO
aRVpCVxzlKOzwc5WIV7RKCvLHwiqgWWWUinV+y/Z3NEkRaD+gSB0gJW1G9P+HpM7GfLfKgVIokkm
k1s+ZAtI0ZqZpyaV2HD12o+ZHkO8hY8SDIXRe/m2pgchWgHRrJQ4uJFzH/pJqNjnFCQ+ivN40koE
lV378yjKB6ZsktMpTwE/ZuiOSo3bmcYsjMZNUubqS/mOny+1ACx+V0FP8uJz6P55fVOk1CaDsvOh
s2+3Nx76C+wmxWmLIwRQMdlwJuIYeK8nddIPk6dwg3c7M4FTQT4xtJdik5Tm/AukVyqoLQKdesWY
DqBAMIv7wFzArgPkhEZa1E0JjFDkfr7FbpF52DDhyxAhN6+FTnP0G9kucPOP0yzUC5/fNkdU5KLh
0olvg2DCaFNtP99j0NUxxh6lGt9scUNeQarXrzggD5QgEXOQO/J1SuZdF/GXfCKzfdgAQb6gMRh8
E4zsqkDDz0fUzx1EQ7M/lTNthAb9yAVrUa9qHccICNAfUpAb9cGe5cWwkmfJP/2feSC5c1iBD3GP
HBNkYyrxGc0/TBhrhfokx5u847Qhk4Wk729P+a9zJOtSw9UZQDw+wOpi4fmV8kJgbupqElW12F/8
5849Tqm66ixCFu3WnWi1Dpost1l929dQODH18BUE3/QIGLWs8cMZyIVv7RXdhYmlaVSUwiigONif
yN4Sk2P9gapCtgI1GZOeKiwyPB/coPZoIo7lEruuis81TK9k9+SaWjfsOKntkVrhb0bXXKPkzzud
E2Efcc/gEWdW9luoTqAvPo4n6kcpt/cF9UW5Rn1oIiMzs1hTNNawFCCxt5Y9sZEPud27Dpp45D6B
c1Ka/B4fRq8PXD46T0MpaDTRxyCOV2nCddNg3tLBcwcnpIdwOWojc1LtQazrIgwUoA1x/g4/fcfp
xaeQrGnoXeRPUkygUxuV7H8JJrclm39kg61A5wlUxYuq1uh75czQ3ndLHHUTJCjFxj9GJQIWfglZ
QeUzFBz2yfaF+CAgB+0iwPixfTU2ISH6VKHKC83ReJsxpgZu1fpZM1CUSaYv1VAvNQ/Pd17I4y0L
Vr4zkk4FEwODL4JbEMwNddUbfzO/jxqFxD7OfpwNf/LORRug3TTgcTLYC/RSmUSx0arY9tH09tCj
IEvYBVJ96BoD0SQNyzGbP0jKhrVSthE/Bm0snSr8Q33m7ccegQovp8t4yzewg1q/FNC/4tWcSYns
7xN9eMEZVx5W61i5h38hD9hCsxVdYoCxF12+aawcwvfx7ErDXUUPsRE5CjRKicaSmUxQQiWMve0N
m6brRlbmvRl1Y5ZHTzRTe483Ud70aTcwOYOSJMSY11mjwxQfxRLuD6jOa1xrK0TMl7nahD3CiYm/
oNm3NBUrhHr5iMKS78qLn0HYwd+Iyw7Q9+m5KMkwPnAF/dnN3F/H2UKyZPHnil74ZACkfEyzR5Sm
Xa1WiIwzDXMkVFP/rPqCgsy1SCR8ZqDw1rhzlGkl6ZJKf6H6xU5qwaY2JYy1mfYWymK3topw9LqV
HuojrviG3VEskzE4wWIjv+IVq8S90JDJc95Cdw3chUnZk9FR6oDOxAQGSROHvGtziNbDKUo5P+1F
i+zIT8ufEaMQZg14VNHYhgQVu18ZLU793XLS02oY+cABIqRJZ0J9LtBASAS44leq/WCSvGiWdp9e
zrxpfatCIQmMCSwHCu1I8Wk2GsF5HHiOOCKtK4MUwEyMSklNF9g3CWvSczxIocRWdYApuPmoEKUn
ZLraO4ZGbKrMX4ORyS5A+uuXfvnrNEZLPwjEoHpCTw73L+UeLmGbG9VoxedpQ/6f2RfSEdAWtwp+
svqSHOO107lltEY9hoB1Y0qkv8q2fPC9IR5V+n/sfiigRAy/QfAQc1bt2MFXRUTui6iUDDzGheAo
1I4n5lxF/EQoSo2gJ12hnuSMClnEFZOId+h6Rki0dIihk7O5LrrUEHTwN2nGsNuz6YWg4PHRX9Fl
wBrhKyl8r1CfD+oe5T8INql9sas5Dqls/IYzVRqK7mK479T+LZCugadIoHeUUKwbjN1cvYVgLFXl
yFxLtLkYHeTc5KgRzs48D4tCD0ZDEdomiC6cA3WR4eHFzOHSEXi+qkXrTxsamVDd/acQ/tw1HnTI
+YupZ4dbO+yVEyuGc2Y5BYQQYKy+FdIoGvVm1eQrX8eLSJKAZ8e3Sy12mAbyAgBBgWjQRSrNeud8
P90ULQBz/9WoND2l9AtftgrACHtzxYArwiVrgOfj1J06aO0vC9nBXersDVEqQcy37Jy+vehykig+
s5tXgDjaNSUvilel9duCMWlIEaEQIimW+afRSXxAwC0bPrGb8irrytG1gTxC2mOQawXkFCz5/hYk
R3th/xXpjDix/q21+LcCrtfPlSYx7tpMRHX3EM+m/C2+QZHd6hhteYwTADSBK09rzO9DFkoRhIBF
55sPzt5JC+Lv6Sq/SZjdPulfkllrSf8BSSUvIjJ+S5+xgL5LTRkZpKGd16UvYDST+OJT0y30SmwH
svd7+U5wtbmu+F7EjZxzVflP1EU9gwGJYNLsDXs0GXEc+hhqG0ltzEBJ6PvcuoCGeK9GsbBEeH+C
IHCeqXo4mUKwSV4q8a2sklBNn+2eyKbu3SFPCQpQAnKH0IRnD/a7AsMG/k7E/Efff6+q18c7Pqo/
6RVQFzbUSjd77cBI5Eu3smEe14/hXRryPxLtcJy0f75Vr7iat5NOJzYNmI2uWaptJuYPAgL98WDA
BQumIFvovD8KIVoLWVNZxLSkjBl8XqvSDrKvf6wSIGArLTiOelnvt/2I9AFgPRKfPqsNbhhhrFgQ
sRWdB69cLUZY56oGqqux1Dr9V/RQ+0mINCpKaUAXntSjtYOCGvwANDLy4Le9F8siNTLc0fUWpYCu
uW5lz2+NA1XtvfvwWa2JJtuE6ggNOKdPBDD+GnB5ceh/JuVcCR7gTlLmF5HqwNRkOqAOqtU9Tu6C
t0GCl/0NKWFYGHoKABOlR9oCvTpJgNkOp5kf0KO3wH+L+P4PVMLaj9X9c4k4+1bhh5VnLlOeXpaZ
1gLzZ9ieJqAFfDQ63hDQNgVx7IweGu+S4fagkkAsjPQEMueGYW4yIojWkg5dEOyYr1cwumyZcjEE
HWVaXoUX8lp9Zfv1SVraa1m5lW10h1MkZ8XlSeQrRfikipyzVkli4CiPZn+3jZnvidVuQsD4nssc
KZ/jsRJROz7SGGafrnTrZ5ClJgd8Y4PG70KuvvaBHTt2Yaaa58enIvpxUi2rgwO20qwDstiCz8py
rt7gyK1Fp8PS2lMLad//U+45gsXPyRvuuAasI0qV8BCbnJhPRqpxDaIXIXn211Hr2+1NB63dS2Zs
B8tTlrv8I4GWV7BJcanYH9cGzVYGNn/fBP2I96Qf74dXG9/cFeJv9Mxg+iFNslTV2vczlDdBB0GD
k8wP3E9OqSlFMM8N1udDFMnqavuQgZRCNoAmPD4I2OMiDUZd51Pldb/1vys4HdOSjusp+eq9VkKh
CSWwsQJVGOYawvX7hcmCK9Bf/cTBjDanqshWEPhpkjaTmFyaRMn7Z3i7MYEmEYjVlW4GGElfSJ/j
dojq/OJCxiYLxASjCW7HdyUHZswJ7E7eWVl0VIHcHzkgbBqKv47fEHC8qSEzGkjLcftXJKdYwMfG
21DaeJJRYXSG1mZyNnanGsxeOBwbclG/6YjbKwKnOG/WwU8KRNLpt2M8J+xgwS2QWfH0s/VqQLGk
pc5lHqZlo1Z5BgTDpbcPU6hF+HJE5NgvL/R2Ov8YUNPS5BjIfI82nbb0NUOGSztZ64CZ5F2ipIPZ
cINTDgNTv/va0gFUSBigk95aBwhxZrfZ7jYlx6QoerIEgXkJwLLMPafA4Fjjc2iT3vbDzdEkxS5D
6QCNJ1dbDeweO/nWtqP3xHcX/Iip/rHk+yRlSo3XXl8Gg+ECsl4uIE6yvnVmxwPAFPnaqnZMZSiw
4osGcj+sle0jsbPf19+XScM5tSEitq4vieCw6BOQn7VcDsgak7viQBiraKHMaTVsPTc9KNbf/lQK
7CanJ0UxXZagbPKxeVF5XZw7mvi/54K2iB+xHmtuAUtT44b+5zmfkaJ1Z+nuy+miuasFgH+JLzF+
DD27YdBeFDllfP/27bz+I8fvcf3DHaeA5TehEAF/Ul0USK0x/st+eRDNfOFmHGvrVypHIttAIns7
5WtJeQCGwvRzkYJf0SYWpVxLMuJUEw5i/D9VAKXGSc+xnklOdkNoXxyY4U9/FoutHGzEn8Xi95ZG
vo4eojJ6jWAFowws+F3yr9kzvmaAImVXS97/Eo8wmPD6LePfJF07/5loU4/rWs48R2eFvlcataM+
0lo10a0EwPglPP8K2SbdkYiHnbz86ephW75V1Ei3dg6MNaeBpMspkiYkyrDC09EMYuFd54WsPqtX
UQP6TOWANcHjCa+agFwZVH8TbCuj4H9ueF+u2u67z1KyD7thMLfVlda+wSACRENjmSuMKBh014Ba
jtQkCiAtxtDcty3+esya/1YaavXDy9rqh+vLWvYUa2RYf6L2lBshwM1Y6tRzurn7WMcUet9zWjNg
Zy2RgOVjYWkwuwxgvftXg+7OdYeAFO1LSFxea3baCx5hXNhaCyLFtAG2eHCZVjezxsmUk52ZeL0B
XY+nk9sSzk1wECwyyCWpgnOWqvcJmXmVQoScyU3QckrRV73n7or80zSZbezoIIzUQ65kNPaNu9+v
VyJ/FV62mRATTiLh2Q91w/glXuUtIL6xoETQW9RHFTt8/u4+ri67hRp3A6+EI9nWYJLniSe0NaK6
V78phSjDvkKfTcdTORpcaIxWnNp/DGdvAq3aQS2xda4bbjL1hS6bxFjZKPNSYFQWIAqbgaekVsuz
Oh7vOhMks13fsWEu7RoFAVQOUeuWBkVatBxn44yHkJCCJdjo2+ARzP5ngxgUIM3BnLNN6U+P79zF
LDRPsE8bFAtXgjtfCW9wwS4hNAszKrEGWzWUNI68Q9RqiKoo0od/xLt9xeZlCLyyZodSv1ce4bjc
YIzbGRRN+6L4WlSeJa7axem1q5LERopIubz4NJmT39AHZDjlB/cb3E6Bhtotyi35mTf8hzywMWnT
HUfoWEmwDqXsd2DQ5dnAgAHV6GBjQJT3tyggAN3MDWysu2pqdUc/C0QBRM29wlGulQLt1ROSwXmZ
adPx09Y8OXl5moywunpnMxoMDEp0JjKdjC371zeEjgEm7udAk9vFhYGi6zx2Q6tLHLeRokxhwAT9
P9xy2fDBKPDHwbapY+UkZZvRCVgkqr4XVb0ytu+8NXHOOFk0qv0AJpJCoCXxEyc6wDZonz9KlaT0
ghtaoZx7wOl4ZIx39s2iI2fgv6KUiEucDXf/OLYZpUE8B6LS2GcyOXm3NdVMqeTYuz2RjNbloiRe
+9K1KJ3cLx3cdqZwuc029M/6wI4ixAvWVgJ6fb9DgShku1EskYIM6KH866JWuMmxbCCSH4bcpKjX
ltbEeS8OGmh4STQUheKw56cwXH4QX006Zf8A0f2O/89AOO7w+tx2rZi6v86s/Yl97fc7Fk0nVmBw
aInnTWDP0+232HfrmjF0RKPOFCIC8ch6VZTCI5CzRTSc8rn3d3uw9a2hGiWH/YGnktgwRb5bp2as
2kzf24Qjg8P35NW95jnQLn2fMjkjMegnMvF1EXZ4T2j4NlJFdmPY2OsKfemuzMvpax4kqwR7HVFo
KGWLQzYy/Sh786kiT0XO2fV7QPlGMJKfRCec3uSrwurvs1p3JtJFf9fPgN8qnQFFOTrkgFpO0p83
wlj0Hs/iT7N53TH1SamPksBXCm81aZuHQ8Ho+LkfnHncwh8fFHKVJ6Ip4vb7HKhObzZwPTPcIIwn
6NdUobmJvlwx9qrR7gdVUqwsi3g1yyxN/IiJHX6qIgK8Qfm+s7PKXVgPfkGJuK40noljoZpjQF1B
hJQpNYa84C6ErNrOtJXtaOb6nZfmdN7drPRpkG6ueewuQr9XLWOTnMAUKkGDAgQ8G3Wvb0r6a8eL
3l7fQECbMW7woVAGICRhbtfoSoV3XqQfKuFGzhdoTgwvZjbDOsG8WAqUc0QbWM3+SEKZrrTghu7y
YB7/1dD/aGTBSfWuwQuQxcPkY72oY1oMD5cAnC+mKojX012Da42JG6DoKjK2EzW7elLWDDMHT1Sr
7et6Z983fCyB4ir7PYqSyc5sVo6o7Pxlawc5d5vhioRexY6G+6tSRhtJ6VVqyq5W3imBKg9c2VV8
gK7U1wLkoXTlnwJ7EpWWeLMWjOKvInr8qADx7OHATkOYIrMyzHJJZu5sRQ6e9JyhYAYrziJ8M+yj
WJuGJsHUJpkQjEXD3OHmuj55nBjuirpplfNDjTv1JloJbAe+rmGLKqm4n3Osf0BmZtqPw2lC5pTK
1tyYTeNTidhoWZ8Vs8N3iAEzyTAwc0hDPyZPN1chGNB5Yz+SbBPPUGRndbS3FbeYeCXLWd59FLJC
D2vSk2q5BFxQNbw3LUBPGi2gC5I3R9HoCvAy7pXD/J2EO4BsbgS7KOs8b6TJx2pMBrdEncL0bxLY
j+E8hnZpWHyEu9i1PNcyp+LmXxW8nB5aiGlfnf9/t96jU7MpdWYlUaLYoh0EjKqhjjF8kBTrL5RY
6HNb8KFfz/gKPjv/Fu4GEvOaZxEzgd+iZ8jW2IS/lGuwiLx3AYvCwvKQF2hDW2HkXbOBrvvkuL7q
G9O2YXoCgnqhEya2FZ+lUrobVvn/VUUCemAI02fRmaed/2Am0oazLsFd8++C8h0t/BZbaOlk4q8a
pcgOaf2dYWZj6MEwIlvExhjzhJy637j9sSiYgQOxdrbC+jpFMMsRT+vSRC8ioO1ZNngFROxqkaBo
Li39w6XKCaUv1r0qZfXROvCw8wagTMVxdoyqlCFbRC+4NpvlYR1GBfP1Dw6Q1kT9O6N37GJSi0AL
rDfSybgJ33LCYcf2ChpwrLLWUbE2QbUjt3u+cF0swalEoFIig0mCfM+lJT1gcy376pNM1M9wjy8m
4IqGE/S4wQwFumZhdfBC1lbKeCT9EW6SMDEYWxCHt1xUPeSUg3KaLoMFCjieY8aVzogeSGxrkjZy
xIuQnLsF7oDsAKdcLYWBcPSQhcblUtf96XaS1j/6kM6KJ0T9hGlRltAmEd0o8WnFFxuC7lQ+Z5jv
NGQ0alEO4ZurLNx57JK7rZa7cboeqKcz6v6f3Vjdxg8gw64jbkUjuUnKn3LLGQH+PMCSlNAUKl0E
9O/wGuvmmzBJi+6BjVpgoRY+SPCPXbtjbctoYE02fziNZtno5c+Shph+BbhD3n+T4bFKzjfVa1xD
KXVZyNI4UnPEG0keB7H7ujixOEnA8TWWTBjuKaffaXRXZxeNe6ERo3XWs67LIuKwngT25vLhHoH9
v+WBk7nyloLJtOclQk0ABYek+O2fqu0w3zKUhsLp7bM662iy77GypwgqDzt+k+36HWy1f88F2Yqz
iX0m1L1wv4v3LbgrYEwfj/9IRNDM924FL26NrymgcCd1AsrgNqrT4DrEVP5FEDoo2cqDYZxd1vL3
YvuPJ8HPW7CWhVnLfZsCvenBte9aEzMGb7wzgBSnMmvr2uoEvYQgWHAuhCVVuJfmcU9jHc8y4Fvy
O2yGJoShVEEA7+WKpQQvTf7i7thZXrfS5Cqt/6oHgBUlroXom407vB/kqUvliV1vubfySbUeRScP
jeM6qUjbCumwhzx5tbsz5Hr0pnBOuA4GEl5/zK2CvWvMrQvorj2vi/z3Nzf8+v5/wC92+ffpIds3
2qqEWW8hZh5RNHf1bcEMOG12vzbvnegiVa7LZynJd8osEY9S6c3dcgfgGIRy69XeJLLTaS0ddn0c
bv88VJ+5lELj3xaGn6uuwQ0Hx2hkQWn81BZh2mRxcmq9DAgOhTcK1gHsFoTLd0J6J2QtEXqUiVeY
0iyZ7/x0UtDgklL9sGDEEi/YFp3zNUukZYVBc61hdZOaTsfgGJD8LyzMC1oA3EE+quz6t+bFDhUG
PP4sYPpkCxETPYmnvy9lpYPXounBu0PuhpJ1C0NBvTO8pNUuElZE/tBMYHRlVaREmtvVwLJyss8/
Dk4sYd7QVDjc4dU0ZHb0xFULQ62F1+i1QvYSHcO+tc5gtnDOiQkeR3eZV7nv5TGKqlvHCRckg1s9
t8Lp1MgIbb06Bz/H0KmkcAX2Ibip6TZSZ384iL4jrapLzhDSes2noKO0C2ix7sU92bASrgL07AAa
1xQzbdgy2xj8vLzrLJWT+ENGSjpvNazeZX588yEE9X9VlijvjtNFNvC6sdW1rBdYHu0undvmE+Es
NqDFyfPrx7ICbUHKRGxUCQNSIZcIHiLE4iIcS72CO0k9zDmCISUyB6urkXhNbTyFK831bjrhAwSQ
DhEk3oELuVvfd8p/+EEzlon8hFpQCF3uMm6OEdoyRTVtstO2T4MGJ0yKnwZF1nJnEDGCcSywpMXt
7NgSB9Wxt/Dz96ytMxutVetl249NoaUGjpU6xHuBKwvmCspb9tp7PxIAWGgJi1ZurXUa6dToYF9D
oe0pfJdNutTqGVdwd6psTGqcjEqk7YuBG0RVgNej8bRFJgbXw7Nhv/INCgtyb6xY5czkhSj7QXBS
alv3zWeucvpIi2iRdLOv1P36HqkI9+Cdtzeqyb8PtgZB309NRj1huK1CSHJwYPEyQYTkFmaNU0N5
oR6aNsSyRCRTOKI2POYNhS+xXK8qGEZw9sbeB+JVLfuIpuX5ausXM9apvMTB6oYMhNdHKW9OiFxr
/h9MgWFh11mY0ACNPwUyVpvPox6eQstxxMigbHTJl/kbfq2gULvbB8GzBjo1RmwNDs/1nnm0y3Rp
dhkgR9/bd+e7qAIiU4BgTQeFJwD4zsxmXLvcuY0VDsYVQ7EhDTUtiiq5JY3VqbnNKW95hpXZMuf6
opnrhCw/P2GdkZ01XO6tKYKIzbrA2lJr/1CcyRBxfxKFBboUb6G/NLZQfmriE5wlj4p3gxMhKwlY
+9qskVplY6p/f939R3Z+AbKeY6TOtmOflxpy5MirHyAOzWchNgJrb4dlo1O2piFdS31R7jtp5P+9
7SlTjg9+fv25vuX2Xw+HBipGHxtWS6pMDVdqvsCOQ+0KhTYJV+RrFCFLtxipCkfoQFRxQXK7Z3KR
slBJzuC1SEKZ93bL82lvSHNB1O0cXrwDXd0tfKEne7XkbX5V37su0un9TK+WxglE8vDIceWAWQf3
zKMYO653SCBNtJxZ84gKXssdIIH2l/Iql3yo7bxGLrjOFhxxE9lMdOxl/3Q46uzXH4aCaeRC2Gjg
UkaToblJKyuen6Fs7VkkteGs9gsiQt5yPfGU8yZ2+G1HwyOOuhixYiNwLCqg6pobC+EBJOtik8ax
euIUHsvq0sDERLWYswSmJP33Hlbj29QHDODXbih2MDA19dO3Wyc4VJk2LJwj3lG47DWzgk9XPgen
2v/Ch00ycpIr/xlsXIPJYhsCkENt/8K5Kfw+bYdJS51u55ibno6VEbAjvVDelH7VtcVeAU1d5+UK
zqBZiJ8M7ykMBMSq1ElQZWuZqFsHB2g//nismU0coJdEj07xMF6mRAoNCvg/6F9PO+tRPFVhf8+W
WfxHy/3PUAOw0cQNKnuVjI865H071BKRP7Ov0GJuNvPMaXP7o0EYn5Y3nDCDBMYJVYfZOkX/F4e1
z+wRPquYngLzu4JbLNlaHYL/90uXchC0R4MnjmDQL35ZbyZxZ/Xs91IxHr1OTCpPP1QFlBu2Jofx
LgB9X3MXenB4ueCph2YF3sOsBpkaTPBb103U1D2Ccz18PtclZyj4IdalPvUkVF2s0HE5JVyrOkdp
ExcxweaFzMmYGDFxbe9DxPaM+ujBpETujh+a/usyl2/elulbyS3CXw87CDAyDMlue/2wLVqNtpK1
KGsehN5batPjrl0zzzXKBDLOXswBE8Gc8leOp/eKhn7nujCwcN5DiNWwC9Mydwi9alsGg+33mW+C
/J798Ea3gWvkzYakqjxOESFY60MlmjF6o7O6VSNWgeMe4fmXMg/n4xi0cocbime8MDAbIa8oZhGW
tQee4nrpUEwOZrVNSujz82AKMJv/qWgIFVIaWxSt0WWe55UPE8CuwY3oqcR2DxQsVrPdLsBp0TZs
zKo9GfmUL16F+gluLoX7Gj2ergRYz5PuB4h9vrtt3SrlndSYGgF0Ghw/jm+mAGJUIX1l7HMHaTvA
SlIeP8N8hLVzEjP3KOjDaGm0DDn+II1/JMTm6/V7jg1zoKwe6vtKsi4sA5NbpFDlWy4uvakRP4KU
KXM60Kr/ROlu3nTqNJfizu6RKknez5Lkn4xWfq89238MXDlSalzI/g6aFbTv7QhDp1ANio90qxGm
qz89r0deOQimqUQ7fxZcpWZuNUyHFqTnA59UMfxndO6t8r962yjiZJR0QiYcozfc9gWrR2RTIv/X
9MGFcySb6345N1vrb73fnmEV5RkJ2nAe3awqs2gKX3+FP+BEsky33fu+PJRawA8GymqMaC80wfyB
SsRtLADUS+TXqcoe5uWd62NEhSEQFtAPe6omIKroSp2q/RppulstnfDuQ7RC7pBtSmILbmorXvl/
sTv5VwCueW55vvuv+54JaG3xUVyeCp7vuIUxATCdKMfozDDGw1nxO7vk329cSP6NE3JIzqaJg8Ad
6StvUEVJAi8h+2swxapDztN1EiQE4YP+UIBRcIfobO5elPdCHQ12+XZ8la4JXbDihx99w3eGRVZ0
VhsTL+N9zCmN/4z+S4sopa9g1NmRRDdBJ+vpOpWa8i4s6a6HMkHp7W5wW8pyIehaoEa14Xb08bNA
GDyB8b2ICjBHKx1Z0+MzqKAzK0kXxBgt7WMPX+ojwknInIqc9bb31BVy1y4F3I2kbv1TqWtMRbHA
FeXh1M9neyuNtmOQjF/vAIz0yvcEc/zh1k2kN/rO/BVuApTg5WEvUIuKgMa2ngZLl5tAWqJs/Tum
c+Sebij/phcwyXfcrsIWdFjyj0S5FgBbdX68pFL4YcDQf20SshUPwxyeD4wuTNKbtwSaCmqJdeke
caBNnatOkXIxBRnPQEvIj1WrTgyFZ1iyVcGasX1to4ugp3YoIjV0VchxnnIzP7ZEwc/GDFnElhrC
eWZqVPngzeCKkgvQHaASpJyumJHEzOI3sF9AgpWZxdvgi9XN3F0o2N/gDWAAJ9J00y17xCpD+pJu
abCyl4sT+3DzsupdAuolohxoCJsqARx3JgnoeIfm0nRkPSied163b0dVrKDkF0cOAiDInaaVUKKP
MnDGYAaSQkh0MlEaLIbr4zYKL2eAiH6uNoCQabnJ+Tlc78+a95fsnO7ox+cOUW1wBq6I7b1bdE2d
ZZdGoWrctOuV9bYK6Ubo6VG21SqAvEcQCbC5BG1tORXpZN9Q5J7X5/hV8UVloGYTgMvcbh0OIDDM
yvFbuMCr7q6sWiEd3u+DC+AaZSpISBO/JEE+Byb2DBJ96KeylfQdDfs0wUZmiZr26AXPHABX5N1c
0911cmtzV7UHEz/W3pQHMI30jD1T7YtxQ1DPmVpCREn8mrWjt/PQByawd5MTU1FeRvzSGmgw9n5s
J1R/g5demXsiYGtRgJr4mJLeIxfuJ0gMvTHb/EYjOqrvnOWRPDPdXD59kCwkmi0iPKC5OgKXGBgU
WxbDwcYKgRp5jzkDG4ptIIpGWOmtFbAPMz7tdpml61sIAQv4tOiR3lMPzCTfl9MkuZMvrnXTdeXy
+1ORHHe3ol9ZO8i7FnsmHANMNcxkV6Lbr/ezVXSakLhfBJ5hbqVW6QflDmbsUEeVwEozm5sQQPxC
nSESDkcA5vzLA4BCFy317mLSFoIkDlCeM0f3qt0Ohj7PY/zXbSwLJPMVnC/DHWGl86QpSY60pGR5
84ok9uWKjXVdSdDfRFR8bEi7aai7sfltPqxoQsxJyu8+P/LHlOzEJC0/LHnT0nlapriLN8CTTj1Y
vU3TyN9RG57CUebcFpWkWg0kfbfRM3612HcnqD9XFralqjMdbUEzUZTWnIbL60ns+TIKTRTnki9i
Q5LGhc1G9JY+4SEwE2OsNOzzVuJmjrpq6JPVlX39rRhwqQ70L4yl5b6q5OoJ/1XS6w37MV3usfC/
KC8Se6IQnO9QtxZfv3A4zT9JKmLCDhguElKMcgNcfFys5YMf3g9i3vi9o3Ys03jIgMCANhITavKD
l2UduWOwDmUQTJ0Veu7BnDPb0YmA8IjcDQvGLt5V7EDJdR5kQ5I++Fk2mruTUvskhJXseRKd5OC+
YCzmi5N2oMMymRMczFbD55ZLEprjribn7J34EwDjXAafdD6p8E4n27WATmggkaYV5ZMGftaEihgl
2w0uV54W0MgJUA7ZiZp+QkFZcjKZeefLbJEv5N9Y+TaCEYEgvi9bSre0+foxV+Nu3jVfIsyIZTV6
EqDnBz9wDNNVzRBwrnpE6WhK6t6raDnj9ykNpXG6O7iSxr6sBkMcZcfIc5YLkQqcR/cq1wEGi3jj
neMy5TNbkxXQ/rNZ+meCrEou7Nb3ypj6Kcjp1yojbr1i+YMItTaY4oFgh7eZCALc4GwK5DT+X71o
i7I6m0XOYsgIBhtQMDCglRQ6h26VRg10tqdqMGDaT7pr5uAvQ4P22mkB2KKSAzZE45FCZECVAh6g
iSffWi54xcvX67bKJYdQN7qaxp22Pwtlh13wrhhvoNjBP6ALD055kJhAjiq3L/XqSCJc0IrdEBUc
vB6rI1Ow4ZOAz2bOoQU3+3w10FksAJAAvXP4S8rhJRNpd9zINoCfsN3WS5298ZqHkkCOnnkqUXUA
I7o3vK0Tr0WJSWRa2KOkmI/3W94iJUWMkFCcMAwauCtAPM2YouuFBBs4EkdriyTVwPl8Dd2g5IMy
Mq/tXr+UkJKslEC5obuG8DVvZPIZE+vJMFszz+NFhYON1sNeSPi6vKigNPTgaSuz2h5FViajwBLN
ItYXa7DgvGAXWshqSuP/zGYPGBYt+PkYwd+rksyivZVhacDVZeqIVCb/+jOljyahBaaNTZnxEbUb
4/0plSngkCtzEEgEBLeTInM+vyQnER7kdbDDSgnfd7fvClGPkKbNmW/zFeCuOig7ZIlFwq0Ohjwb
NMHazEk6qd5QmCCvtx8SDwTSdxTFM//ouy/JHB459WVyu5xGraPHxMfhBsfdBABqI4yboudMdIQg
zegBjhHx2Fm58sToWR2HUhfsFmtv8jILd/wvmyXIeNNuS9nBxp/ioRgwA8cNs5+NGmwS1ak8r2Zw
wM4+5pnYylKtkD3v1/ugF6CciucE3AsTQS3FEjl3uhCterudWvHaq3bkc/jvjjWHdrUPcKIS1PFl
rSYCXKMdqRl/rt7H3KfBVrJRkOyKfLeahuDUd+lDlw2YMh0DZV2u8S7gdJWEpm1OqO4wDRMvmHaG
qL1KQk6zlY8/rNdiPJoGukJf87f6N4XqwSmK+MTD3xsmVo08xXTISA8dOJCQHCjgQyJLZPX7nVkd
9WXmTLpaUSc22tpx/a5+MLbbseYs7xknpQQ1DbwTyFnMukErhcPtVSkqA5rEMDuuVNJHMP26ZhRX
ahHxWEQEjuOdEfva4sDcm9Nepr3TOAjUxDxqk7Z2/8BIMJZRKrJiEhaN9Ff93EUeF+DVNzlfkUux
TfDfIZRCJc0TTASG9j1cxPXE58u1Pywe5NWaViqGTAPchcaV18C7rr7p553hXrIUWcW1vDBfljyD
e7Wd4AYk61/lf8jaPRbgVfLyhC0je3QX5fhBmgv72gZUXHEIJxFhEdUk8RahnDPwtcRefJh5uhB9
ZjX9j5DYLpxh+XyyxoGOKEbfV/neXizY7CMsDii880rdychT5xzrNZg58FT43EfHixbEZZnBY4ko
8ktf9Q6kxWKq5QmaZYJ0k4eugUHXy1P4BQyuBTnkxiM4H0+1MvWtjDe+um3VeaghLZoo8ux8G86f
kZEKQCNprvKnQfo15ongscEvG2usuq19nEvCxCfrS7rXj5jyV3A+OL7lFV1I8vwxfeUo5vFYbut1
OIjLAJhgtnTi798F0nNCbRZ/nEqqvfmDsF2gfQwYNvE6l65vhhX+oOvTlGGkSoGx5SkZ6EEzQV1z
++iAW1x3nLropm0JFfD5VMHBClrbkvDlWylE/PP+5ksKa/RMGrif+6k6H+UdQK0wLe4P94ss5Kor
2iarf7TLa39/O1utwcZWorTRlkA/EFsZ9ETJV4W+R7240qqXpFiLUmMD+AN9MHnlJk1ZDOdmyrg/
bi8WPV5bIw+IYhOs2WCoPNSSGBgf1f7ukMow5D/RpHYbM0KsCr5yw21dHcioWhVXbnJlClyau7yA
dvV98m2HoEbNCyCTdpG45BWc/hwVdb+XM28ICzi4RDCpwGjElURhV+eTIQdGYcfa6675mdys+f8/
rN2OSwCMeKbWekNN38STPpZLXDCIfgdt94f67Sva45UoDEBopMCPkV03/pwazk6FnANu2jcK8oXz
OJvCYzVtQKnU+HCCTvj2yWeStihG7nv4wKQ/knLm3NtumyKhk6rIJ9ihf0tKmF6FNcX6txgpRdGS
Lr91TJdWvsjqS0M0shwgaZqZoD1gtEolWeDwhwjK9ykFh2ACN7vsc106J4v7McgYuTtYeWylM29T
xxfgS9KN6vbKpu6eIhxuNOpsMt9c/+iMUXFZlCkK+jfkXnCRtckJHNScY/d/ZF7z99oB4Xac1Zjt
/0pOveqnRlFYEwcYt9Iq2pgYkHRTa+KtCxqk6Kuf8zGVyrQc+hWeNJEoAQLX8dq65zFuyp684AFD
q7bCoFR2kXiPWD4kN3HFtQzAE9QLT86YbDoxIUXuJDnfZi9soDKhTa5CPbvOlevEhk9yi8PUiYlO
Zy2NOUJrbUA8S4vW9qAAxbcfBSRbkA2RQL02oIflgRsKaveAcYe/kUleRB2Ux59j3+EVT/CCiuIP
kQxcd/FlLTcnglyz2mUl6/E/dYQ8G9hN/GvZzpSzvMOa5q8s7cD9Jb3WvyEqIoVj2bB4Ib/Q6VtV
OwYb7KCVtzV8sunZz+C7O5AsAJEQliYucHOE7twM7+YqgDqWqbmZN74fXd3UE04a6IDLYbhwdasl
U2UHWJKar074AXCMGuFX94EnS4GcKRgWINnmzOo4hTm4r0+i6nn3W1EV6F5NP7hMgoibswUYnqHK
pFg+J8gVFadKhVfMwKxKC/Hy+HmKbR3/iIwlyjhJQIs72K8Lk9dJbSzcBe7nzNtO68VyKSN5fyRf
+BTK41E4EMMQWGWbS/E2UhYzlBqalgkTl9KElolWWApyUl/TuKDz+O8h2OSRLo9GXLzC6awFl3ZS
DzEIlrRHUQz+odACjhu6MkU4YELp81JBKzR7fIscGJ8RnqLZAQ5OVl4WILbSnAP/aA/dytzj4BSa
MErY7KGa4rrY2JqgWMUTGJPBQ9O7jDxbFc+sA1ytee2cHcfF8LgzuQ0lf/Y2VXVqWVRtTbQlGiRn
MUOOjRr6NLvQAx/MREeXoWm696n1gZsOPJkLB6jkkY2ISstXiHPkE9dR3Or9PKznShzLPFz80GUJ
mHD5sIUA4MN4RgmhPrG/uidyZY5bu+NYBlsOepMnys7uFlf2Q8kHIy+dPFEc6xJtoRXZqswpVls9
WefuVNarFSfHJ5aSI5CBdgFYIHutQizZbLZgYJn7NYEjyK4g2yuOHUlokzCoWLfPAnaSGMlnd3hR
DuPOmYCl5ZCdkcOKEyPKFIMkEapV0blpoR2UcyCLORryfsNl0TvZdLOSfk53BD3CWZvOm13jqKQa
fEGGrf6072IKZkwiPSDk5BSjEZbHfCWe4vP5H6+09EpnIZMCe2NFsaMDRyMzOIMeT/hfZbskWDy2
H+7OM02hTkbOGP7m+HisQJYdUcA9fhtfPt0EmXz+J737noe1pjTpjgZi3Ikrp+7aDuAiyRH4XaCe
/tMipvOuO1UJ0krJ5elkLYmsX8Ic0FNU/EaC9HXsuh1psMPZScg/SWbPDSIA1n+Nn1tycxLtaMOp
JcNsqzYdS5jaPTfuMfjp4iBFMiFQgK9GZyOsgaJq9zxkVOT4oTZC01qeW9FpHpq7zjQ8NuwuL9DK
MuB2OP7xmznB0KOf5KiLr2lnD7lOkw8wL5ay6hml+S+51uQNRVbp/2u6ysbot2GGAKLLed5Y9STo
1nDf/yadzJOBU3+xeAq3SczoxIc5pNT8Xc8UGA12I1eVAM1HVrPfPGsVN5qlnc/afv5tSqyQGrNI
VzOjWBkD6faGo/0rNVvOqlQhWZQsIxTMdyQ+ezoxQbobi7aut6yhEv84ENib+6DBhSEOQHeTME5g
mSZ0sXASVWJ6NIDh/LTmU02WX00wT6Ln7XmixB2i1V6eu9nlTIVo+b4PPyZ9ziMD6XtfqS/2giX+
WoLXMZIqwh3nJFIY2dlZ5sGWx9goV0o0Y0STAYUc6J5RlOcA9wuXypNnapWHzN/q4xQDzB4XpgdM
xG9ezOY8BIcvgtKOzKLpTXTAQ/DQgoa3JTdYg5cX30e7f6hdYJ3qMNndP0pcE2qQhodmwNWXwaTe
bUhS4wKGe+wbV+thKGCNXtMn/Tk1aaboFpZiiYzWFIp/jl2TDFbghP0GSAEbB+e7GwjlTyyZHlEk
qceTvJ0c/16QsRV+T+IRGFIJxFehlFgkp7ihKw/FJUXtPAl2LTJ8rKltcG33RuPm/Dkh4luIEazZ
66JJ+9gb/qTY9Z3GReJfsdFwzOkr40AY60GyM1xYNPD/w367qeLGKoLpllt8tXnsV+yVd0uvLxtA
xa+eKZrPDBl8Nyo9w2m4WYmFWns0qZQXsIBxanEehPUsTupIFeE0eevCO7ZFQp1zNZMgKlCexVfr
Vo3m4L0dezNBiSxR4Ne/OtC/EN9T1FFxtixu+7j04jZsgaYQZHovJaykVzyIpvQYW8HDgbi4GoOi
S1YNQPeO6TDHhZacVZBUgHcm8Xvvb0rEjzH3YZvPt3TT7a8HLXXPjiNa4DRWP4C2nLjvu6pUnKUD
iOt9vf368ww3/oQ1hgMNf/yEIkToA3d6+3vnZnSCynUurdl04d4fSkuCqNViGG/YsIjVcU/Z20Li
Y+6z5gtaOjUlz0KdfxfjWB5MsZPEs3rh9m7gHS74AYBCs604DKs4GgW8GpfE9kd7aIWR8NMhRcgg
sQ2QgRbLDXRix5uiQT5BmQbJwUEMoLjO8Xl2hK9yd1w6VDYPYh6T6CixAeI7V6WsLwPqWJPs8OP3
5ddQRNHufQovuJqQv58QL4JD8dm38q8W4wmE0JnpmjXaaSt63ORZnMOM0yWMkT8pBBFySnDXDMMn
hccFoJDjoBjUd2nUE9NyPjtysqsi9UpDdPU0KjDatiwLx8XDp6IkEB5PXk5yBKH7+jSSEERYH3P/
Bpbvj653S1Uws5QVyl8oMIw4yZYRboH+dqBe01/zWuEznFsqucvi7wKJW3BFFyk15A5HMfDtoYGc
oZHkf3J0jtMnc2Vjl4ReFoKq3merqlixmDNPZIiFQXQQQSSSeBmcBzwNoqx06SA3IKQPsYyu4nGI
FO5myDrnpPr5iHayay+IRUl8ohWujYBnzLef5H5sGCa6ZLa/fF0MMjSBXiRT597Mp3dHBnLuPPu7
IfJVfti40+s2lYzm2eTwpd4k2I6OzgGqA++J9bqiGOml0PuMRIq/mOi/ffq+275vKJGu5UM8Yw3+
0I2G7cf+zVJGu8BsIsDFA1ChtQ+HCHH8lapAaGg+Y9qfyZfuuD/lP0WNZKuCpZ7hPEMbRA186okT
xJlFQur9n43hCBPQ7FU3GvbF/NC3wcO3tF6RZVXdQwia1fC8JbSoxsQktGD3ZqdHb45AxNiBL5g9
E4dlH7vl36/iJqVoRqY8trgMM51tAxND1/ZA4z816TlebjY8hguk/bS4enfKG82v1hJRjbMIeygy
bI7VxkaeA/ClRTZTKiWMTTqV+uJyoUIJ3Vs9yLiGle6/MS71MztCTs8LI5UY1sji1sb4QXlR/wQE
cM1i+r6BZKuoLHTaw5e+r8l586wi66W/SWB8mvYGhQqHXpCAjpgvmrywIA9QtVXK+ZfZtjSvdnJj
bqhy5fIWW5r12KmquK2nkQrCP0OC1L7Nr9FCx9qLNG2l4Ws1xAgGmHoca3r5Iu/c4+5ZgzywWYfY
g4sVn3z0RPgv4lZqtuuNYuxghLzG3zr8JpipGP5c5MzhPa3WHKvL6KyKdlAI4+AbSpDw6g8thXun
JjrgxTSDlVY/8G2d+M2wtBP2WzRRLkoVAnK/oc8ajRPdc8vb54iftecEXOZSaxikCf+tBMsmZfoO
I9inoaXiG7ubire+wSoO8XPcouDspnZ55SQab8orcV0p2+Xgtj1lWOXyr9xBYIl/i9SalUxnckpw
4StVlIParRlLrUGiQVaH6OuT75usGazT/Nzni/pcznFlwAm8qcJcyPmQMuFqK2+k4uYzV4x+YZyk
f0bEeQHGdlt1kR/e0KVI7TLXKUpM4pCkkKV4Q4tIt1VVAZZmPnZhpxnumnTEAuiwPqQg1AkxChCi
Hn9dREi0Ady32pEcTsPa0PdCa8Su3/lXI1OXk3vuh2oXe5EsIIH2BAklHPDw0U2kaQcfi8HdQPAZ
8NlvrBcCtATXVRs+SQLHtw2Q/xmyp1EH7OM23xtZHlkVhsxf/CfmKbMUA6TSrJ9CVT1SnQElhotf
CofPouDcQ1rVzysR9fGsqV9cF55OQ2nB37n0M9UY+kWCspSExpK2dgRXPD89hHWPpGD6opNBG4NS
C+7egoDKqTJH2/ylH8I2OYgX6RBRH29QMIZu0XMrk2iexR0DwQ6w4hndFzG+zZocxBnW5ThWmeS5
Ld4hNsH7bb+DsRbvc1/BRe6btgnPr/KiaOtuy0zLT7hkNTtY/dBoFoxHDx8yMUekcrmZdExbVJze
GplgUVbxielQ1cBBCyI+SWndH8e+mRRkSUcX6Aq7vv/EewXmAE8N2C4NRuyXVpHsVN2KpSEfeZu4
SHX15IbDjKCAk9Kq31JuMWNGpHSpZEaemi7WoLJxNaNlhWcUJEHQnEjSUIlohaVujsbOV73n28pQ
INLpjQusPfIcgdV1FF5uEt7W3rjiMecTxubZ5/vhiaYenM7/bxz3P2pKAFvEimRDh63Mhws9xCNM
C6Zd4vf1l0zdjPuhapFACg9l+iSASlhQF2xLzipvBuE3yiKMbOSUjHTmTSAfyDTcrDL+kskb8lOY
U8f5CHs8Kg3dBQXeXL0uOJTwOBfIYsAShWHGPQVCgGZyGQWL+dLm1i+e5tI0Q0qQ2ZPOP3fUGEg8
ZNKEiA6sB7kyCyJMG06YLSZ/TSqELQkx6uGUQ7RnOe7QFyTI8rV9pozo+TGMoeR16p9waB5hClnm
dz3/fxNXHGNEpRlsKo5eA41Atv6W3sJkBvQNgo5/qinaoz20KMgzL5Sss9T5DEUNmGBlYQNElgzX
jlKpTbh+DlcVuhiuECuC7EK1PTWgh4/OT7MxRFj86mm7vU16fyRH8MeGbPdEEiLvAnLQF8IGqxYI
cH66WkB3jc9p/ebjArQSy3zkwRq7OKcQWS8YgdhSjt81OSJ8nzqYzlcOCN14eKHj1k5IvAZZR6QA
qNO0j+D7zFGqU2o4ln9J/2hlN0+9cm5CKL6u6Xv1PaD5Og287gmCk9F/TwKzFT/W4LwaP3LaCW8z
/jF+OFN3EqR1TebtwcG0DTMeJoaf2O/kx67/gqhoZLsVB0itZncDo3YrDJvPNwJavnHamVtiJc67
C015g4DsRwS2vmUAtV276C+nmiJKGexkRV3K2rvomM7HeKGuWIwULeY6VlbwgqwXqQjhq1IdvfLM
Fw+EBelquA2B4qRe+GnI61RyV48j5zYN5NL75TRTiurSLH0kR2TJ1U4DdcbOwtP7cFAZk+YQzk2N
rfJsaxn6uv/qWX4SziPL47/9vizgteB7Nw2OhUaFKPed/QBvHrefVRQxdTX/Gdu0WMbvOc+C7GGq
IoJFAxveS6oILtesEX8VQkB2jD9qmKnMfKAsW2n7Fn5UpF7GJK+9eoakkLORlqmxtmCimfZJI9Jh
AZGtKPJmVao9v97vaSiN0QLaPAGFo8KXNXIKVKxl2sWFqGWEznRB6RVX9uw3g6Dgxf2r6/9gpl86
UMEshDLhO/cPF21LKcUi92m58/ilM4vGLf60igk3EPDrkL++JZdHCwiJul07D1V91sn4nTfX4Tjn
p+YXUv7C/WA209CGWBi3sSP1YbVhdl0bVEQd5WqDvVw2ArKIPnyLzpSn0EKNsVnZ/iUCDsw+E4Jf
bsLjNhpP1+taujfUyS8dnf37OUPHY7VWddRbDZ2hLZEgnXa31zlGQXBV665SB24R/6SrIpicvSfK
o31onDuFm14mYU+s1P8xgZ1ashcWy6N5Ns0tsNw15FZ5WUGyrkXbd9QKuMSOscey3ETxM1t3rn/0
Nia03PnKPgBFB7wa0mZjmxIWytiAPJmaIYw6qliJtQDcNWdsq+PnpHJ10oqGcPiQB+kc3Pdp45aj
GlLCpbLbek26K2bThQRODR86FVfoTiQtqBBgDkCljYs6nJkPQ4iNyO+HwFQfbSoqs3d2un649zf8
8KGh/yPYaWCtboKCWycX6AtGraS/KIyKLCOuDlOaS2rt+/YDaiKQAkN6il3veOpQTGav4rALv0x/
erKVEBmHYGU6vaf/m7XbEATRbFsoFSoArV0+GRMJmy6jQfUHM+DgWNXF6B3/gegctf5yNz4wx8p1
r+Eso7oSmnr7L/4VqyCenKnbOTRyyRUpyDyaOeh9lMsXif8SBe9TmHAS/GaGWl5C8pnRcirxjj44
1lhc3L0y0l4e+K/Rp81ULOiN2Sh3LbTtYPD+L/oMYthca+yycu5qTbm+decS+x1GznvA6mW6qHe8
XHTt88iWLEsVkAtaTaJw3izKl45oOpHrwJg59XxkTb+7xTx/fmQ+Yb+zy+KYhg1kCC5AOb4NNTHh
zExON29JIe9kGTmviW6jO4pTuWS7ahEnSBwAnOh5sF5pMRGSRYp7hcW/9H6fzXobY6JbODHXVA12
Bl5n0lCtibZ+3WLo/AVq9xl2jqpFGVrQ5w5+m7wlELIrLfd/vuP3ScuHz+ZtPSGOUwzS2nbAmcLx
bP0dZ7LhXnyx3WFXv2oyqc2sSTTRwrQ5pUs6x5bExGr9sCBk8HbZ1auIoStmfW0JJDnMsyn8GLt7
mRDK4JUlIb696TQi27cbyeyiOmBN7LTJRH39S61M6dpr/4+0kKUjk2CqKWdoiowDgDfmqck+T5WJ
mfWYwvkOSad6VpecZ/XIu7EYyDbEhnNij09NURKTQL2GZcJMXun644opfkhdRsLOFYOL0lUz8G2n
WCGVWPy6RLqZJj36jkp/mgHi+Nn3i3FcUad3b53CVf0Ao7N41HlpgWWxymTAogGqnQsZN67mq29j
7w5ZYcGVLC5UxN+270lwUIR2cfsz85Aw2LUKP50FbBWNlBe6FVWOXl5hdxriZlxgSlr1oimV8uKV
bPSTvs5sA8leICTVnqrTOJOi32LNpI5hsIHelQX1YLo2VfrBPA4AbQxZd0/zX8mRtEOWc+ZBRo9q
qUEXJzwrb+CNPhR9IrAR/axesFkqF4eztQOQnnFS59JCtXHV6F9qhpyrrX1IWdsKhnf0jC1Yp7TL
oxz10abG4DfwV8DV9EELjwSdsS87Mmj5akcYWo2P8ZJ2l0pHrkWBbbf7I8vc5IxzUj51ZAhPUhaE
ple2GAV4EGKLuEzPUxlxwBfClxJ3K/E5POGaT+E8zEXWg+1C58SVAdQEiJcnNHzW2yxDYGnrrEHx
bAzfaVj/wb8yGLg5DMWl12c498qceboSbNUKfM6dNZYf8jvX+jBAFVvdFzemdiLCFg84u+kNYOKw
4uwHtOzTHCC6AIKhW7RTGQ9ZnIf45Z45Bk8CyOum8rDsfG7/fW8GiTBs94oVY3ITWgL0P78e5Uht
dA4wck1z7mzXTl6XYkwPdDzbFfHKjTX1Li9lJocRXzkJv9jl41X6B704IVIVTFLjEB1tmfYoY+Ut
dEcLrlSPYqVyGDm5IYSgYiGxPPnBL5Qrk2WYDEdB468zn0VHplVCuS2nHEVD7TXBgeIbPn55u+VY
ybkCgX5kG0rldH4L8F3ovYjdesfGYZVT9baHWpGBETharCnSpsoNrm/CwsC2eEJdIFi5JX/cTf8q
NFJm4IPTFiJkYeEPMxhhd0g9hLhR1YCOJFVAu9CqaA7EjJEFlWwDGZoDhKWqTb2/97+jAMqFjywM
CY9CbVmbnYwvtrW+UmBkBcriGnb2vbsoZGoVOYFtHn29Gm2zFjSx5qpoL3MSflUb8dyt6YOWZyQN
bdUUpNIcTBK9RI2H3/2coNzTPgHiAQlrhvNrEhK2VnM10Qv470CSqApvVmCGkkrFHqxRJIIYtAtH
kSvgEkcZ4KXFZSb/jJyOz2kW9VjUVTfgdioK0WxmghQn0DL0ylgBRfkaRcAXqobv3FnscJI5cMAz
t0ntX9yyP+IqoTkRAqsQju20/OQFM8+13YWGJR56vYKfjI/SEbXz7Ut1tEhZbJrDVxu6z2J9WBP9
q3YpwWQJ7otnItjL2tfs39yPP3pB2VlAOGHksOMchVBX8cBNPXFD4XT4zJVQ3TsXqrXZm/85RbmB
vL8G35UNr7EO1kvhggxL2S1qfrjXwC55PWlqWsoLezzEA12pNripcJWmRCIRIdmE9G14KHZiZDC3
QhoT2Y8X85IvVdloKmXA6RJAafeXCDZdkIbspA3iT227PQbrKEfXyu5Cz7OWgZWLR3MsY7Ond4WI
JOQ2depXheE/JK2bc94XN6xDZ95rrRN4W6j4hVLo+NqZ9TNOyYcXywyXWPwsQ53sYQQKMz7x86WM
VSc4d8PtvF1fWc/WY2ggc6wbvH275LCCD08IGeAEcoFX7M3tBoWyYCwSSUj7+q2MnQnLNxqF2IdN
JF3BEgyPhbG2ELA+PjEkE7tPnHfTBJuzsDgxXp+g9bupjvDNeG2JkCPhogoQj0Cb04/UvaUAKrmw
RhRs4LLx9q4ZFuUxigpFhzXXTnDZVVfMIM5CnMpSLLAW+lJfkqVWy3vRmmwBAYDa7U+O3W4EApLZ
AJUd8UjjI+xrdS/chNEl5ZHEU3lA01/m7onMw2tW8Lt1Mj1rdIy43oiAdvteGZCULzieZv3Xq2JF
36MqtNOUpSLYcgVQ0+B5ecUrcsNNivR2PK1T/d/g36mTXRRtRYEeLkZNo8+FGOFUMu59xpSKy2wH
C3QnxlJCogCH7vvpxyISnwoLM4cj1ptIpKYbSWOEsblgdzgG2s9sVo3I7OBq/WbdmSLNVcOyO037
japZBMz9UH4P006vtqPyWxNc+rNUS4j3aJz99Gp2jTx5IhXJdmotW11+heevUyJ3NAcQn2yh0v6T
O3ripPr+u26Psg4avUxqz/S0cj+E0L0iZA74exjA0Ae4psa4jgLAaWPigjHlLEImJLG2UyqUqN4x
Q7vS2kEOjrtkD+yosMWL4jq2EdbQe7QA0RPe4a17MMvvthBH9rVnN7jP4/V0eZsJhz5/CEhdbTzT
Y1BM7LRECJi5MYSgz4u+ncKEaxMCubv2ZnzltbqnSbZ3lvSPn/H3UBomtYsHKMK2FdOVDAIadB7T
viy8ymKWSPYTxKaMY9+8x03AsjPXhhYiFoikfMglOYVH727w5gJxumdcynZ9hwZ8T9fLBb2IHXT2
xFLM6Q/OJIskHZuqwUSrnAl0wBRHgAnopEuFlQZOswijvu4EoqCu4KmEPBZiP8pGfTAND4V6G88a
GE0+x17W5Y3I4/IXlu1bM21ZJD/ONFgdWEFA0mvA/aKtJBhiEdK6JLOSaxIjt5GqqiFH+1QJz2Ug
PDz5c8/zeS6v/ULA9RRr8aFtYjoc6bhVNwnyBsCOEYppF4nZIjWOvnTH4stf0+8bwGoT8k6RmP/l
RNHNNAv9G9lLjhpxgocKQLvmd1lOOktW+GZRCRF7boYTuo77iXxWStfP77vsNUoeJ4a9Zj1gYbID
KL8rcwQItPpomtQEuoRPmVVEhr15799sNl0jSyBziM4fkCVTqZS4aieyaJzWQpKE/unDd7yOg5g5
Uxa4IV4QUEBodU9dkT4AAeuBilRvEoWyE6ovlrFtoEXc14qKVo9TYb+Ay9OtHkxpE5pCg9Xv8U7c
du8guQ6WRa3DAhuHZLurdAZJe7lkh/GWCUT3/aXzfOdjv0Pwb3R5wN4M2bFi/mqPKBVVeBOk0SGd
FEBZSK8oDMQoqXiLGS3si21BC79E9fycd4rSOwbizTXDze2NqqxAiFNyEoBwm2faQodpvpChFaj6
2MJd1BXsatdKJxHy/o1kW9YnsLUUGzeGODO4s/KJyR1f+wlQZ9I+bJDVeFoSZKuLKcj1DsCMOpb3
USQKFmj5IIVSxKC+HUbaP7GEpf7MaEyDA0sX3aZekVZNxR3wlJrB+rKxL0wcqEcjw9zOiEX9Tj61
KR7zQXvXVVRzOfsoGQ6xHWQXVA44rp7qCQUAGtH7inLmekNW76TbCKpkCR1IZCkaExnHdQGrDfzc
x/Z4/gy7gldK60RdKukU/TRvKLtvd2tywPyJ4B94/4dzXe+spYmAdZNNjMTZEHtMPIZ8E6GWbvbv
AyX8eFlRA7w36+QOrs6+Jx40rexz/UgP+C+ZeuiqFEtZyU6HdE3a1LmnxGuFjmnqS77FsvmGiPZs
JEcR8rQ4R5LiOIRCQc3oXFhrBJG96LggCMU4Q6IfaoC58ftwGh1t4MnCrd+lRi8KN1S+WcN06F+P
ZhJcFh1EiKLqx47+B8vtoJz6JfiXz+L+Ycor3bCfZWVe7SjoOzCzsPFy9DXlyFxi9OFQSV9AVlXH
3+JPFePCWisqvmATyoIOKErfL5EWPNv08zu/or5O0wBTyfW4IBoCOS6rjTNeC/Lj9uEBwglZVkzg
Fd0UcAkrW4uoWVYwiFRbmrXDPwX3iDBtoaAu7RQq73uCkDxP+JKDntj4hzFO3Lzcv30KXpFFE7sl
rXY6cEiLnRJrtlkZ7qbUDJnOqiLfSMFL0ZgAK37+psoTpaILXcupSeLulReUVedH1VcwCnj50mwk
pHZ2MnbK9jdZuFripbadxarUPFNPjeLnUA2UdT9wKcK0KX5C67u0WQGrhB9y0U2IHBrV9mIZNTzG
zgR95Bpdo/f7EX/k63YTV6WHBv27MAcA8BigxqZmuLlHB5aR3Z5VyI38HiiTtl3y0gj+vBVqRMeI
Dflr0wzdyKY+SC4iFkMHYja9EG1FlGDwER7y6O5d9hXL855dVCjjuExP5vVG5aPh7l8opm8rKMMj
6OB6qvF0UbxVm5wd9MaM9BG5nwdxpvgL3uycVRl9Bwpf6+dccn55huOSieb2ZPr1DLQo2B56Gq5u
vnGLJsDqeepmPVu2L46uXWtig/XhEu6Bw3/uNsc+PlSfvko9AvwgCkA01pjofIjwut6d7Jm6jSpE
wTry2E8w+7POwERtdA4MfrpWTf48WjEqAEv5gZSLF0OrmMcowNfRn5j/db7jetTIiWU2lPvmmClG
+jAFa1QD5aS5lJczjcEEPuY48MetQr+1ctZEGavdvo2T5QfqS5FSX/eib20+azu93zIqX/+vHYa3
6eUEUml+q/nS7cq/lxfRkYQNQa9N1HL0tnUT4vqlibe2HuOT4r4wfnITRvvauueTMcxC+7RHX8yA
AO2fV705d2z2WIix+HWNBCOwP73WwGaUyhBIEPfgNclwnRaJU9vIWODk7HOTGWUBrzdl2anmYIrD
QIExog65qCqeZPxZAL1hcFua4muvY/d5jv8JSBxxq32rIZT6jM8UgM0uyW+GA2CND+FAHphVXMce
bLWtFErQ+D5I5ptIiBV++XVJGxOlukHFpgah4OUvbHXfsqvZ8oCzmds9i+o0ZQmCyJ8WhnGFRhmV
xYa2W2hz/egttf5qUHB1P8d55RzpiKUwIGessxCMhN38IrdFo7G86wQGCwLkyW09CoBQulHFix6C
DIm+xT5IUzO8xklHtoE36KUTNOlfh8Abyrdefse94MeKhMOa1j7PX9QVguLWOWZN7dtNRkt4GAW2
fa7kSgbpDLxggu2MBzdlUhtuZpFYB2J1Sjx89JSrjw3Whk/hQaifB80QHIj7eo8O1MxhzctviDXE
skSR/sCtF2MX1WdhLiv/mnjs4tqZDCI1wrjblbwkksLx+rGhTGBKhY23iySsw8x2xDLTmQ194Qi/
xyZZCbxO94cA+we8XCfjJfPx8peXgb0ePhuqkYMF+gIUEGEVO62TXcTpZOzFuSkTMkSFV+UBlM9d
SO133uFJxBB8JION+ZirH0Nh51w0yyQNKLDmshsbA1SUTSdaELZUycAKJApYPXVXKBx4iVIAOYs8
mFnVoNYoPVi6lNNJWZOyJSyxxSr1gEV/0jpL9bTwuqqUb6vfkuZLe/7EIWbq+w45xJCDdpUcapMi
/mjRMlSL234LtF94G9GGbLFpw2ETWq9mXcQCJt5IVCIAkdNSUwaUJjwmz1klSae2U7cYlz/+iegl
phia+x/gkIJb8teAFNNknlJwxuXcVfZ8ZzYYu+gWIIQc+FI+7aQLNEB9RmF1V8+zFz4b6f00Ul2X
renCqMkZ+C9Qw11HthFAZX+8jDxpuFZhIpM+5GAJe0zQXetHuHWsroMTQb4SgaNqWi4v6W05NOku
dBHoboGiz67ZnB6hRur/fPPnPOCWuXcFeOjM2tVkZQ1T/+MYueL3RVKWLY0pYjExa5hcto2JsP+6
z7Zh8dxGPbTkDhq4DlgWs6ta7+BgU2cW93FTnO0Q+wALbJpH/I4vj0IJkLxfFnXUmO/LS/+Nh4R3
zT7dATTx5IXEVLLOJumRbdiK7Vp8IISdtRu9OoRu1u4qn4qPCXU/eemNOXSHqRTClIZxY/wC+Wt/
m7+WZG9MVtIkq71aTrVXBc86sBW89M9cbTl2EcOhHPk/t1F4NQ5MPn4vrfnV7vB8Bw8YODuR559l
wWKF/1Pu3pfN8ilbelpVaLwlhLATwTOA099oik24aw5SH/q/MWQ3zuDbgUIcr3PYeKOI6H4BEWpz
ibM9Q4CpSgH4PqPuA/CQX8sO0rkkjD1cgFXZJ68NrL453ig3mstBPrhYfySLgsxk9HZH1xHAf+gh
6GlnN+9w4EdbQ9Az/8sgB8pBNc0BCJ+08VDC7kDKMRL9o8O4lnGPqWfMmzx6CISuN8pXgNgikF0o
h3lu1c93Qvl0tCkKQZE+VhvW5NN0o/QQBxtE9EAXj+/5ipNRpJpoXVJ0+cOnSrShkbDteM6xmOtX
Y7Ywkm8sSUYAVgcWD8IHdikcbg2e3sXkNRyv9RRhzR22sU9vafaLBy04kcNMdvGzVkzAgyzECvdF
xR5Ng/LCd8norlccXUwf0d1uKSHaqWxTvBRBCF3QGDWjR39bBvOmesQ6UjQrJNMCwqWLz0FpwQWb
Eh6/Y2SBy0lROvwKWHlUb4w4uPMozxIBHUgKmi3dnlpjksz5nOIu82FnWJk8PqfIR16pEj0qN4ml
VP3WjWdguPuJ9zBnXPG4CP3ZOPAEhwUU3C/DREGwLYt45sx1HeCUv+hM9J5FQg55JOqfXqFrzYXd
sQodz6WVsNiXjmV/GkxRmFz6MqQu89a+8S4Fte1iXx5GYJ/Tx+ISTOOsDEE6VRgn4Aae9kcR3NZn
Bz6gQd8DUvF86LHhRCaETJQgdQFOaXEzX0Wd0C2F2SnddNOkZN8rG0euMwKJzDviXFEuvoMK+e1V
dWMCpit//0R3J3FqEsMTzhD/Bsi04bRRU9e1LQh/zAbu+iKLXPXUqZJZakxAfOVApNpI+83H4xh1
EyCyYd8QXR9ZQAh5mdSU65vs0F9L9XG0Q83s9WiOsTK5luwD70GfuMOQUN5fmn1LzrnA5hr8Z+LM
CdKngBzOpZh+hEHU5V9RBW0whPkaUaBTA/lBNsTKChy+ug1cdQTqaie9Xtb2M3p9ev0YkoNeCajn
6KrmfoPA6fDG8bQ7klqSrrojuoHUFAI3VvEKjdnGypatAfWaSVqJvk2uYqjfoqVxMd2TZrNl+RdJ
u/FAo2dMzd+wo7c5Plhqmc9xxCCyzEKt6V0KQTnaVA8EfdzPW9TNap6i1r/esbwJYbR5JFsdqGfg
Ar9NaNcjLmPBUR3P+hIWQDilBoyyAKgmUNj3Sv5P0bEKacFBJ5H5dhMTMV+3+xROmohHyPc/9A/r
AUWSa3KzJxWwliXLv/0NcrLoxk639U/FgQo8pGFhn2CmXtKS51yMkgJB8mKXYL1lZTXLZaZV/lS/
6NUpJ0hH8w6gxkSw3Nus6D7w8Ax0Vkmt6y3GuqxrsYSBMDauicNdJyv71VdnmSdeFrYLhZQ+Tp0W
aTjOxe1ZVCEP+8efE9YNG42Evd5r/zKjwUk7mKh8/CIP0ju/mb3hfM5wlh8BOS8QMuSTFubkZXHN
SQE74dRb9f66dBE/T2E4YOAwCKP1LHc0Cf387faFQRlCPc1kawxopstd6bYy7+woQAcI8I7/hY68
YX9fSdA63Th5++serqqUOyX8uDYu6fbNn55Te6qFn5NzsWqZ6Y3d6yxdvv5MzbkErGXve0fKCRFd
ZPOjO7YpnWNeHAtSicARSIRIKoLGkkNhnqz3xcybUghcPOEK3ABOkQcFFDByrIwRsQ1f1CjZFMv1
pGj/zdDJWMxQS43Yv3rYMHTlGbhp2BQJowvFf3LcqUyrdq39Fvwr5m4mr+qkdAAuMs3TQ16w6O2j
aZ0q4llzSRNaVfnWK/eyEY9MUSC75VOHBtNyI8qbEZorh86i92uUEsj+iMoRxy6v0krbaq+pjTPM
ShTWzTMFQtOR8E4s8F8XOkPNJdRLEHqWZE/9O2G2b7p6khGe8d0d43q8FEMnR1URBX4lIkU3fyVk
jxs6ME6Rbwt1yh8n0TUOhGXIkKEkmG32jIQvLo0PaLRUs2aAhvi7SxNapcc548g7F8ITngnGl2Xq
LcJv+uQBB04N2efNPwQ0RBKU3XnwaJbHOjhpIvJ13pAtrhGcZxYW3V/kQVyJv+HtZW4WY6Mkfbql
Cnsg2NiXFDg0kGs6no08B34ckd81BhN9whY2Ywia1G6x9AnARLG0I8A896DWJg3D0bqP+wujI3i9
tKEHKibjcgUBdVxcl6Hy7lbeyA/CHPEt+cNywKgOxrISKSTJs7BXUtEesphgRfoARo8zGHEpmnPi
7rPOg2ZrkI7sPmQUAOm8h6f0igZtuHVmhFj0WXCCQ+QtGEtXSaK5tN/z8h8SCDurIHe8NVF7CUz/
jdUNIruO+v09sH8c1D+/FnePkDO7Wjze7hD1dYWJHoQgxNQmyKj/fYL0ed1hPSra04eFayBq1llP
dAMOfWs+mzRiDQTpjVn+9kN2n9s8ClUsPhX89RVzAcrysftSFgT2qskiOObRCFhjfWN49dG8EaYN
u4mEyqIBtLagdPp4YZ85WBMMfyTauYfijLYdKr4tuxV/PRBvN90xXCQxa0KsrFowQ8ylCqmoXccl
Us2ic27VGf231XlvCVVtlSdeCqJxF0Eua/11q9mum9qjI0r476pZgqsD4zAtS5+1ZOlRUeOtrPgU
NRuvTCQDiEhDpC3vJOg3JoL8ONZaoHUD51RauXylN2q+s+bLKFtufQzWnb04Pbd9JaJQWC9YxUMI
yp4BI35OdSCC4hlqqLw+qOfoMEObDsqzsU61Ig9kddnACfox9u2k2Z7B7pCCWqHuCBq4oAa2TowX
PpweZ/gAk08UDw5rSQwQcTAg/fMp8dRnk4Py5qtQpWb7VLzAKuZhZQftq84ydnRssDYHfJB8UH7u
MJoe4e+QQVVYmTpYjwJxpg9E3QeoBQkliRwO5NRezYIFpEoF/SQRuuAIGPa4+716dXTSH11545DK
gUFjBua/wfJDfoM1u35X7AzHAElU7qGThkpdhMXVE98AyYHaN9xoPUejE9zyEZsqLLV43QnC2dra
ethBKqQ6CWQ9tqZVpE8zpp6VK+dKaIlFjtuwrmgCqD+tVTQnr1SvGuB/HHNuPQRHM6Que4jnambM
XpLQPPIltDNVSHLZd2WOvuWsO0++jzfQQp5rZL5M/q5jc9v2ouNwmLZE1Jya4dvbH9NQ4sCGs1Vr
KF3y/HnpEEEffUP1lt7n4CGIyKm4sSDh8/L1oXU4jPxhQ/opjSq39+OBNV2EhzkAweiDS7Cc1Uw5
iY8+3iU9LG+Ti1n5rkWHEFVZZed8ATYK9QsIQRKjN70tJDOjMdikEBT3ZFbpVcRBmGB0jcAu4Tnp
12ql8/SZS3de/12cxI3x79mHEBJEX2ZXqKpNPpPCErBObMpng1O4thIdBKe4l306VNGGP2wP01/O
ZsN77gM+rR2YCEU/MTM66qhC3eYP4eC26YcZYz1IU+eK8N039JChmDYY4jaQgGm8bk7Q3AWViYsf
+GbLojUXuH/vXiUdlnk2gyREHs75gAz8CgequQt9nQs0R2MlC5ouf/GQLZXKykL9yqZhL8cvCAqq
UTbYfOXr/7Kfo1GODcjHvdNTDHJKqiBjyXWqQ8jWFF2tlPtJm2AT1RaiIEpQiqvJUMVB9/o2wvjZ
meA6qyfda7g6epBf5kKES1YowTlBRehteCON5b7/2Q2mrAx2HiNt71OxHDKhMzOjdOMEbBvJPfYP
kdoQ/S20ycwFlrBg4VoFlOfC3Ipzv6VPlBCTUpkZkBV9tRaoG25uGJwi10OodO9JF8kyNJMCCw2g
BP1MosULwCtQPJDYPPPXl0g7URKdeY/X21coYkWi1vFLQyg3aC68FdCLeoXrjYppjm4mDS40anUo
PP9S84tC24TsnFY08KA9XDgldd4+P2BH70wijGWYJxv0tmBCsHR9bv7ipHM6LjAoPACgk82HbLFV
xnfihMpYQYS9NaCRYqcnG702NKg9UqXhj7idEpKEKMNccuNKtzyhnPYArlnvt3GBWdC35ppq+ib5
moPcOfjDGPCxX9LO9RszuqknHnLC+Cc1ehN2p8ufYqhwfkZIVFGRRsc5HEm8lbdmjJk/5ooILwoN
RFadoPkplZiRGiknNiGs1k6yv/K0JuiOlmSpzNJWSU1aysJmjTWMRsbTsSXRHsXluT/bdEwKsICl
eW61+tAuEoDzj12Z1HiOr/k0esx/odeiqX5yEZDN2ukyOucyo0GqTlLMeUmkPpnmEbAznsu/FPN0
JH29ukI0DQS6V/0y0oDehDxL3qI3gceXxYhtzMCqN6fKdEorNhxMb3x8T1NXaISWRCi0hEE2su8X
fRXOj2HuMs4Oo7/+WgvUvdOY2S0zHw81sMpdaxFeJ+h7ZLYxVH8nKrgaMg621xzAO0/pjqGRK44b
ujHTOB3VKNjNd4NGKuPG5Y+TTRWonejzaWlj+J67RylrdwOanma//no+BCZGYU24BdDZFmKIYf4U
5QfmisKlO7FREKaIIHHDB1tDd6Mor8P4WEJOETp6qUH8ilZhAveLD6Tem4p0a9EI07gMvk/Kn0ML
pYbWePZq63m9MCictaOG19zhHybj8xWLP4Q3P6ZM2xXcrAILOjULiJ4HFWoQg0Kf6/RSoSm51Ysz
kM4BmOzmS079A0CxpT4LuQWrX1jPKmikIwGOs6wNRW1wJStRD/t9msseMCv0ZSLOmSk1KxB2mJu2
PQDziHyFvbCClXFNB+m42TlscGs02+sn6Er8tGzp7L3oGB1Urb1QH0iWctOgiBPlR4JhVeYHwVmG
5kNhjOILHCw6hEJR+x8KyjunvCJF/NpDvZguI0041o/SqiSennU7d+QGsxYRoiYbmen4rxyafT+k
bFm8uYEfXBF7Y7+BUara6OGD/9SAroSu7rL7cCfXymAnERXTd1YKZt9INdBlxuAGToyAJukgbfxZ
fd2h/AL173QP1vwMgMIzu7Qt3D/cU80N4Hdh/9cTUx9VXs1/u6KSLIBjxFXRMsknOcgxD/y+bSgb
cC7EVpNd4+TZBLxvmHD6rabu+PSp8fzJULQaeYWgC5f+OFJ0I37phUkEfNlkbeDnaFAxMMmeOJrm
45rbO/wpxStqLkscpSP45iwm9ql9BHPyMf3lHvIIMdpWtGc9FLGY1SrqmViwdS42nX4VTBF1j7Y5
Q/syGDm/kJZWxEpFdh2Di70VkTl9bu9s7uhK54XvpSzEZAuXM+/zKjN/rpTiFmRzvyuUJn85vS21
qLqRSbHIfoWp3yuDqka9ih471vZOhKgqXSbvZ4miQaC5n8Zuouk8bsqmBo09eNKWECUM0DQpvz+h
tsl/hl0s5rdZgtoQNrQIVJbWhksFUtWRN36ARFQIZKuccwI9H2n2JfJbr94EQ+8py/ALxoTvoitt
O3t0N1qZ7NejJo+ykUZT9UerszBiTXsToDOloqmVglKxYp234nyv937FzuuWdxs3W2ZE3wxdJM/y
j2QWfGcwWTU9aUWXfETJvu1HtB8FFCplYyGCLSgwLkX+BF1LtTg87EShr4bOtn9H2Ue014FJkhRT
NwVR1/Gg5T7f9XmFpnSW6smMXc9LmvYRDxrN5748NTIpxXGKZquRAv/10CgY+m6lMDzlwSoTaFNM
+RsbWdKhgOBKugAj9MVfq2+o6eeEDmqJIJZgrrPys9ysmK923UIl7YLlmz1Ivd+CKMm/tswqSW5a
X/MJhCFNWgn9fG+p3b6oe+EGz3Z0n4zUy/q2/sfoy/HVJti35DO4m9wdtqfDywDePDo+jPQvju5a
LB2lBVGKFniMK3oBe0vnE2/o846y0s08u/x/kQHGg4Yx8/mIfkBE84puci1WvbgQBmxwfyAbFIdg
TUg2LauGv6AmcExTm5ts6Tfk0vsBJqjPRBGcuQuF6pG04DIcRqpaq5Jrfw2BFRUwiu3TgSVCOP+S
45+vLc+CnhBY/FRmyOzKTtBq3GEDEEOADMm8Yp0Fdk5RDS//9BCYqJ654NIoB2S/SH8LFdK0xx+b
xuUsr2kH+yf26jxVzDE2hxv8/H9OFv5ld4bjKqaRwRWhY5xwmWu6dq6Lt7ACJVJ/PHm0Ea8/+6iY
9YeyR7nqOATXB85Wj4JKmi9glpEzYWwDMZKNNLPOm28hpj5zbobuSxmcwkr6n0Dri6btJKrsnB4w
Ff1GaqbNp11LEtxt4P9kyHzk6AGCxIfMTiYZ5SPExaKouTJXne4ZKQSPm4RtK6JaOxog0bvo947c
sWYckcGJ/jLhkXDrfwZD+Cx5w739JyDLWmKE2PAGi6W+F9DRo3Nvm5NW1bmzHGFHVgWoBgoY/Q5u
k5P7sQSriyKrjukeLGsxclFLStn+Vh241x117RN4r+MxXTi7RXKawwn8n0iWa9KhImPDNPZANdAa
66yC00O/hD0gu0zhBaco5C7nTOiSSItTAUhyHVaCl/gXCzLaZrZ9FfsMRw0aqLWJhxvrWmBWktyp
EWftsv2KhPYe1dUgL1dxN63IdwxVMQLk2jUCmd9HYVOrfPwV9VWL0kiaYzhzDCP4OPYMUkwDr0RN
rgFaLO+GgyN1r6qOBaw+5BLGY9YEhJIzN43kln5YgxshAs4xr8T/SiSR1/bLEKJrl6tziFXvarGy
32hBQ+A2d5eHOfP7dCSpVlwmXD7k2RjHA5AEutRRsZx7uvZLU+ZQoZU7jj5qYuaCPFwTXd9UFxu7
3/BUV/KH627fm5co685zCGrT8cjKQayUfU1CLwZTSMq5eZ/Ua6W2Ldstfx8amw8/HNiMoMSrdF29
QFOdml0kwRiXonLbeHZeUF4vyVzfquNTGVOJ22ZR+sLAJDzXIfc/tkgHR8mLW37dKaFfo6sEfnxP
AQ6ZaqACqLJ3IEaLb82EPNlW9MVUtZAGFsyQXIk8uZxtzdNxmVoiKKoHw0PXl5uZ6iqVWQF2QuQ1
O5C9xwJUjxGf8M5olD29MuzlIw13m2uti91yWYdmD1QKDTscSFA3mxfjGvzeRxAHTNVhPHPGuZmj
IjTtsW5cqtNqPdiMnKkRGFB6QAZNmGMzdtmANK8sMOSc3cl4pUyY5BGok//rsIBuITTzi68o+WbJ
hYkqP6ZHZKN2QlxVV+EzNG5i0EpnaP+Bf3gqYz8Z1Tq8cnCpCVl0e/V/NegpJJRTcYEsRzqxmpow
U9mGGes3vKsjjgWDkxnMwp3AyBR2HqIWxJL6syXtWpDPCm0OFT7bq/9Zj+JFgjZxt3qSyg/0Z0Wa
5Mw9+aDJPgY/Ja2RxYUqqpMMu9cXe6Fomw+iCR488JRHS1WfmHezBdlWYL+IX4BabT8EAuk4+aTe
RJf+9kCWWPEIeMIQTNAix+uvzjqHzEAZw0WrMcnSPRivlZ8FL8xPidxmZxRkO9mo5FBFijmw57hT
699srhxHyjMJSd3Mh/6JNDGjQ/2kUTBLa3TNSd51xqxeBvZ00qtKaeAZkiQ7C4qbXpZXWKPyxIT2
cvCFCG6eLsttx0TdZolhm7iBODhRnbddILrnZLNaOW2m1wsveCGANITpLrr7Z32MsjRHxUgapD7z
YZyYpUzHpnCCpR5oq1kFrTuLAQkx9Tr92uZ+oUhpF+KWqwPeykv3qu+7jTPkwSlSCUGTHH6/yLb3
o+0RwebVdQWUKrdJ8ZIB12UKi4WCCfxTq50+GBSZpGzctoeaAYHS64cLe2jmKVwOQeCmedyLC+AE
m5yETDwIGRxuJjjcOTK6GsRPxKXA9X5honFcIXzkjBMTcA6wMjD81/qKY0+5xH2OgHvHBpeVU6+t
HbwXRr7AMXPZ2i42afZIiJ6CzjbSn8mkA7ycFE38ON9SVpFlYdpydJL3w3UgMEEFiSMU065INVCS
X0fs0ipVfn+Yw8ktbMslpzhoYqINW/PyTQ8CEnuKIjlzunZZ6WCP82EpqOISQ29RCW0jLbUSwU9z
Htes7xIKe7gt/Rm3ZJ5uwBSI3TJCikJlHfDSPQt/xA1zwd012G51HpofLFtDf0EdcEWhk2bYAljL
JRcPMRQDbTHFdBxJSNoixxnOvj7a2jYHst1qUfqtgscvhD3DMEGJpnlTrGsdZx5HQfg2GheUCPiY
rGGq9U9nX6CeKx9m22YxBnEsAHZtQlI6RPLv/QuOjOQi8Pz9IWLwE3rTSNH8lbrSZunINwcJACHU
TceL4wrcCrYZB+DqasQjF+rL9bw5g1rkgcIWOOV3LV1W/xmGHq8kTLP1FTGSXWWeSo1qRCFyTI1F
T+mhG0cZlhUsWdu+++VP5IaqxOnHEQIWsBo9/z3EN6XWEwamGMO2vxuTTytNNcuAA6OPmoqZ84v4
45MtINwoNTRP9TG/oFMZSY1YscFCmJpKG1rYeoCMb4lAS2LMGIponm/lTWxitkm/iQA5lVeU1YEN
+T9am/yEbCGtTnOfZZHAerhv7eN/cRDzOKd3O2T7PrRyNrvl33hJufkz7llRAKCCaNJw57yLVrdG
cZPLbjgCje4mTMk38NROCaXhMGNagj7rPFZlOTXf1RgdQymhtBosH26FRPfL86tzJ2IHbM/S7AkW
OmOamvr5wArKw1e1n4txBnJ4uk+EuNfDfgNNmpU6iPFSbKC7H3eq38KrjZxIOZIeGkt5UL6VO8Fo
/DHXWnBySoPhEafiZ7J7WRqUJTFY48npdJyX7oK1hZTxPngOMXbl5VpclKQCpZGGwXBAQuTJVGnl
afRFTxMmtfpfJzjupVOgWGv4ROJA9vplOpycIE4QQsU2nB57dD5HYIvyPwz2Tjb84YlOjpk4DhLw
Mu3ByfDsGOzq8ri88KMIc9GQ4Hpp7SdO/N4wvfGQlK/AR/bhfENB7b+Iys5T71PNzXAJw7bGJS+D
AyJ3tYUwQ9BIy47pZwpgohhuKwkl4DRB/mygB9sCJpGCAfbRLnqlEFoChjMKGA/+QOfj3udne3ty
Ca9lgqg7d+heaNfeahLDs1thQ0ckMkmsCB6vf3M1jxVxKOXiNUKRcKSPQlS7sSGKS+a4t8gLCF2q
zd6f22rzWnyDMF4YZqVuHWP/a+q9TjfVUaV3xmlfDg8O4nl4UUbk+B57xcZkXz4yx++zlzLQ8DNI
BtffyjRf82udQlF6Rf4/zOJqbcYdEcopZrUUTccKECermfND/AlhlLfy6Id2UKp78lblCcfe4kO1
/RsY7t8+gUPucQbUAYixnF+FTwvHB/4nM6+9yIynlm6yMN8WhkzBkEcfY1GN27MKV3YLBQg4Mq8i
jGEiSeByy0yjPN7eELc/OnRDO37klXxoGkneu8uMb+YJurf7wajnBVd54ENuMUrIWADqGd1Fln6d
gKFQNRLLU3b2Y8MTmLrCL5STdcpEj/RYxvEOdlmGVtoUcVGR27zQ/8pg9Flrn7ECJADH+CQWXfAs
PeVLRc1unD9ZibCCN86f8tITQuTNv04TF/46Dg1i0IpLyTw9U4Ko5pI0TqFi/w91+qWessbhyLQH
hqqPiLK7HtdZGFDRasOAurJIoC5/k/eRizDEMXfdLlr8klEhvWgsUFsAqWvNHaDBzC6YKqIJBa0B
ZcyKiormPvOhndb+15Gyud3IEVubK283EOYeJg7tBe+ODf7FYULulYpac13OzOdTYk8ietKLedSs
3sHdMmgjfW3lEPncETk4Z9gL0o2T3+/Z+BmFlfqe26PQmsB2yQNszjHoRGPE9F6Kw/T08xrUyyIs
F28XSI1sidXRhV1djufgae8SD1JvKh1XzN92n/aPXKJWTDaVasACkDrqT3ORapx5KXeWrWd9KMmQ
P5uF1W7ghsYHmVk2vv4Sq2ot35bC8dSm1EViOBFUD+9pS8tnm4eF0RFfdW8r+z4PpBBK4ktYlB4U
k+tpIJcQtSjbuQVKmdrnPLTNNfAbcwc5UQ5FX09qKEnFWtTJ/gcOQ/uAgy40Q7tgN6hCh7rmVkBX
25GutYsQ8SjKMQ5i7Ar7STywjKw6FODnXGrWoiaCgonxAjbMtB+lVISU3Eh6ua4nEnU9qiUWjFmu
BQwVu7b0SOBSk8NQtYN4C/SExfO1pWcGGwrLHCxNFhXKdBtf2cNItURWBKlAl6aiewsKOD1HGIqf
JTL0IRAXEzXtg8RM3lIU70Ha1fmU6rS2S0rAlQXQom4k4H9I+RM/Ux9GXOpG8RMAs+geY9AyYf+n
jfjLtiiREVTprd+CstA/j8yijUH5djRtM/Wnh0bnZ+Qxygze/7Hn33vZKTR8ECNOUulZs97OAN1S
GZ95ehG1+eSLrlI9x2pzFl1R9C1ex3u0jySrL8uG07TAeTXM2U8HBLihdNkUtTD5Sjzg4wn0zeM5
5dy6FU4Su8UzBJhTLV+1h3SVpzMtiVoWoCBy8a5mu1rSmjxfHCrX2nEvBLFZ9Dy66tXgR10j57xI
VPaoRJ4wUIDe1qM36QHa5g5hf9QFxF6pLv9PynLJeTXsCM4oE+m8U3iRg+AE9Cf1MWakdANXi+1D
orXq3f/vjCD3FVpzxSO2E8i/0g1WHFmA227gTUERtnd8VMDjvsdz2fkzMcQMc2qqTpYhL53K7bK4
PXVNYxEMOVylSPbjNEb85fZEYoTGgsCT29jeVKHRKMRHXxGpIsm/sZDuC4bwsz+Ffal2fLBXcvak
0TnZJZErYQ8z6rFTxIY+L8WY5sN/Ebe4GTm6Ncj6GSGP/vW2i+q16nbInVAnjeo7c2ih5UMEQj7v
mttZFRcpnsnpvlCpW/OTSJTJaO0G8knmn6peVlhJ+05W39V9c1WSyQcB6twN+ZHv+z7orIFc8sOP
MSkmcqvV6pk4T0y0GPfeJtgHWWbFyJVPJjDz5v1VuC2VJw5LOpht1Ka6eso1ccxI+NsbDZC/wmLd
CHsdet6oD5HH11SBZUumMFOmLL8Ld+UaLtZPlX9+iRpLmhS8QSPzK0fi/AaPG7L9QA2v8m+HdkvL
WIp4KCwpWZzY6NajpRMGNgDdzc7dB+gW3782iCnAFmqoSzURDznC93SP5f/fANPasDmDlaaIo/Qe
lCuAnGnCqpCU27U3M8n0flGuCFXVMWtYddpZm0/MwezXMh3aKe9eB6N/QgHfYmaCInf7FWJ6Tofc
SXghggzLe58BmL1veOrhJVt/83udGfZlIYrlhqCnBI9n8yMpa+dzCi4GoSKmO5+EeYU5vrdzoI9e
wUdOe2kb+1xiP8BNrItYqRwCOThePzMl25Oh93ZA0lYZySgb1XG+P4Rpx+/gAPtyPhMhm2x0YQQx
N8ILecmFqpDC9fCvTZfH33bQF4MKXAM9azzOHu7osFUx/AEJNt00EWcr+wKd0VZp3CipBTTej5Sl
cUrUm9hlZgUJFNvP1ADSxiKGrEWvpXGaKFBwS5uQ0YBUwy3qDJa+TPcgkKIVHcf7JQfWwGnnt6kt
yAcWJK2vFi+13f9ChzsGkSraRThFeLE0aL+QRXdKveb6FXH/Z7Om+byFutugLWHLbsP/nzIxav48
xPag3lu1TZ/dYOnZFjK23ba0sXvi/OacC1fDu9RWF+WnsbCj/sdcfxBmyksxPKK6LEumFSdcaGE8
v3wtQR4RNDsqGdJWI91QDmk14r4Fp5WBCFZSxwdfiLhuQJIVPhHUJ0IIJWemxVodXFo5is68DvWJ
Yy8BXmtGYLeGSqZebw6XqLdiOjfmcbZP0b+nnPsvflD+ERXPNcCb40yZNKia8s5KJykNqgjBzE3b
3lP6Bf9DOxvIKnUMfWkUzkApGjEPERa9JPisFxjaJu7b5NLbVhegKAfi+BdT/2TD83QPh3/x/fOd
R1v+4CBnC5TvIMUsH5HA3/5dsfGxSDcQnAiHWSfLLFV+wTw8LYraKgBgPPn6fHjKKPkU2Ga6rYcG
YbYOHwo3BYraQYaq1OwmJ2IRpsj52PBjZGUGs3+8oYp/g+4/zydPcKWQEnm+WaD66L7+Ec6X0FIP
fvKouKM87kfkyKe78FDVbBs1Ske7l4q8cBhxoJ/1EK6xbe4WBGzws8KavXFv0mZnzWHJFMdKSwRR
uzCwQ6BU6w4v/wcqhIImuZBSFnl9aE7NmDOHA3a9WkTYcAa5YI3FpVjcojQ+h3vtNNOEDKLLRKHY
AqvU8PV6TqpMcwwcY1HyHl31i7RYac9zK6FZQTnC+i8ErVY3CbM/OAtti7q5S7RUVNaVlUapdW9r
nv4Xob75mvw4MeWdUboJrSiWfYPvGNtDJiH3WsB5O3uXD2Qc15wx5IHg0fgR/3/o7YdOsd41r9WP
n8jkgKSwjqZtwMII8UUQFljo9bJ6Q2HnwSuXwkbCnSJrsM7FsMF8bPkJLDF1PgKubDhGqZAHdWj4
kUl5/rkFaLjS1EmKSwkcrBbNt5FnNXGD4XCaxtF0vkd9zCAfRYusypyNvWT+bYdigVLCob+c5h7H
41JTAqUOGzYg2nbhHpfvS5uRd3zJvcAXQg8ynSfJ6D/8ZO9pipwruu95Lc/xCUy4hhCXhkKgvfzF
J/vbO6iCI1Yqh3ucnhzuzBndinsqouG+vbFJPmTexmAwaZV8UQf+AoXxlYcw5aaZsNVjAaE+GU+c
Ao58siqhDoaqwgiu4TRBvUEZvl5mKRfms9eGYOxW3WEGRPs6AEsruFECVLlulY4z3eWUzpqDb7Ma
+s9f4v5rBlvIIeSWv0+Q0eUX85GT+WjkyQ52hms6Th0AF5Akq7weRMmXBqOxnVYraTXsgab0Wqw+
0d6rwf6bU8D/XABHM25A9SXtQGKKgUTJlcFhpySWU0FtyYz/+r/0HAL/7Rd76F41iV7uKVStm3uw
t56TvOG1iuVyuhLWYw0JzmwDf6BAyITT4AiBjTRrtIh0nwqJLEYUV0p/QqnU6IYAydkZwHPCzqc8
ZKY6tW7w98VAU/GT6ascTS3WL8K/D9DAJHp/ZH7qWjTW55SqX0H11VZnVP+1UdrUkj7paOAV1Pd/
E8iupbyppGfFIpgfEnkV7YtCtzc6DHYsvkJhz9nLLf9XgLkxgqCQ2Cjhqc6nXwb8s3p1ZZuw8V6e
MAWEK3HR8OZS8hJnzPfq7Hh/2faRj8oHy3b9l/JuDMkJee/d8nFem6GON7LXv75rCvlnCuyOwkme
FdCtEDGKCfG0J0GPSMSghfgUTjGus3hhVJ1uuF1KP8EXy7PrktGJSHiE3lYuQ1ZW4xj/lW8vA6QS
c39gan7UBQDOL0Cyja91RUsSj9o3VryCOnYugOhTcQn/snWnBTegKDxYTn+mExSiX0LIwZQbqv/q
TL2E4/BhuLhme5wojBYO7dX7mhBXaU3QH6TEQtZRW62iiAZf+WA0/mRGF6rqf6ZdVBRZvZ23GuIA
MLv7RXXzg/pOlJgOZYFpPeOlaOUwvZWh8MyxeQEUMh3l/rxZ87CHs5RYT2IpChPzMJkFUYLMgqMB
ul9qIg2QogZf3jKTTvO6wzUCKxUgWMuwBG+uhSWrNsz87K3C10Gq3YMpyvgp77oF+9VnBpOA1Nt/
m1K0uelIWM5MAy9HOFUNAbsDY8zxOMz7QY8wBpindEdrrX+4HcIxvgsJ6ER6cW80WfZSqBJbyY3d
eoxoHeIDZz4x+WlIJrtSbSJ+Om5oWfL/q5cmgNV0KnwAD0xGuNAwMGH09JAncSSCT7b4yOLDJzs5
TGlIoMeCV/2DJQsH1VyAHVtFkZNSlKC4/Kys4A/2WGJ7emlEopROL53pc1Q3tBvEUC7VWlsPtfnr
YwSyeyQTjX+irRtAid+boptRXnq7jPnxgkH0OilqUJ3Cn6m32ElJi8rywKJF8CAN2a3DmBr0rVZZ
Sv+bcNkm9JXG/nw4xXo5EEZiOFhVa1cSA3vcRy8BpyRyEA7JmMAnUHwnUKG7Km+LcPGWtPZgyCUQ
94o/UQpZ1A8jPSSBu+lJZkFV7CEdbDj59QCN9PRRLz7C48aZYoQrZW3YtWSkeThRr5cvubP1Q0+T
ulSLRdyUkYdudUkVy2DHVvluDBHLPiAdiB1Ua2MTyeVXR6iH8zd0qlIrWBbEYb1DsJTQYcstcwCP
C+14bCjYlo6vVUkPK56Hnid6Y2nFZOCpHxoNmrENCcepnY6axGsVstCTYSU/upujwEwXdaTJZlqZ
BzWzWMqhybyvnr8/3alJABINYXqY1qy4J/J2w8dGBP15FmJ3oGR5Hc20wd8qvwRY/oRzszguOe59
5NBhokPKQEeX2s0tSBkuY8J6s6HLosVr7LNTG335sG2fLOY1vFaH/d75xHrgB3KouWHmSCP7fecw
LBnd2BSS1rlCwyZEMjzuMVSw3E8iwUIeDrMzCNhE3rsgd/AGp08yy/T9rzCBUcRuwFwqzvuJXPHe
RN9Qdg+oURIYxCQPkYi/Gl7BoxbHR0kbw+Tg8Bfk3jdOGOn2+0O+GX59/hfLY4X6lc+FB4kNde1w
BcBcr7lMOzlQ9j29OzwJpHJHI9m0fEwJM6Gr/DYTiZ4gg4TFr0mTKF+0ag7OVlYs9i41Rg5R22KG
vo40EJxHlqv5XhIgCl1T2IwnYiTY7zx9P8CXpXst1gLjsksTGPlTmua76yCuY/VcmKiv8JcA+Amq
kwkvIiu+InXToduEZMkjcMGQp4JiKZlNBLTnd/WIJ2FZKlgacXniuIoi99+WgDobFDGFu2Zxve64
Yekpf+jRFWu+ppiKopMKAfdHupLYkKx6s4jl3w5dJJoUnKflH428GA+pq18Jyx1kkrHgf9El2q+L
hRQ7cyqbscnplY+6Xoi5PnYVF5s8jEWTi1T+80LV09jSPlTkHfNMdTOq9kPM0CDmAh8tovWWsrb8
SFWuHja9t1GED46Ii1ob81WjhMTpYKAamKNUGmdRu1WXlXGF6jqwC2IfghjwRtUudThRT7z6Tt4u
Spek8c8kId91RgG1wuiBtnCjJuLj61824Q+4noJcjIm0UBHYd6j6jC9VYAYmxFANcQ/JnfotAfEc
cvuRjFHzZ2rXi5hNszC7reA1uacdm0iI0855n2/OrnSLCDV9u/rpkQ5Q9+J+UjRAxfwfJVlZ1zq7
axfwYDJAE6H9bOExSQ5+bhIG1iJsWnnahGXaJN0E6tc0jNSdsoFB5tyIqcBivt8T9Vfk2tnO6zCi
MDc2okLg7yZpsC1BLZCAqSor8covdblk9lAG//iD2nj3K53Azu0pofFcuR3a8X8ha9VS6Sgp1fHv
wAK2CKDBnS2EUeJg32TVTaGEW4ypgk7CVpF8132CVQjjcIsnL80WppTaxtZ5PSerhuVRx5o9qUil
pgOYHlSogKyKjE4Pc28gFvGbtgytm06vyfUbXOsfKAQNNKrZKg++TYlWYfp0n3rk2+HSI5hdaPHe
hwieQPwDYK9n4uSNehjZWc0WbV5+ApU6oakoSUf8eyWv9X4PvPlM6HOCVqIixWGJRA3IqMPESrdj
bQMizM25zY1vXcqU13GpeChlFC7FOgC0fn/pQy2khstX0tJpghtUVlXjck5ulnPZ/mCJB0intP0V
u20bA90X4l6ihfIhFo2V4l6A/yQ1v3vaUvkWWeJx+6v6VlqMxK4QG1gS5NsogBzR2B09SF0sy1w6
2KcbwV+eeiWVqet+r84VbGkddD+H+4spaZr/paCCdMrVUcWW7ABucjbPj7mzBnZe3ZRd7nssRIiU
qG44eq7gHd9mVc7Uc2WvVkLPiW+n8JuTEVRN9mhSIe0G+Q2s3A6YyFZuxtz8q6h0jCGyB/kjizAI
whq9Cj004fnNjNskECwQe/+pjM52SHaHHwH15AucfIgS9p/1WLeCIZ02prUcbxBsEUVc8Av8ck4I
mGrhsKIvq6BbmO0xW+0LTiNMIZzlNLjxOkm5ra+LJx8ZufUd+P0dPhx410YQGJLGc9uwynXsbPMj
vOWId7iRmQcfvuWQtcSWKF90RfYe31Dh5x0wA65rh8jNvA0LHHUsbI5C89hdn1pReZvs7lFJJp/2
/JaP9qEl+mKJ+ZCEUBVV+g1QQyvGmA0a5n+sSIDNUkT/MFfiT67vpMszkk4mTjfdJGNHL4J6A/7E
A/m37uzLnf2aiSp2w4bWpe7TiTryoobATFZPjAqr6tecmipgko/6dIXsBfOM+yImPWxz0Yr5eVgV
+3NIRjk0tjN1BiqiHGWsa7/x7Wy0Um6ipOGX1XsqyLzrtzEZX8Jn6N1DbVAs/PUjgnTWqRCjR9Ok
68VntseojIf20qjR7nAtcBSvhBvGB20j3Wyud9DKXhzW3z6fUVlDaskU5JfXs5l5Sc+/9fGM4zct
pG12ZR6JwqBymd9vlic6vxsYvDjU8S7mxkC6CwH27L+T8b6CaD+hsTfwgdilUzfiObRtW0N7dPqS
yxPsHo29dHc6JD+TUQF/aYFczbPHe91gdpvoWlDvnfgYhowqLsO1jcdQiaxLZxJhTiU59WymWC3e
aNx4hKRSZlOoKqmtJdDzjLrDNSjo/fvQzAiwrlP5WOXjnm96/qFi81ZjiX+3GazRFMXX6KyLKt4b
HHBWO2QW0iug2NV5YJZLptq0Cse7/U92/b8a10bLlS4OAnJow3BQd5k7oiAr4XaQL7xYzjeTPJOc
qAYgjjpqg4yjkKTK+WczFHxiAbB+3Ey+wkjZTTti4aTvQP8b8xC4xP9ewx+l9FOFDjxGWdY2z7t6
8rdwisBn8bW6VhU/pM6YZAx8YUFhP9KGfIOKBybE0JOPLXsnw+F1o0dZplLYC4PRoZ73EFR80Q3Q
Wg7mXHYiCnnHHdosWnGRewAauwBvwwpxtZEgGrpXdCp0kisw4lqw/a8g6udHl47/TYWh2Kk/C9dP
rhV1B66wFJNT60yOtubbOtZvlwxK2F6ugSkDFF4PQ0lcDTjyeIpc+GaUghVmBTsXvZuOrhjNHN8n
u4aaA7iEYbhqJDUP2vibWXXQJzpYfaNcIxHc70NYNtiQp6SUFvv/GXm0/NrAiWpsunWl44XgFRHu
WG5V/NsQNpwTYXSD/Tg+WR+Kbr6GCj8fsge2Fqyl/glyPpEZTI8SfYL3SSyagyqYjeTEv3cIk+yZ
ZFce4U+nbOTIJ+Vq8yCjeNrgmIlZpBhib9iswMZDZQiS/aTXCFzjT+ZGGLU23Nbox6N6B/MxOlUs
7eRbugYaSFq9QR3Qxjq2xT0uebeZ2+Mn7tttiC0KxsL7LgjWXE7Dzl/o1gBvXoq+lEwbHwwOxGe2
tS+gQf6tugnLl8kzLuLNUt+C3bX9tmf+Y2TyR28aT4JCEDN7sp+1sm2WVHX7LrGjZW+OclhjbzL9
OkIsUBHIDJ3w9nb/k3GAqUiQJ4CvfEHLREyIkz11PivH7IpqFA25PvBaoNtWw1b3F93mBTFk8339
A/oan7T8zH90Ll90iGlUlUxvJbWbIBN1tG2KJxbht1nSnw7zx7Ese8YXAd6CDIpxvNnniv29+iWH
vz/LZI4zX1rQB6yzwfVNi3vqpvSRoaTPO9SD+ULxrM7836V0VVPQa9DY0DABLGnKWeS6Pj7PB2sO
AOl2pBnrsVaaYgU/O2X5HQAZF+QGEE8x/jrkwZ+u90zB7OUTvhGOs5IiHX4mO9zKNfQG0iAMd+aK
u19DgJCewFxe+JkP2QwQc/jDCcbztw1zIwRms0ef4zunmIdkFhjtsmA3i54S/3IZAVMvoq2m1hSv
mGSbtj5XNCqJwBwQhKGAY4gy6IHgyc/mKxId9WdUH32Zx0jvDyk0PfEl9CKSv3TU+FawzQus692I
PWAFu1sjfCc75JrEok9TFYuHUDL7gjF6jJVHygYbr3lTjyx/U1j45d1WIR/1GpUzSSnzA/hfWsUJ
uuJTr1y77OUMtwzcG/PmnUVv/Q04ZFrgtV2XEIN+a8Lg1OCT+nIcRwZ5S9bPgvQssFGwxjELRMgB
B6U1W4HB5w0jFt54iBhl9tV/eUI6wcFgBJyy7q/HZ7knBc7hCqQAgywaNdH3t1SaDFbQrOGzAKnB
nZ7tcK2oJIF93fzXIlqPquhD7W1iULuvYyIH8fFHuNFbDmtkzWHsSglwPt7/aMHQgI1j+GMaeLbc
abl29W1eacJbJoh+MVr42E5xaboUAURz4Pn8k1j1uubL1kX6P6RuOhzlt7Kn+lTANTCZ8p0i57sb
FtN0wEDEBLhMH46Yrczk161RwCB3Omn2MzDcqBzDEQ6C6Yldfw/EAtkPwtUia9vRwecGj3Gs0fMN
XjoIxn8Ss7qmoktbCM6LzVNmG8PJ+rI5AMHzFcpCyjiacVTDQR7dxGHdOVG/gezB1TwV6MTsQH/H
O/eCCbqO/6vJdJXGVfIpN8ML0FGxurhtRC2oDO/LIP251M6OqjKLVXfxq9/9YvaZNppoviJtuuIy
fOlqj6baYemmou/w3IjUnefctNWobZ2JFwU1xuYLv2F5KgOZoGuOsPbci/CcsI61hxiq/SwhT+vi
wr2EpBQ+rFd24zkZTA7odTZT9PI6A0COCBr3PiWAzZjcq9i2xWoGI9A6Q7NvdcDWtEsAykaMqiId
4fNG6qSZ4wdvpVyk7YSm+Kvpwt2+4kGl4/1WBnu/wdZbD4xVN+/Djw9dTVHhQWjb1k2DeclASw4w
Gp08EdirgEcv2OdOH/fQeHCe1t8ew9BQphMQBEPCZk8DxF4wrwvfSmFuqMgnRhqsfrX+cE35TmRl
Xlh9fMFpSBg79V1zBvuXUORFgaJYjnTR4CNrFSZeSLK8qEIAHZVC6n02g56EyD2nGhnoIShNP3G4
lWF7+lGQPPIyXmyScxLJcoEyvdwQFwQW+3b9p81NB2Fr/VEztye+S0Xq9zso7D9DQFdEerdSDTk+
h25dDir1QqY76e4dnsFPRPUWrcvlIBf4K4WFhlWtAVeIGFBhNPjt2e8Nl6CFKFGb+R+Az+pyHHiT
9Q7ybt32J4fILGTpEzw8yJRLY1t6qHcApyQVYTMjteMJClrTuifg1XOrpACLJwKhOFvNJGrytL4q
CFoaRJa+ZYlWm8MpxlefeuYPCF0CEHAUpuuyoaEApBiSwtzwg1sBBQ+Tru4r8wj8zLmb+od6VExf
SNiO9B6nPWHyD5eHwAb3R2IMKGGQ0Hj3KHOkRyBhnSiBRIdWcLqdUM0EvySfSqy17j6W5tvbtyZ2
xN+2tBEhbnp408wpYaK85CTfGPq8a3Lfs+XWcB+AqHf562tysTSf/Xx0ogcRt6Fa1r6Dv1BIarSa
BMNAhsgWxYyLfj0yZHlbpP6wfnDZ1Fhs28KoPr+tvtn0KR3H4JHZ7RV5gIcIY7HMLiZk2LmKae9f
wXvDJ1q5G9FeI2lLD4jAN6doZ+cc5Wm35qYYmyorLX+/jM94fpzi9/pKJjBufeOdRfg2MgV27tWm
i4uCOVrdIWvacFrDk9fTDXo0Erdl1/YT+Qa0oajx+/xkN49k7aCuwm0jtWe57EnehfN4XHYTNc38
x27LY7S4cUE322Y87pXd4zqXrsyTT4eqg9iN22zXqgB7BHiChdpgwnRSbYu8RrIE3aWf3R6gBoDx
s3MmRa48NPOGFZqbWAFmv/qTy4/y48bDtn1U7L+XL+gIxDCv0rLX8y0TtHq3IdN0VxcCsOtIdtPY
E1GX9600bVCVoJmgUm7rQZNWBvB+b48PEGgHd8Cx2mp2NiLTgUYSPeUVPBZDr6iRf9SbtkmVPnNB
ocgV+aRoUH5FDNFJNLxpHR29RKQMg+u6r8t1vLSh6OuH0uAgp+9UHFydMgnuI8GxDQD33j9/pG3d
508P111w9BYvLW1fTQzATrL4i6N/SJVHMVlK4SmtJ9ZrVPBbPowVIxG9s6QJCIi/mlC+6yhAt5rE
OyWw1KWrhF9wiWLDM3YidoXr2rQBBMRmQ7T2nmhMedRai03EA/wI9tNoXE+PB0RxTawgmpGFDYm2
eazl2LFExnHGc85Imz2v+IqrjE8MJ4i660wZWi+t7Zz4zqKmP0enQNqv3+mUbzkMShQDRhQ8HhPL
dFFbz/gztwWi6aULMJQm9IMOE0xWkDewcqnXzHi0Pggi8p27SMf3A+S4HjzPBTzV1QxAc+qtJ7WU
ldtOYSaVlQ47Z2VugOOf9N8qgcKnMREwC+uIaGnrdlAIO6P0aNqKrD0EbDnwpJFkUsDuHl+1mDru
9GxijvJPioLPe31LrvUjD0HOFC5wfEvlHuXacmO0ilBLbSUfpIkA9wA9odFyNmVffksnyNAyZiba
l6wfapnIJxLZ2V7pl6ABHRdtzqrekuGfGpb8hLk7HCI9hAxFq9XJlwpTdKQzzKKVs/2wiz+1kZXY
8uykMUYlknaorgRCg57BDTTVs1bur1n904Nlp0USG7K3qxrlU0Eho8x6hNrTJ5RNwsXgXsadzQW4
I2My/gh158ov75Lh7lsd/v0axrtrtN8FKONOGbNJVFk4n+hClqv+jqMRMw9B/FySVkj28yg2w0V2
RULHnN6viObXr/BwkhCo2tefTsULifK0oVn81Tj+gzoq7rtigXmchlwRXRgBnRZFufYAhdV/VnAS
bgQPbZdnbls9Vco/UbEeA/csEvVqPr7VIpz6tHqnSQeIc6aPMowyBj+MKygn+domqCYmi1/lJzJ1
vE4NZPQO24RmlBSOSDotNhepJaPcKKGRwCZn2cI2dHz1JBx3jTrNxCu/Y4vKqeG5JlTKkBnSwOPr
p1Zd16MIoNXoOa1YLoenuDWYqwLgqpxgiGq/SDFKUTd5p0jkEuiesukamwGVp+LaNm3HqszbfYiz
PdOd5NNDD+awzZYG1HdxfOVbvENBHwPqemuZd2EZmfGTbSmosUXrj8bhTwK23UtJJJvbHAAXcRG8
LIZrb3ZxOsw4kuJm72GNLdV3GdC/HUTACRBOxbPnq/36JAo/pXPdlgjo8mAX8r9Z+T3T7NWsnTsP
Rp07fDutGg709eC8mkvFCYq9hDcb8dvOS+SYaOVIDlW7pola+1ysrRgB9Hcp8UNzkxOnG6IWHcY5
L/XtNhCgSl1SF+P7TmlNO2jO/R285D6fmbyBmMhAjLHT1DbPo/ldmJ9n9rf6zJhuj/tV/3/U0L5x
mvWdsLZLi1EXjEaeTkhlKxTNGXdmmtOnbNYNEkB6+nDM9Qdnfw6RiufSV+BCLtdcTqBfK4Rj5IN4
LruRq3MXtL7s+1ezT12P79tiYC7Gg08tzWoJ+YpVh+BU8bcrzvs8SL9EUyP3/XX89tEnn+B+1Brw
HUbMrTsFXAXHH+gLeQ6NYFgPceGqg3WzJcVfA+djJfGY+IZ5mvb38R6vZkKVJyOeBxvfhhb6cUI6
kgjopohAg39RgTN9yojlmx/Ev8B0xc+EhXxSJQ8SiQB3SitXKRgEMWYSfEklCjNrOf6jwjTzcBq6
TtoExBqV/lqfRYoD/sHzL67qgNIWq4iR50oDZ6+cdgO6i6jNU0iYmqMOYlgwnSCQ9jO0SUFEMGuL
JJ2BPJBoGHQhsf/b27aZPBbLnR6saU1bufsww5YUYxyWXS4VMwtLhW4AqPwFrVMqo+vMe0N/nLPK
hekDe1HksHupOJ9EzkQzuqd5vuz53V4yVVhc4tmqUbRQFGay2wX0ieDJI5T8kjf1pTfg1oDka0Rn
Hhtfx9G1PsabgRCXnGMPexJYOJdzfNWksbhVfZVZDHH2UpzGYUIWI5LL8GzJZtrOCBscDbCC4Hc8
UTAOJ/YauVQ+vhlpqJN4EZKmoBmfZ+87Ce+rGQnutsJNuEFp//ti/BoW+KTFhKAiFa8QkC+SiVjx
uNxcm2LfGkKQwvr1i4x/aCiH9cCMoQy2g0LnPvL0Iw7Hbr98sQLI1kM5eV7eDKL3tqi7mIKwkKg8
lsdE+akCXOKm9G+SkgiMAbHYPUHLQkKMbEvilvwNRA8Ad7KvfhbyG/Zv6Q/0VMtzR4CHRS4Khqnp
j5xpgFFc8Zis8/IE6LmcquR1LGDCQKKUl1LVB/O5CG+titTUiAg59+VPKS6hcv0NAtuTk776mwa8
CjpMwYKjQCgaMBRHY4J2vCkryadC+ZQ4OsQzZ7iYluxK8gEmBxKYZ1/p5kuwTBMfOXoH9NoE+Zvy
zyRkyDiKdM2SdsajnLSn8184CTphzMweoOkKxHYtDMfswneRiWJFHHr+2a9+S1xrxyC47LtIi2XT
pGb69fzt/NX6x/6yIm/5vcsTmneHWOpvtbNdZvtvYpafg+LjTdy6KB7oLUxUDgYLbX1h6knR46eG
tFHsKMLuPAtgl9kfk7ClG9Zz1GS6A5cmZp3ApS4rCZPMPG5UREOkrQ8wR2qjXSA+pceOtfrkXRud
4r0T2EFG0Po/kd6NK2x4HM7ZT7AKm/XtnRW873KrL/kePce8dSOgqQXutsxXsMDKrdFIMNVFUJZR
ffgcQEnoCFAslhGL40KngEWaHzVTyBMw7FFfWBeuywvJMP0egyfEtreZu4BoNIfjdDYagmhUmE+Q
HlpX6TomMYE3v18cVJu3q2IoH7tV+GlbRQIWXMBAwb6dSOOGJ3ByQOWeynvrrPBTNYfvG1mPSsy9
CKTMZqpAWQTs0y2w+5gmEUyaL1+RyOYo1hQSTgA1EhKH0T/papde8HDtAS5BJveXoHuHE0PcMHaq
5isbYn4xUH8AyMxfWQ+s9Zxw8VRg3mN/brX8Q3Z6RzjtAafzbnZGKZYoJhbZpVAcQmsCLuvq4wYN
Pb0u4nguhJXje0yDe1lPezKfDFE4ZGmEMPxXYbzu/h0XiNg/1MVxWKInIPhJL3mF0/xemiXatZ+l
wEeUYpkd9N3gCiotMRS9DYeDTrOHniUspA8LgV7RrX/28kEdXM+PSd3iGhd6DsuiXeVsUYskPNw6
4o0KXaRrGdR/Eb8xh9Ex8BZFxk4byi0/lhWMHK4UkHjbgWJjZojejHIBCWVbKdBMbZC+S5t9s5tz
DHF39rnYVmN06yqe5U8DO48gSMIn4+t1nVrpHVHrmqLp09LtAb2LXDM1hhPkEXb01k5jjwaus2w2
ANJ0swGLy0ppeClCMLhzFHii4s7pbJNGh78NfNiLuchOMFH14eaL+uLBvAivhrkevdZA/tjl/7cx
NUtEV7ttuVgDxmX596Y9syHJyNnksztxPN8/z7zhFMrfBS7RKlrUgIL4L+OC92P6PwFle6gYPkqW
RyCcb625AiVtVylvCtNObQtuQXNNn7IoBq9PqTWQTSr6XcyP7NUyZqgVLUBvUkSzOZb7uU6wNwTE
WatXRKjIIXwkFlwys8vr6hSiUIbfXRnBv8pOqH8krAhqSCK8gjpTMboygkrE+kFkqRmRpgOH9+2t
6oPJIFQiL2l8ezpDym3dBC9dZ1sZaTVOWa9FOt0lCEgeJ59PVZwCi0qVLwhEEwO76pGbhnfF9qMM
4BGC194BxAjXXU/yn55/YZ6iBAZTQIzA3l1EjIGUXsY84qJw8tHA2el910CZ2TMSGswsa+GmHMdd
hcyUo+nwQTTAVr418HY1vSUTTL7SX+Hfln62Omq/qc9Cv3DK52OiIAMXz5jlys/pWawhf8yHyGMv
8eS43MYN9S8EAhBm4+Ih7oWViu1+5iXSOJ+3EqPiIaAc7uNsNFLLSAUYrRY6yY1Sd6M7lcT0KnQu
0MW0zKpLurd0Q5bU7EyYcM5RiSqVuYFLHPocqCvcekRtIsPt7mEMaipfhnPw9J7jRezEjc/Pk5Ie
mVSVxwR6kEcV1K7zQaG6owo0JFopdt2INR69kvnfJclcvrJrpdIi4sOFnxLuYgMOFm+IgMZZXmA0
vsQor94FfPX7aXvnahhJ8FXGczxRB0TP9qMXb1uFCKGV3lG5AsVC0+hztXp44tNX0DU/qGeCHTr5
yvozyBcWQdHf/D8Q9q8+fgmYs7nB06kfT098Ys7uuuF/apOHbXn4gGzGrJr0QgB9sPwL2w9AgOVd
SZYl+q29NRTrOiY3ICWxKm2ymlFm/exz70PCWHE5dDT2mvaUliImZ+gPeKIR6c2f+H0qD4HQ3Att
E3uehiJTmRZ+R70H6eH2uRecT4h/oU9BqOaxZTh3Y5T6lI1J/9RvAtV38Pq+0WKa0wzWipjtvn67
UyAEsxCD/insjsvhQThFgFEPlyvWo7oE6fy/SW22WGXY/Gh7MZswrPLq50tNjRLkyuqWtnJDrk31
Jh3A846AqCur23n8VTPbwefDI72sn2jfP+yu5iwXf1YXy2TdmgSdCjr7kD7NVcFLWDEfVfctE+WL
4rteVXQ07Mov7H3jky9bX+up+1HR6fVclzyV7pTrnlH75xhbKVQq80e19ouyYMpgj9LMN7BEJBo+
YhOjKp/n5fPk+Hkri2/QrJUvWYBz2+ALKsUjkxuceiGWDLOmvK6ViChzDRtwX2oWXVtDhEz9KbVM
/p+yCmvZ2r1DT4Gf3YDkwUDEEssk4vinvC2WawDstBbMfrHP61BXwYK2kTJ5RymtYc5BS/ZXAb6g
e4iklY5t50O8riuaRof6CpNFv8zcETHp24/v3duym1zaUuUXS0OiKknxKYao4JktTjFoCaXr1ANR
kHYbt/VRF0wjr2EznqxdHKllhai9FpxR0e30T53r0CF4tDusuhKUP2Ei2vMFiWXbX95UWzu8B6+j
q+vwiQ0P+anC8L8Igt6fQUI31+DX7XwhmaK6lXDeM5suGsO8Y4BlRHPPTyaaUmVlg/dyEsl6VxOi
e6wAsmdHvksILMBfi5TLcHeLDnoFroEibveHRJLzUIMG6KGCPfpsPpIUBHyJ1JR5E4JydXJMbDAM
/9HUT5twLuHICyWreaMLB1QAwZtmApL89IiawO0gRJesaxcnl5L/CNbc6NLM0Aujqe+3lpXsj/aI
oy1IYxYmW9DWlpudJQDZKUTArVjjBZSuYRZfGpsnaZUC9wyuBY0avrgmGl51RqcynAtXnlWlPqrb
vBTqd0+FdGagXzLyx+462gJqZUfVzkcXMEIn4zBg6b8kCjTDglhYBT6gxygXfuOH+D0wP0RRgTIz
b0oCJIl9sDdpSbp+B0Q2NUvhdrSclNUmsRC7u1sQlZo7aTsCNEfgMeQ6y0i836nVqm0K3Bh9gkui
NvQoImE65/sYS1fbHzRK0ueqWU4nmwSFPBSfrNrCIzFUcVz1gN/mjh52hR87jvZH42KWPMpbcAwH
CcIOWdtCF7/wqZfOp+qWhutiBywJJgDXf2opCAEiLrQV3DqjBW6/gBAF/kSnd4bB0dVsXFPLdBVL
pMi4IhCSK7I9/pM8lGLsKSMWUzGE4fmfWyQ3TH2cwVUAPXYywrgB0u/IvNCx4/tbYtogiqVIcmsv
pITAHvpe4zPFnumLBQcGdBwPnppguC3g0Wiqwmw3WWf8juv+SdYp40tbuaOqWAHw7+lob3Az0hUv
K5OMk8D24wWpD0/nJmpmPZ1GOw6/vhW6P7NUPMgBb/c/K4re2SHl7qjClnUiZls7p9cY9qvBm7NS
C8vERnxUzPJ05XlFg59mbE/3SZMJKVSAdbQGiaIVHUSfOsG6EVtdLiYzsLJJq6oSA3q/NPBcPIJL
VvyElecyP93GmddpHNecHzZyQPOd2C41Yc7ikYZDJerHPzjpwdAakGCIH2XtPmzyXFigXYgRK9pq
LA92SlZ+mjCmHMThpHVPugaQtgyhFcl1F61AGEc4yqdNP8gH0p/RYLiR2btr5Uao3qe31f0vpMvK
m/mk0M7fPAlI4M+GBFLM//1/Ls9KbwCo+gMhyY1x9epd0ffokFEsiezXeFeIOYVe0JEK9AalzlDz
3EJuGyCdeu1EynHSHBadKo0su8pUo2Srtt4yTKOhCas1drbV407cve4pvU/cKO8A+iB4XDLUx9Yk
DBaS4uS3Xm2Cx3vhb12f7ZIAAe/063yz5S2sYl5rDOei1v8bT0LDXIbOeMFThNBZUr6+XzKYYwxG
FYdlmlCUokJEAuOoVWres2VfTtwrRy1M7GMZcmywurQbiq4vZDBY+biajM0mNvfOhEiSeL2tb6+Q
oR3Tn0LSWMqCckrPDlU37ONQNrPVhy3OWsoLad8XoeEn7a+S7/CWCmYxDJR4SPQHVJJD2fv/WF/B
LBLg3JiHjgOkj4ng0Slmmd1df3m0/cQt3Pc3V1klMXeey4cDcgglivbdf9yG8fsUPEHs6AdVQDJI
bKeONWVo4sZdmGpnHgKx3/b1YmUHNAMZLkgA+sB4c6EbJexmBDXRLn/WbpAR5lta9rlmlYmsb2Iz
t/yDE62oe4uoIXva/rqNaQZKxzrfLFehQsHu3vW0Zksak4dMK3SJWQ6yJdAiFahJvhQgraJbx6W1
eCYNPDO8Emru+a9hJRRtFKALH19DxPv+5QuFpx81kKdb+3uNN4FDBzN69l+gB64WINrz9s5NiVTU
0vD2XinAPz9EVpf9rhzSWQe0Ce5+QtPZHj10g0gX+UAy8zvTOeI4G+EOi2RH2BTkHx83La+hDiOd
9l4T3UGgxvuTqQTzjFSdX4FNLTgHUHc9thMDRiK9Fwz+9H2DlM2iu5EKjPTYJJBufAvzgMOO2caP
j8S5yLqvORbNm4lnBFoWFsL2cnuX94WUkl8/rC8NGRNKsLP+hLvr84RgTcH12QuOczereVpxJmGd
WD3bvg7tV2k9W9vs2FgUhQrUlzGqL6UCHkVxNO7Jasyh8Kl+5h5Kwl+LXUtp2QJSMAVEnJEhaLj+
7ILX3XdEn6yro87T9KzG6pZdGHdL/aRqdmxu31/FgSA+eulcHFfk4TemUu59AyqCWdJkXAojDxi5
4Ti8ZeKfo0Rv7KfOEYZO5n7ClA8NAzDZVf2+OVW2V3zQejC4pBq4YTk7aXskBFWxCziw406SINK2
YLnnvARSElJo/uwP+TcU62VgHSwWEny/aN2NYgU0M/J6VbqqQ4aM+Ej9l+V5IGlz/LPuUs9dGT8n
fSXV/L4c3mbi2idGVusris/qs4jka0MnHCG+0YDONpuXioa9D/NuXxw4wknhUif1K96eSXeK9vZ7
h/1LkK6X2ZIJl1YIZBEVkamPVpDll3/+X6PFArZA8SGYshDHNR8Dl6lKqqL5UJaIVBYeZqGVtKMd
eZFroG/sBDgtK14otKibQVWRzNu36eKSNxR720omBouu/c4XeVwVyMKk/Vet4Vy0gj5QrC+t8ghN
XeJuhHHD6BartP+MmOFFcjCbnRwu734gQE4BClTI6oJxWlpsYl9lZCnTdmQWkRIfesjbxubqUbMK
4+bzMHHJPpZ0oVga1w7gyOi3liZQ6zkt2rac2zgSbXc2ZbTaIrAOFb73nlUv2ZBTsItM+c8JHotc
8HfEG9rcbuZPOYXY1h8kEeiDD/rUI5lirj5ucDPjHXfY+UhTnTIEYFQLN9sjPSM7BewiA7VLpo3q
xEdAyynQuxUSKH8AZQRqsG5k/LeVI1O9cPrmim7d+ruHKOBKnjr/4mxbrXJOngBuuMaSJKIz4Auk
EmkN/py9lJAgZAz1bQLOjiMCgae8IgwIp4Imbi9nRFThTK1J1Mq8otXQZZOEG7nE5Yms//AY7vL6
Jk1g2Cv0oofyFKjVb8WDd3y1TolpwXYvuFGyLmZ9pWoxOsQx2gXqxiDMBqW4hG1txpCNSaUfBAvN
4GgZ9AYxzH5bNb2uEn3fzcpAQ/Gkn3Hdm/9WlgN8PHLijteMXpNhil0Wd7VcZxDLsWWGoKjEBtyF
iskcKDLYlbscO1YXoSuPAl2e0eMgAb+xqCja/q6Nvfum/WBbSPqNixGQRBJ1hhshUiWa5ZVQCzQY
JGukXwcfX+4368+SDmYdLne0L5fLJWIbeZTxcs485vj+TabzBTXNitJL2t0nxVXWI3URZmy7kFg/
MJbgkWPvAs/NNc/I0hbtijK3xQYv1y/yVgBGth80aCa8HIn5oGI1/RmwkMydBEvaq1DAYxNnXmu9
drkhUBkSJvE3JSOYGWicHYsSa4yLxjAuLKWl9SLE7p4/esw9JDSgOQuoUTcQ42QlUYFDIGcBGHlA
OWGNRsFbPZeAPdXMKm/eZXtnC8zJH9PP8z/0n5ImRXtTpcFfrVC8xdaj5yjQWrN6FU+7IfLX1Nzc
ejvSc264IQsBW0mayGYi2oo+G2lot7vQ+hw0Mli2MrZaF02XRato5TXBBaUJk50Zwq2Y1/nKlt8+
/D+Xr9IbDUa9TASb04XH2bCXinT8KA4eFwFYKQobUBOxTlKzTyin6soCZU+EipdFZLbculPioO/D
d4mkzR/oow9YN7c84SWCpsV6TKUweQ9GQ2I9bIpwwvTeJpb9jQZ7JzfEOj1voyrjFP6BqiUWhbYJ
+9m4BrdgOiog13yRYBR0wCvqAJmnHu9gzjjO87gANKfnZnM73TFOm/zXGj15GUXD6+1KHqf6451G
gmf99fI4/TbUA5oMiNmTqJosXfujkffCChJQUxCdADZk5qujaxAkGDPBevN+y1BicYTPXxtyqUEP
XS/5LBp+mQe7MiXsMZNaieT3BXc78FrhnDUl2veMXAuHknryj0eflUV+8Ytmh56Vf/4/D3IF3fYi
aEJQVfObW+eOfdNxAGuYMpWOBlJurGlqF7z82mYhoODilEMs5w/FRsGGb5ExyXBN5/VasvcB12j3
YsQxrTykrg0cq1aSnrQ+gi49TIemGSDMv40QZtu+yMcv1AL57d9UN/yWaEpT06MVx0cmhH1zBNPu
4e37BlRbkanUniGMGfW99kGZvcH2BXA3c+2iJuXAPh/kTzpxAmKOfpyj4B5n+OZct1mDD/l8iCnI
9l6WJPEp4FZsRRM8Agp430ArxcN0Gxlu/Un/EB6qvRkJqzfMXcnVL2ijBiJu7it2T0ypDy2WbUQL
WV40SKx+pQQvPEmSJHcis9ZnDULfXDYLYuBs2HbGhU1Xv3KWO7eSe5PO5bp5XpN57DAwiaqmER8s
pxo+tXyAJPpP7imRR2F8/ZbJOBfdai3zUq71aapvpQUK49OOYSiBs0jfRhE58HhdjYrY89Wv5JBw
6UZxG6qVMbksfihaot8IYe/ViRP77SOHpi94x9NLNy/tnBgMWI/JxgjHRoSjcAL80tW6A5jw3Q+c
rmMsqgcuS1dQ2MkkZk1UoNErGJnSEhB91XiJmubeNcBQWhS+5mGhXq+CnxO+br9dJ761EFhNGQke
7jLWgLrUCKfhw+QehxcYQliTvZpVQWJzsqKUwdFyRnwwXDb8GkaRrFA/Ui06swvtP5fKZRKRnVSF
LrQfkoFGh7O7HyRfizsicmmFP0K//VLB4I4NSI+248Q/aNNaE+zvgF66Uaw+BgVGf/tEwfvvbo4j
uBlLVbof922wcB2pOZUAzmKXwVvvNt3o1mbd+GF4PC2GOo7jXqO2Ml1LoXG9uYdtQ68gc7fW/oJZ
YtLGosKDuPwUTw+0WNc9BjVMZu73rJpupU1kBd76S8t8/5q486SsnGIMl3IxJ8lKgzTAq2A/S/pS
3OFvXZeamq6nyeB+vtmB2GbGtqJBFsFhcFELIP1StNW+Sb3bw2XFDFe8ViYquz/uMZhZmDU9wM8J
TNSbJBMsWdOgExHR2hi06oPjPmhZPossQ+NpSRXGEfRjRqI9WrfuzbsZVLY1PctYDRoY9u+UPn9h
rCnTEmhyFaFrdW0cWrUuNxAoENBTEcMdMXHcn3AHg5nYQldXUKbSIdYQ66dDMRT8061FCAgcIbaw
7cdlqtNReJl8zyIEEUOqIURFHKCI2FqrvZcVOjLwq4kH+DLwu4s0UbSusXEojye0yYwIkYurW8kf
o5mQtD1yJnmTD40c5yyU+28S499Y9uBARpiEaFvFkqxip5wo4PZ3Idr78udXcsHz+VDJDZwxSJIi
BozaxwBbwQuYi/MXMbaHfZIYzGIQN2Akc3MqzB5DL9AtbhTHd4A52PVBXX6z0Q0taGjKOBOrpADV
49JyjfD3hgTxTzAzz42hmR61BlQ45lH44seXpF5jpJLHeznTh8YdqzbBZ+HWPd136aaTY5wvMFbV
dX5Rw/Yxw5e/OLlyv/5zJZVKGUhUDwWBvZ3KgE7SiGwDkf9UeTyy08rTEbo3a+JUR0qRq+faOUbs
dDNhs+sGVDK1fVzRbfWGBOz6RlDLTVXCLAj3j+rWN7H9dW8PjcurqDsMjzXSMEhpDOdu8cUei2e4
0OEmPezdS51QPeuZbNxmXNtH+QzdHUcoTpAEWnVr/TJYGvZW23Fb09MJlRhO6HHa8D6/ct/t3G68
7mTuUfBquGlFUdiOI1Sr7u8qFIiTpXOO+fnY4+2NS7pylb0g1VFtsAiv7cdRKQiOVUpGmJzYvhMq
cm/xAp+gPQdV9NzRpjMHwq9YzUIATIPkvx4Dpe265V42kHJtJGKtZIG1UW2ET+Cy9GQVxS7sVlTX
YmPISCGEknZaMFQCPa9CqP1DyQYHk/tegjBGmR2FgdJh06yOqyrmUhTBqd08YPB9GFHQsy4r/g0m
Wka8tB4vESuPl3T+yC+4pUJMGoqQBhqBH41cCuQrEwedpOegrGNqkW9Eu6yS/VKjRry3Cb82CKkr
qBSAfCZ2T8uTYA2C5SLVmPew/fABvRwdkBfveGC7EuXsXRUWmW9kkx1erxZDTFe4g063HJcnNkr2
H6o6YK6UVDC1Et4Sa9YY1Kkj8laIB91By3cUXSNYxVHSFS5bYCA2sUF8FOR7uCGUqdXB0riL+DrJ
xgwezfi558geG56ObnwH+JN1fDkCTDCtESPlWCPCbx+QMfshW2YTKTBNa8sqTSymgpLcvsu2PWeq
lzplE15u9zX1Vj1kHNT8T7lizZ+cZLH+q6j8w+7G2gy/4GQl01X+jiMOCB30gbruP5Ar+NTXuP4O
kHrsGDWyvwEmej1xQQYcdTJBtkpJyXZUS4ZTEpH1YWRvFmsWPG2cq06cpGfqK3sp+pn6qrBb7+i4
1yVaJb92MmuOoD2dzP2ekubr/+Wz0+blwPW3V3kyJMcAPhJ+cfvTjcbtGZE7ySRRuywk2397nSud
Jdkx2xRew1tHGhL/XXbs26p37vAZTZGIguc/MTFIVrCv6R5d/dyvQEpn2Kv8p94B6XQZo/h2TP4o
XNHODHkDiX1ZAtgHGUBuq/1kr/idZqmgxV3mS4ZDz2xp4ElB+5EDXR+hZdlYQxeXUTfGgVAaD+Qe
ifiPzyC7o7LFEih5sjCHXxboyg8OlU5NcnaQRVCFNqLtOR/LDCavKr4PWPiurZJzdHg3GwJPUd0F
CyyYxkLKg8rhOY9WRoicCI7sZDdSCdSWOeFmM3dUjIkbZZ28Pn23IQcJurvFY+cEMU0wldaK10YP
aHmTAHO8Q6MAY1KimmLbM4529Ob7BeyqnKpzzhA8aCkVX0GX5M+jknBhwA7f0rfX9JbndlXLLk3w
BCQwLvwLUtTQel6z/XmziwEj2DgggZmKuGYEm/4sjcvrLiri9yXShdjJQiKsLc5PsRph/5bKQfLi
rUBFZUC54CZOhtLXtNyMRmoaqyabX+r5hTQdndHLXqdajai/X9OuVUY+XsuTWcZJU5k7HKl/gdHQ
zbKuoDja1Qz8a2npBtkYeJysj1PDtQt+LBv/9/4bUiP4Cbx9/VsXQGq9TDFJFCjNmS+cqh6jQqUm
JGLW+SHaP0ARjBNvw2QdLg93UO0nUku7I0t0NJKg6vuViNkJMurLrK8anZDpF0zWFnjr4xkD8Tk8
xmaZE98/tgaGHvsb6guwIuJN9AXmzpSoRPnUorJxxAb7TmUPWveg2SU1UTGxXabI4HZisFfnMWYY
PjsOgwpTvS/8030xnJRgV/kITNPm4IBCtEcws/tUKbM+3kMeD8aXzu7QvlnXflgwmkAwxG3jMOdh
nzRT/7Qp1juEWWWrsbFuqAZgmnn9VvQ+LcVzDZnvfVoJpptQIMfpxYEVOxigRWT/JKbQjaHYlUhh
e4QB4B//AhaeYvfFlXU79ZrSg7CFprck7s+PMqpr5VC1IVUnU2pK13aWytqfTKGPEHcxqR9Ur4L4
BVndijIm95RsYQ2EZUSBiRoHiTjCow2DC4ZsDUhBVXtL2sDJCwak4+ocZD1Rgi37zuR0n167Jhdw
/iAJKh7BGT19NQF7xFJREeQlpiOnGzAO/hSM/ZAkeIy0bof+xJ0nVmgq3+iWeSDqJI998EBE5mAA
XQJt6/FiF8hUOZzeoousYD6LA1jWp9wdcqxfJDDxnEX1gm0vlArLbzyAneJZbAtsmZZ9tKnwbmCp
zqX5AUc/4blV6sahE0vyFYM1tXrzEDizk3Cm5rSFOPL4TkqWBzLCMOfmsdem2SBxdBRkWvoibIlc
xL6lTwOZ8dTfKIWvAecPOlYrfeOBF3O1LAujarCNUZxcpbs/aGzbFaCnLwHCFA6hf/DIRnDi7c5o
2pv31eDx6eqgbtVTst9d7GrXPZFEsn0OMRMGilowpHEX+/FrZRh6pKk2PTLfF1EL4clp3cbTgSHM
lfUUMHJOMi9a/YU8qTjWwSQ4FeR4q3FUMfyqtIRMdZb0y7WOa/nC7UnX7gm7/nOt6tMzf3Bd8QjS
r5VTGjsja8XIxkQaX5R0jyFtymbwezh9x8SKWuBfomm3vHevnwO/PyEuN68FlJ6ARuDKF9YK6m55
BgybG7N8GG6gNsEQxVpCr90vGpAR513tDUN9F/ZCe6w+YOnxzwUJUoIDNSoazUviyjuKJhQcyB3A
1afQfAAYxHWgAvNinRW9+5kAb41yWvJwyQCJLa9EPSO7DkP8Athy9sb6q9x892NRo8Gx+ot4oL2U
x/vU4QQKZr5zYL8DTNKzsympOPYbOg4fei6WNAzKea3Rd5BDy8MaCFGc9i34Re3Prb+M+bQkQi8r
EI1+OG7MFeyydZePkXSBSnaO3CCUnl1TB8oaOD5nwfCopUKZyJY2BsLmielpIWrKLdlkqfl7Ni11
KN1h4YN1gcCRhb91YEHIE5LUk3gNcZtNJK7PrRV+faWYpaad7Z3T/XmalcggXJhOFdfC4bRIEkYn
R8FyY5Cam6c2RUWGtva0n+Hi6W9ASdWYSVyIbDT3uhfDPaqbWDt6Q0Og1HJnmBzSsXI2zdnR8uW4
sx9QXCkHRDKEvgHA9FF8nIjK9XLLwKzhYMWLMj+pHkuytWrKlQMyiGenGk9wj4xqOtyOG27ESCZL
a32TYUIrYxmInj54PzYZ5JhZhpfmnP0TYdGLloCryJmKKsep3X7jH95SL8Z6Tgq2n3o06kYYS8cJ
TUgVHF0QXkGgruhPTT0RVhoeyLFf4CYpZv5dzUasH1dQd2Iyuk+JNBObR4iSCMMLP6zq5jx42vnf
LRRxGbqCy4wnUuQVathW0gDs2Eg2UKbh/qhQqgBpJvXX2w+Qbma1oPiShq2VNWnOw+PWPrgbQZ6s
NnQk+Wdp7X3WFijutLwHcMTmfXBI11H+aUe5R9wJIm6kgSzPTB07mE9pFGVluJKaNH/uOVy+/ldw
tPF5jO/FPVpWLDD99HQKPTHQXpQPqzDZK4P4Ysvl5MOABGgaUSQ6WZX6L+acCBFbLw3wd+X1Aho9
MC7ZpPuAg2nCl2mvIA7/pBQEuy7LMIz7+kiwLCWBdOsrCBBCpFPAjBMis50by10sovZRk5QaV7g2
pMGT+0GoeQAktc+hGyHaCGr5h6A3eE5OHE1ec0YCVhjogdHI8Z6AaCdkD1NihKw1UsflAEDIY1y/
Dvgjqc6np+SHy6LuXY65v6ae+kfiTFjp633cpdb4FCxnNApUmOOKOiKYzM0ZcDmsvqAerut4gSfO
uIskokKCi5X46O3bXvHAn7XBr9ARbS8FLA8dQ1u4xD0HwAemrJAA2S9W5gC3nIBk1y66KeGtrT+4
8zdSoFyooWhA6Ud5eLJ11oT8R1gNxXOqAYInPZ8MVhMM1SaG5q/lWqtQMIQd2EgHa6yfqTps+IR8
MJOIN6iwFltClATShXSiJ5op9TBDg6H/lsamWIN1qNt+2Bw8Cn10Nb7NzRftuJC3TDayidHbJve9
TV3bi2nWCw028u2sdn6Q9AvIPoV4s9qI3KA0mnRWiJ6oGgJBpaxIviRF7MXdhHOjw42Np3LzEBaD
rZqqbQgLc0rp/JsR9Tu7s76QUz+V970bqDfbEyXRkbuu3Otz11IYy39bUAMCr7/erBBbl/wtGCQq
fVCfAAi5FDshotEf+6jpkfF8hfbgv66PXQcIybhdZP0aLb0Nh/jMrWiS1OjsHR8/ED4ASxvZox2o
2lOn15A0zdWsFUFZQVYb6il8a1FOmsGNf0Zi8jSJMS+7z8oqdXu7bF0+DyJmpscGH6sz0qyzRTfj
C2s56FzCV6wNdGfAnlCsGB0iSr8+W0WJa+qwT13EpIKuiFvSsoUK/XrqQZgqLn4aZbnDie8wwiub
NvdoGzFBubultDVPtYR5xQWbcbqd0F0VbK8L8SGuLK0pJQYdJ4UQHoU22vSXMZr6fInP9MgMLb59
2l9glWtmf9KXWBHy1Wmsfge4QqvHwIR5hPjWuYQPXcwpFajMlWYK+H2W3bp8b1WdybN9PGIPJSE7
b7R4AnpqU9ldBnPHIJIVx/nRBVeLkOmX+N7fi5JuGEOVc5E2/tX+ztsymxaIni3FpORZ5ETt9Mgl
lObFfXgq/Kvg1FnT+MuAdNSsGVjRnHhug6mWcQM2ZVSznxtwjKMx4AL6U5f1zrEYVnicYqobmbAK
pGX/JZEFM+d3ZS+u0MxvAWDUAURu2dQfh8vOdIRdfOtGvVAbbzq5LIu7TQB3o2n9hdXRrWUXrA7B
Ho8F41wJO2ELPVZT6Kih0PnQQTSGONqOX/sFtrKhPTFamIkZ10hMIwWR/5TTZpRlACQ5KRmuYeA4
wJjYAR0p210lhbF077d7lD+dhCwdqC/xND8vIEJ9IofhHfxzuukenW2g7fV8iykQMzZcJCuVB/Ua
vu5XLhDjq0SjHW5NL1yiFatjzqT2IHQG9CkcIEI7rj5p+MkYYpYid7spg6dFzrwiSSkczR6GsEbY
s064Q7St3KUxY+h+P2JAlubc5fy1ICOnbmXYuurDV9jjtjzJ+0vtgjGQSRpstsWi17TxcnOLjdB4
mwGgQA3+3v4ExHJFB3lxoRIw5lZUEacUmuspqJjlHWYflpNLGyqqRNP7bj03YIKQqoFfU90ek2iN
hppE5uDd/1R0S922v4rRRD1vL1lSmRVZNyqij/t1yl3tGE4OYFgpsBJgYwSf+gc+vtP4ApYZKpN9
0DOY96DAJJWXm43h1f6eDS1vrPnSCtAzQ/zg0Lze3FkxKwnp5+wIlORAkiyPXZG+L9pMbnzofc+g
5kFWsqnjziJqDqOPm1++eCVarTvLq03Yi5a6QCcLwtqGPsAkxyRK1CPP/kMJ6eGSsgE+VwEOOcmA
m4ksOeGcFrxpow65ZNmUct4z2MFBpTmOdjqHNZeppVDoWvxtlK7wdjJzKlHaoIpTC746kzB16uxo
0ufIxCrNizr5zRjMMvj52IUFYjYrXcEMebDo5BStLoLAXZwtN31Ep7xWIaCQm+VGm96Zwap46Dwf
Rprd+T/Uphlglg6twBGQEvVShOpP4o/vF+FxcZoC6I6MTquVgs3A5qtk21S4x88zHYYmZxrbBkm8
WumbS01s/L3J5YzTN0USnNhLoCiNPU6eojLanZs55jAnPo/xOBnW2IeZMKqBJfHYkHG4a5/oDSH4
vEDY8Z91ES8syiEdWBZR3u6xkqoIkuFljEuOuQjAJhQgZf0EKK5rHZVMD0IOJsCBnv7vhzTnkSVB
DA3/aDDWTC1ZJMvfIcUFdRWobAENXyVyle7T58boI6VfG2S3EI0fsT6ArBpUHBIURb4R2lirZsPD
bslQWMctMcf2dzijntA39yiKzDlpv2PEnh0JrC+ndwAiHRTSvWxqHa7ggf4TYUdWpkYLXVyDGbTf
FNJPGO2IihLawg+dxSCUXoEX4Txv92tGEUZCTj54YoVrS/7DAi1vcCdUED8D3Brbj5pDWBT76ZvS
iLypf9sqfm2tKwYkobJSgbUMLrxvNYvf82XQx8jj78l9Jpny5m41J+482a3OnoHWMth3u8FdoI0b
YNIiyo+NHihbIzLV9+opmO/eH/fo+HhnJaTP9PRqXochhmJrkYZ9I6BecCePk6xYE+4142v1LPrS
TIMRtvuYy8JXNXYQp/0LX7Mwx1CjExz9vZMlnu0iGEFwZeHwL1KY98sT7jGDLoPhn8lw1vMh0GnQ
8zdxicu/E113J6FKsAB5zT6klAwrLbaxTqaq+M1KZsudernpsduCwWVgEUbhhFxiLqRwuphxBHvV
gTV9J3AXLa25X5SaLEpxjNa7tf4I49VLlJM0Ov+x3Ai8UIz/LyTD9h7uHGsFYfNXdmh/ots93nEM
43Wlq6qmdmrejmp2d+pDDUbrmg1WPRcK/lP6haR5xXy6WLuvevVUNT1gyxY7qcx6iOR76yiUH7w0
SxZaK8GdH8BjKjbRvam0aRMMisIlgIFx1b475Elqsndw8NFrumzMYO3mu4wgjpu9IHvh8ebe31ZD
B/TA/H+Ww8cVqZB8suOzSlYrC6n7wLZtOrSelaLj92rmeMOP8CB9qIOYAqMZAvc6A3FUDxNCtbfD
/srKh63Mf2kzysd3S1oUyzV1C4QqpAu6XbxOuADVtQnsyePOMwkVxntvwylo9XU9IXKl0yGHeqDu
SP9WAEYePODwLA/VEILBmaHwyRNXh0ZSdAcs8uymDgUq5BhJw1AnAO/1RfQREE6OpaVON4DheI92
WHjrfoQAKi4FmtE2jw1+l05qAdkJbHP/O0+boH3c6PLOUbbPPw/qqzlFsXqQz7Ei0j+Yz7Wp2PKp
7s+Qejj0mjM+fZ1Q/gqz5upcfwnFqaqDdYaLB3YeQ4BiIXRefYJuKaAZJaIm+GO8hbeu27ub7UBq
0gOD6zcCKDLK5b8rDqVJkGNfDo4YOcVOav+Uat1jR/fIcQcAqdoBmPAv6NR24gngoPe+PCBVUhVf
3fefZhKBKmAJdhMkDI4mK+1ewCQXscOVEhG02oD+l+frV3JHGzqeCzpfRqs1+nfSbrM6gUlsTqZx
XPw/k0u6Ba4ZH6q3/nUnx8y+g/2ZvpKuNAor464qIS0S5tR0jiA2z7pECMAeoGGj0tPumormGhBW
p9GDYMwcQGExo/0w3Ytv3omk/OITmDu2R6Nst5Yzu81l+BVMBgWAxvpWg6a28zrg7w9Go/eDZ31A
GjnvSQ0EHpY9etwdDwvD6B3imBAeznBY2d+84J+PLHFbG4i8JYpvvctgQN3FU/Ofl5zSLBbwZzM/
Q+AkuuoIfhnBEcpyMDKSlY+gR19Kmue5/HWj+bskaEWcpHME80meHf2O82QUS5HhuAqOilM5x+Ea
0fMZsecM1dc9njTk6sQC/652slQ8pcN4kTKgSX0gbB0xQI7HVOza24g5k1hmCYun8nsBI6RxnqNw
r2VJZ3yBoXhr8r2tD/jE9A+JBE96P6NggDc8Oi0CWqRQPhcODufiHYLZLjOQHbKEh1XGdnRwPLqp
2IdcExjQERG9UK6ANn9BFsjF9B5EJDq2yt+ccB69KJ0KmZ4hWHbk6MOUyb1EU8rOR6a43ZYbJXGJ
wej9LYOuz49OC1817LJCw1UBXJP/Mu84OIQqXF5IR1/XtVpiuP6XwqTMdDBuSc6vMgUUcuLbKl0H
SHPqquoWbfxZDBAcgJ0mIH5vIvKHq18aOddhQAh+BAD2NtVWWXDk0wVeOURp0VDZEPWjRih4Qf4Z
Hmxhh+JWn0riKPzML9Zi4qsIC8jS0qyerImRnZm6XnxLSbxEiIKQkjxHjMM8GQm21DQZ5unGhzuw
4oR/7nVEEe+TT1xtUwCUlEPN1YyQg0oEdiLmTm/49TikZKRtexAynxnsGe3LOcUQx6WEc7XEFI0n
SucK4Y+GRyYCunvZOUfC8KaDgjCtjz0/EvWLIwwXfkBapQe7r6ANrxhakxKAITIOsMDbPNnmjd5M
PRyc3FNr1UIpx9IvFPdmQcDHc2qz0H6j+LnW4hN//YD0qWwAlfyM24SOPXIZdVZh7TeME0aaQ3Eo
QFNdqRcxZIvng55JApHW0M4sc0J3sG/17aFYHJ+pk7OALKqIpl6kCwNp1T9tcpe8BEglY76jgp1y
4VKTjJn8ddVc8KtSSWtx43vqJ59tWhhNcp3+ffAryUXOEEhJR8AGUjWfmShpjFoYkLu9tXfWj9me
U26ypVQXbC8Pg4bcgcBQ63w6f1H/QohfVHE+kvquLUFTx8/U0++7bzNqv6JDiq6cDJGzCF3eTo7Q
FyFdaPARspfZBc8iM6ob+wBMwbobqit+Xv5oAx7NWGPanMAH+xuRkhZz3Ywmm0JXAs6dFTHiwFBV
PpdUgPcbLd9u6zQhOw5PFnjRHotkEk0SDm3ecnp/6Ya/5h2b+9fPIgMVajrMdoPl44Y8yUMeoHCo
KuseGI2OEhzcZRlXfXbcDSfF0EiZxPauJbmQ5qFzZJUHWriJ0cuB8O83RsdWcMTPFRjoMs1JCpY2
TP0o2FRCSxEwqwmxLxDFIz8ao5cdmuig2dHolNvqRBQz6g0TLDhsKP9CfpBfcBZlZ7BPgf3ULQm3
zVGZWV8JTG4Fy29jjL20Wn7PTVrObsA6hAFTyNyS7LRgyQNE9sObW9N2dZHkRyNA/2maZEqmKMbq
iF3mycpodJ8aUHHaDBdwWEIAnFM/OCl5ZIIKgdSEEa2q6pNWvac4j5mYEcdCi/LZyYYofSGUO2FW
FsOlnWEAUGTE+P4CqHZlsBVRbNhCnwdks0Rc9tsX5xEhUDLMinnKptsVum0mFGZV/4clwoUkHpyk
jwFAoNMlrLajbbnWd74YOmgrVVt3zjSNsVhkvwwvT9Ul0+FAWPup1QV5Ha9KiaSEYO3ZVCgiAzMv
9WEuCGL86GSOZei4PyZ5A6rkqYoJqxcn+h6nIhr5Kd2Imy/4TxkecFSxOidtkNokjEVmm9aBJupg
EOYFMdvmLlJXErdjK541GSGOFgx3OLuJ6P1vFp0uv9pT3+LDUevzcJ/oCnZsz+7NUNpxe/02ZMyK
hi3VyAmvwDiaifkXq6RPGZ6r9Yt6Jr9IBh+OzVp3EnMInwRO5TfyqbVWuC8Jfn7YzkahwfbybWMR
UVRql7HyyXqMKhbwiBFmD8HFuCi4LlHM5+viSrs8bdCbd7Frgpf7vGOWgFmBbyXyBMo5Mhpsbgc/
hrB3Lp0J1YkogoZW2iD4BvQdC9ZaM/qYAsJbDgXR+CW6l7iYSX3wn2I4nhSYx/DNqtGExV9uYXq4
zhwpDKaDa6ZGSGwzkJWGjWJ3zusYEF3t3z7S4JstXrPk7LNoNWwMC3ylrxzm4h7iS0yRnVcgfw0E
4ZqRdUxNZGr+79cjpdWv6Tcc0isiZlomUctye0VzMYnE2K4H1MsTIA+eIxqf/jN0B1TEmUoCG9YZ
g/ZDUA5PoKTC51EWNSPJxPXfzCi9CvUPsHa05Zc10dbmBWpzBkIccw3Sh72MsGKmeb9qqzq0h9jn
2hl84lviD9lTxAVuyuc3P24hsRuPpei84SRyKmBOlf1+BBgNCLFSOuSVZHbywjEV3M9igSqY9NLr
pWpK93iZwCMrrMUTHLKApdJMwVeJUE46GwMOMSpFgAykyQu3Nw3vqRHvZpJbvwvjmhRevfZhMgDU
2OguCm8+pMQkKUIuhJf/9jSZXV0fdsVFZ6+d0UMbY3w4vhmbZQGHuWUBrKXuDurlG3KUo8CnLcAK
Zs/wsNPvQoOi2PPtmcEm42QeffAkgsnczvK+aECC7MY/A+x50SF0SuiQm+9XKs2pCER0PHStFKVS
TqM+96mFefDUwm9Az9O9yUkgMMz6a2SpVBTcNLM14/EwqLsbdZeklkp+r+hJvkC/Vr5gBWyoG7L6
JGVn+JoQ7yCaYi4IMZtNN5yCd9x6fQR6AFQVk0S3KXDAxx+ToJA7bw6qQt1WGMpiFaQh3jcXw2sq
gmlZZ8I94RuZWq9+wHvjHsuUPQ7PuJykVQ3do7F0CrkDT0nnkb7BdK7uXpYt6ywHEePM0bp3q3qi
uyzOJZ74boO0SWxIOYGTdZ+NX1lFMwM0LNzvKf5Z3hAaT3R7qzKL9OfRp6LpCZxc9QtxhYdsOlt9
8VoiqAYIZtBEMkj6l/EqgE8prTobeLE6ls3V+NldPGDhnNKZbzsyHTVuUW4DT2V2SBglX+/ePl4U
xeVzmTYbBSxAo6wM+n5dzILFRbXD81cflMB8fOxqVQMjckkroypwAYgUqsxDD/qLx4dLkkjbdtEV
VHWRQKp8Lc8ckLSNyBbJ8+A6exRwxzjF5FPodmBA8n4n89YuBgTZa2rYBnErzg2dyo+pEOJ8btT8
IdMFBWqCwaVuqTlOfaMO/339OnjFtCh9s9jfeLv4C1OB0UunY/XgHgwlFeYWsSS8lnnLd65V/iNw
Cgffrni35so0/qMN7r+BIRNSZW4fDUHK2HwMXr56ONtEBo+LTV052FnQGkTreaWKIe6v7x5J3DkH
ssgOwiuO/PiIOC2THJIsGpS2cwQtPIfsS1Ut1XYrnbeqXNszh/Ed+DHSkB7EIiLuQV/poOsNr38E
tGVp9BGUWAddC4V+jCF4Bm49QVDTIxL9/BiKJA8WCG5Y5kLq9XTOcXZI2qIMyft5Xi+ytmX3VSZi
WiN1cS6kdMwmL3xtN+UhUGxnxE/Dy6eXZFpEjVQyty+v8r/A5bh+2ZmkZ7dHWAsN1gy2dwY7mhCy
zwwWjZK17RA31Ut/xrxwVa1qw/tA3Ipf8OTMruJbh5wrYy8i4Ud/9caQYZn6xmxX1fozXa4Sqf2T
BE/dwbmZJcjQBcDKbLrNrRpzQn9sK3aTMkNWmxf0+dOrFi39tFmawfyeAi6Vi9UcpmdpHyYEFUPa
jeOp7E/k3BRSjNClx5+6EJkdygObrehqBte/SzWLWE55wErfoCFl76UA7YPKjZ0Xzm4ATHw2FANj
e613fYCNZNwR21zFsEdBlXrBg8cgzSmm821AADPloWAnJm4hpX3Lmzeib67vj0/1EWT/PDXshEOj
mInSqF5LNVyZJ/wnMTg5drsxYwURet1Caszc0LVgLhovX5RC/edNV0RN0jeKskOISnNpeE94t8Il
NZRnHGnZFfKY2/jQ7JQIeOYZ5o50ZITHXV38SVphYm3pPOB8HVZlcwBUNrvb0jcpxSW+Tp6iMyNy
0C8vfGrnFqLrz1B3zL8H9GXv2BoMitXWVCg1JBJ/DrvF336OyDLaj6Mn0KsYvEujeD9BkPg8TXy/
VohRYKm1bTN/MqSG0tUlXk+9yOlKfIsM/b7vXx+mQHsSui4efA92sG4tpJ0cVzLFM+RasRyI8xuM
Cr6cFgJQXymVYZ4QqgFYTIPscPXk+5qaUnNEjgut3AtoXvre4mKixArQpVHOAsr+/5j6Cli0c+jj
cvyEz3f/pO4Hk/OLD5PNXp0KPppmxiQwiuNZPY789yIrmX3OFS223vEgcjDpKmnNwDDqFMGOB1LN
9FcZYLc47V8XQApRIS6vG1AMKZgtqeJrsQalnzy3QixcnYdPgea1bU00zO5eW+kQJu9Ktc4fHmA9
VpcnjFAOV4k8Di/0tnjYQN+ndLUOdU8Swf8Wld34MJ075S7LDgOWCqIsE+eEk/rCQFQ7IGqG9m8C
KjOx0eI9gZURWM5Q/gM0vqLRJW0v8tQ+7LyoEte7/TgaKS5rpCdwoG1xJl4SN2fv60pMRE2BsZ12
KjMCXO4Nq1CqiseGWdCYjhrYrePqVErnZIO9yU2XZZYXJxa0GvBENQ05VyjsqygnJC+npLY+BbeN
kpW9cUOcZIjcvyKYnVeIvonT7LTxV6kvog+Ac1mRu2Smc8OhDpBZ7bbUbmU3v3zGDi9rpkYr23Xp
qkqa9xQ9yNKINk5U6/eob41E7DPWfrVHHDX6au4mn/euLKUo2kJL2Xhw7uy4+TURr16Jnzl9mrTf
lqt9pSYiXa7bxuSPQ5smGiayNEM66NB/6g2KUDJ7hVxgAQYEQH5BBESV2LmiIRKY01J8onyGNMeP
XTsxaRLytUL4lUO94Bpbs5SoIRs45Tj4XFyHCaWTD9vH+LOAPRXBkiiVxMYKZApC4NXCA5zsy8G9
KVhSn/bH5hP/xTm/bSZQsJR6Wtz1FVYkdGgmo1DpGiGfLs3ZAGsyIiLWtjxECRGjUnZJBOsq6l9R
5BjQc2zpjzpB/kjpOjk2Eyt6UdrDgiGeNtTstfYtc4GORHXXx3iUOaWoXCHgYCZT5c3a8z7MrE+g
/VrvLf8eoAkMVS34kLfLsySp1uyfQPPpgCZg+YEgTiZx/vnpY/80Atfk4pRrdudjN6ZloCLLtMp4
rvFERsxP7YLB7bJUUPY71+i9qGpS+r+fBTHcY7Eb21kLO23qtJ8N3oJ/Zz343rfMdkmJvOVJEWUV
Dr9ntRmndighX7ZywtO0eCBB4fZeSGfXEuR5C9ajmheJT5Em1jRHyCiB0vzc/28jtBzIakvJkloY
ooA9Tz4o13MuqCXvvaeZCDEaBoqnpfC330D/N3X6EE5ggYlP6MmOf4x6vB7nE4ui7WB0RTF1Wskc
S5PhgyAlS6wj1f4bHXVmKex/EtuVrfUhJ8k4qzP4GijhxfI4pJheeGPgo0vuko79qdAu9viJsVPm
s1+8RNfdLplOg107nUnK6Pjrf73eGLZ+/0nAcVxyOB1J5TwC2/9HdBf+x/vkUHZo6OF//cMvfmFe
tazX7eeCDkw9/wnQp3O1dGhsSc6UFyVutMknRx1T6+ebzrVtHF3fV8fd6pOggh4VeE48VNExeowm
qjdgLoubm0KRlnU9Oa/47sVwzB2yNG9RaML4x1+l4HkY3OTXzFGsJ7AIAOSdHnuhGym8VXcjE5dD
kCRLWd1yyGlyyFGA3PgvJtsqJaCNOXwKsX/TQZZgosnm1ycWEEb8wU5XMxLmwS007Y88eGonymwZ
OJQeSRrBPc6XBG8shccPShBaYp/7qD+OFIZxt5O563nbcmu7TUuwgEeLLWCwqEZeJnFR/GN1l/Sq
EKKox90BbVfJRuJ26ex0k8WtMH8BASuFB7ES+yX/qamqx/J2xJi+8nJp6Pb9BSMwLO8w4HL1AI2u
Ds3gorm2DY0vWiydFHbuHhGeAldlV7J6OV/XTOCSKY4JKgPDrG1Om+ZZT5TRUIGH0KsBhjUWRY61
1NLgj2KdSnxfkYSPBUbMiDJPv2pboYIAGdPHrlDMC10A21wHBYiXKI6xkf/VFL7YjGSp3fWgyFef
FxFjaVcqdkNdjeQr7IralDLla2X6Pj54d37iOJMSg7fkfWMmYJd/ybyiMwCEjNJeLo94OeyjmTjV
4x4Y3gd/bvhJyT7y5vcI7hKkjCUb37omIHBFHsi8EfjuUNYdrzEqBA63rSqrBn7ePlSkf8vwtm3k
6plmOecusSWnPFwVPy2V+yV+cNC3Guuewhhbj5mXG1ufVEXW1H6GxtYtZh1bgBaLyWzpLcqxx7fP
r+VUWnd4Ca2ArXja9mVNrhjEotGJD4GtlwF/WlXpvn32F5Qm9DWmXOkQn0Q+Yf7IeV1rVBKrG0Io
gCVHkq7tJ9tvAo2wPSAKs36/mdZKFe2kcfrwhpV7rzFCOgNcgCpFrPwTCLURcgn9nLHomS3bLR0X
jh3/hUEOPiAmvtu2siOLbU23tYcbtEhHJ0L2JxTULe+kS8s8+NRpRlyP2Ui7em7UF5bvuF9Yzh7Z
WHnkgy0JIjQBiTA/vs6OSmafmVEBY6xowltvBMQ2dOKiD2tfz3LPmebiE4Af+hYz9+5K7PPBafEd
i0WWvLWr77dJr+LFvuBmrRY2fobT4auNz1poAkL7jNnaaxXi14VYQwMXwwMZym/isTr863ZhVk/w
vCmBxVTMoq8x93uT+d2Utt4LkSERLdgLQd4Lv+Hsb5j676UyuH5Hu8Xbyl+BkZpOPu9p/LYJzWlF
4Og7su7ntaiV8tkHzyQJa95bDN08z4vDG4sLZvnFZ9WlNeiiyHlw+TDS9tX1aEB6vHGHO3oK176i
w2szUadg3q1+wGY4Pnpx+KtUxKAAopXFlgPa2TtWNrLVdBmKww7teAu1pfe7wXdPGVwFuq4HfToK
z2oQvt/v1gjjbu7eBJV+BINl2ZfGPes1B5o5u13YUNAvQ6Sy8heVpPZMNOJAwUgUOpdrq+hJOdWY
s1Ucfjh8u2L9K+U/wfYkRZn70ZsSWffvA8P/tu8GpX1xmP9oO6ZX2b254+fopuLa856xTKF/vf0P
HFbztl5Nkt+kWkntyJaiLIGAkDRFiOFDXaLFIogPIt2F+VAScdw6X5GgSoXjR2mL55oCwTcg6X0h
JtF9s+ti9pUtMBhzhUjoBsmEy595fuaXH95noh5TcEGose3zlUxPao0aG3E8pG/a5pv0b/oyjCx6
0cYRBCb7b6XeHQnKW6F08TFX93O13S9vCvzFdp/Dh5EupJRAYDy9Tp+UF93t2L5sn+XQytJ9XWTc
QKVAn0uRrzln9AKMx3rQKON7NQcw5a2U97bAwYZSLXeK0LJP00N/J7MDt/PPlRdNs80a1lQaMcCG
zMH43l42CmWrnwvmZ9GRGFv1kCfdCpcdrghbL5DEuvXyDH1wuyOk8yKH66pXb8BD8E/OGFUaYBAO
s4/oDpEfuf/PlOxrT51wNwrEuOLS4wfZXzkcKysbNNRKlBTOihMDlMkYiuaTjbOoV67Tn5SZIFn+
1gbvCOcmEqDIfa3a7UTJtW7fbD/j776YlqNkQXXjPWY6nZ/2FZ1H0FFwBQcAMH+hAx/ZfVTtb4Fd
GHwNK/5G+Yw6jqaBCc9rJhoCVtJs8NFiq2s4y56glwCNc8o6FtFM2RPFBFMwBF6jdV43yhCplvUI
215xZFRNYfBo1ALWCAvrISiOPk1ibqiwvr2yL+Hx8fH5F1lWx3/kKruIr6OehIjfT2bocojgGhaw
pktPeQvYb5HKuIw8r2M67vArJsz+MUDmnRVkeD68w0oWK+ewqT0j3XsGeVNxnCCKwgquFKH3DEhe
wO4nkFBNp3DP5lCUmtbtrWzAGatqWErgcdjZ5wMLvvn3KL5VY4BpRkY5RTrqBpEim6wzboimJZXV
Veo3EgZjumkolhQI74FyrZiFK1Sk2gy4t6PzS6gx3GQLSrSj/J+YP2HbR2+S4IUJQYivN/KfBm5e
9rpKZ/MLpbPH8pP3ud03CK0KmHI8S+2qdbqYrEWAoZjXAjTBIcPkaXN8s6U8LF7dpzmwGUq58h0R
RVGgkbZKjjhzKwVrXu0rN92LMWa60In7VXVom7QwD8d9s3wPNKwqNxHh6uVtVEfI759M4zURETxW
ykdEz2etRTw1LY+xnddRyIt5vDgfwjiBzjqD6RkauADK0DYxbAEB+wdV0KWBHDwVsQz6nwig3ciC
Pq2uRNLpXeGJOVAZOvm9wHALI2kV3gPJqx8FJaKf0M6u1JJBpnVjA4odjV3Xf5/d42Etl3j0HsQO
xSK778JEbcvzrpOrFHATfI6ZfCEHjK7MdRn2B4sOddLdmgr/geIJ4QWIz9i11VH3YDmLuKTe8g4v
yPZQzMHA+T5/2mSPHkMXsgZ8M91+sl1JGcwgRZ2o5SVJ63n690/RoqLh6ou4+J0msZaz2okGRiBv
KSjCrEzgGNKDnx6jr6oOUyNbYDPY5187BWITL5Aqt3FTA/HF29IVmjgzcKNvHxEK3jbuJC8a86l0
X6oI55/LTpfoHEKPVqq6JsYdHg4aNSNyNyfy9eGulzcirnPf806crIv2S8yO3A9ga3lpgZjayY0t
TefpItomP0GzVrNe7hsSuIzKOMG9cHt3SaxtT8f0N7FF+bdVoJlv04TP85meFVGYuhDQbB1fVvFc
zP6VMgaaUH4q6j1+r8qKyEHeKS+oRXASXRd0O9f8HrgiCgX0bP/ly2bt6wQeHeg5A0e9JII6biRv
kCgfGnVumY0Pj3NoxwsFMWqJyBI2KpqLhASCCFMqhF4sVz8SY0Kg44hpnKi2ctdBSUEoZNmHQ6GJ
6yEVShGME9nqcugY/6rP6X6KSHjn+rml6ruVn6gXJ0zMUsVg3r0Yx5CXGR7Y1F4ZlwVDyEl0mLej
WvIRTdx+hXY5VoQzSSTm94uSzRHBLL90pvILBjQ2sdX8lNm2Vcd2l4AibqggZb7W7zJQh1+Y/a/G
ohe+omoaMXRL1WLzt0BilMDTNm/XG/L/S00G077hicLgChwlIiWhQY41q6afPaNt6mG+4n7Ex9/s
361L23SdlBsnsBOPqL+dmBVqtonBaENkgjKje4LEDyOQHizgcz/G0zH/oSkQnZbQjq2hoqow15GY
qlnBJ3fahYxS6TENHPMatLmmIXibxnLSuGWle8dhZNrl7FPgLbmhV/z5/XWbh0wfuwAfsUaQq/gJ
0MzbnSJkanKCl06hFS53CFySoZwScQ3zQC1UqZY12R1Eln2TiyiFzdBIuRLitHLVUsw/ZmShLcnj
MHZCCz/MGzMICTlh8faMdAIqPqAne5qrgj8Tu+0Qh9JpfcPtkZnyg2vLrO7ZDuprrG8VfQdGX3k9
Y1cNFVQcrrSi9hD9/Icjq2grlgcRLcYP0FRl+bXLYH0ZE74rxMUkq6QKibqUZlEgoe1/eBfr0LDA
RvzTdVelJHDF9uLO9zOKouiqeLHQpfaTumUzY8DXYn1OUBbtSvYCdKy0hnKHlFlHLoM1Ew2A+RLD
vUmMB09fgrSoPwm5v8Q3qwljvl/2oa7fNgULoUzyLUlxdz2EIbHSwgUX2kIYHenYL5v9ZjhKR6YR
Z8wZwWN/P3goL0/rj6vNuxfB2KWpxx//acC0l3UQ8zfyGbYjHUl3d9wdiOympJpnz+c640Bsmx67
jWGSilpmEwGVWwqSPvoWSkjddEAGZSZ8+f5pW8v8JUB3vjD5Wi5xDuEcJKViAl34mEA4N2tqVaOH
bFYz0/UpqraftSbDUbTuGQq37LoFzO88yT40mhLs0DvUKQBvw91z5qMVqnjpfJUGd8cx4+XTOeBW
s+ShDz7Skse+puzlAKTeED1Zn0Ov03T+p5uWY8Mk3dA60FcI/FCaFbU4/U4H+r/4MkUb5vnBKGhs
Xx3tRYXL0CWnegdpMT9QF7SfwkVsotqmLPyw0ZG+N5J/eJGal8Ee9FszVrQhl87SoPrstWTLuMmM
NCZz9J2owahganBC1OR2wPHjS3InXFCnn08gB+V6V5rFWJwdwiys8IKIfJvG925/AqkGeQttZwzD
3PRqYR7+XNVmi+rifQnJcuVaCJTiFE92oGDh3aic/45Fk+IhL+CYtSeUJLO3fFhr56jAqCXfgko0
ddmi5zPHt0VZmKTWpCC66nROC7e4J6bPRIa5B5q6zLtJ2YyvLhxDnL/vsYCwdOaCFRrZIA6VGOuX
aEw7cO4/FlMn5pJHcl2KwAE9LxxLmkQH0/00f5wLQWPtVNGT6D8Tppc9YG8yNTHM7p6LsTsk9i39
8IfYdyiiv2vZUh42hBigDBaFsXaUw151cXiTT/imukJIr8dFTKbGcptPszRaF0NsB30POi6D+Yzp
uSDjJ0fJZrWcXyPWcM1Id+kWSoM0MrLAMf2muM3p6VGXGCTZ71Xjz+ySFz93RZas0pImttOHqq4L
Nhf4UM0m+8rGiER9TBz396BopgHu3xNo/etFTqipYOEVRnrgzDMYrdW1I8JiUCy2zb4IoQy8eTBN
bdLv2spj3N8NjHwKR4QsP9i16JIV2JIj2B0LHJh31Pec04f46R9PmwNgFkZpgRQ/V7Uka1O55FlR
S85v28ABRFny5v1tq/6QuPB4tuSOfHucAhnZgEVsrbBpuKzaH2pDdI8y4q7NZI/Cl3FXE/n0ubc1
llDHShcbo6wjvE7C1KspX9wnudPihaHsYCTh9INft443zIuAj0UVkrL5iGiA+iuiOffavsiduCtj
wEf2vGjOOxafvHLARNyj2ybFZJDTL0K9x4dN0ypWqVqjsfFVoqwFtE4lBAVbKa6H7ozQE1S4zK9p
Wlq+6jcRGl4BzJL+EFhbJHrUxX/b9BMd5CmKFx8FJhh+4F/1CHch12KExpwSTlAkKfwXWtUdn6R2
dZU7orEwNHEZcyUbmZl/c4KFc/0KL4byWBYFBgDqFi42qYO8GveQeQrW2NYmEmvyNYDqSfjnQxgu
wWe5XassLfexpbYmen4XMYyqi/kDDfWIgP6VFlZpKHK2XbJ9ujJ3M2S4jNliyGlacDwvHVnqpgQ4
XrQbakqxq3pGjky5HGKvm/HsiAgFpbduDWLPK+Wxg6Rz/+0PJaJ9f6I8QTqwWFieZJnzUYJWxP1l
CFRUE42B+ovvwD8Jo0Sam1Yzi0Lm83hoqep6HVqrJAybkHiMxjnSjeMBIUlTEZAvbYcJg6NJrzSo
pzjICIZZ08TFS2/qsddDS2zYU2Iw2/59Gwl37pmB26bfiH9qrItd8GhlrBGvGOfCvrljaBX4vh37
1oOjdtxfxKMlEVHRLplQctAADViEcan94dPFr/ew+F/dMpZ+ldzRu8v6fTJ+N66b1VLGAxodvIX3
0hVozHhXmAcFPDTjiDUx2iYAbsk6XH6ri07RPg3l9BOZrM+YxpNH4z/PmoCvta/oLn5aOkqp4OkE
e+OL3MRkh31ufvxwLtutcZExFzTtQhJrVbvV5DZ7VF7Bk7XB3UVkZNaJFaaYPn0WQ9kY1QoI4UKZ
qzDsA/XS86CtZvAnsrInxouN32sqAujQ8rapb0xUSaRkyuCJ39GiSIn3wBL9o31ozqYp+P4OvAFl
TUZOWkDq0oaFoVS5KRV0mtMwyj7MKW7mK47tRiQ40uKGGvZexuYIt+CFaRGWDtatpEzeI0/w4dps
+omx/61ChSKu8LFmk85SeGr25Zoi4THVZIsFPkIRCQml7V4zy0dTotJ+4pAQzwLD5bWgec1Z5aH5
eer18ny/sM4obO6Z8w2XOT5BKeS/TCc3B5RFQBhr91T1C13Qw2XzXapDMThRZPgQqxPpsKedT1VX
my+EgQ86DSFzpulwP70tyxCBsJy6uj12xwCiDVPU8fSvLAKoq2K3LgD2M2Rj1jLXIIxqXTQ3wX5J
6lu4s201V8NhT9n4y1imHLk5oNyifC4nOgqi3hAVykg7xROyeMB0NlwLojn271t7DDR4geJVpHTb
4R9DCu8QAgvSeD19L2F3IvyRxHgQlZw85NRmXY18wrM1seaM+04BsJ3wACrmNWnpQsXnRs/YPh8A
GaOGMMjFhEzh6HT3LjBDy+BKmMrgj/jBhOtEElZYaO4KSZcD3AXinXk26B8Yb0VoI5gxg+c3h6yF
XcaXYNahQ97BcygbD98cr7UzC5V00QXCNz1odMrNMNQ4ODhzhd85qMUbSJYDakvFkyezuEqQBgHb
suYFiDaaP1K4JhroRDzSUuoAExLKsRILGfGzSIxJte9F3sURWIe8/CL8ZXwQ9wUlPvxoCoAOHNLA
qlPLXezXWnZx76xYvMxYplmVwrfTwm+J7acKcuwFzNo4d+VHSxx8MuKtBVA/sH6sVR0e2YrUuiDB
16+/RmByB9huCwLDGZGnfMFiVw0cMS9tRTTWvDnDIWIzS0mWBd8/kTF9+K4mLXDo1cXwZGvcPHLv
uzL6JB1NXjpjNCuTzOcRVtPd8rjh00TyoXqae/Y8bxUZ5PcJvLG4vSY9+8Npn/t20dQMjdS3sNVj
fM6l9ZrxPIsvMVWBA7DYCu1WqdXGZ4lcrh/5tCUcf/5s4H/DugM+QyjSezZw326YPHu573AyhEcl
+AdR2lxqmhuOArdXxmGq5ztMtXqLIk0alasMbBITy+TPEHMbkRj0AzpM/Zq+ATrOEL/5HjZToDti
Q2BNr7bs+xrKptZC0iIM/Moe/irH9JgW3yFAn3DO5snV6V8apoqJMxAqiHJfFdB6qQk/Gxe0WqF7
B7NhoHFexr8IEM/vxiGIADSF2B+G1eW7HHRAorfWH8ZPIt8T0iUWQM6wPelT9ploWEZi/cDe4NE4
BB6QtvdR3FbsH956wlOvesC9LtKEbsixIX+Mu6mNo7pOlSIHvjcLI14v3R04YU94e7wBzpN+Yy6u
+Ko5T9VShNpqY9N7hgcncyM77tot6LO78CsAxfFq+IZqvMn4/K5f8chcZLGSqbIHV/lRajlLHPkU
NjUQXeztUsbqR0Z+PG9j6trVLU9pWbvLq6UQJ2HfIHWRat4+yj9n2qApxkd1HdzRQ8kRuH6YWwai
HOpX6t1u06DGHq3FuhdwA6n3YiRQ1GfeU7DzZlhq6WIkYJTcnNh5pwuTgBGghx9cHH5t86d9Y1K3
ykrsYRCJWTDeSx1UpV9Q3o9EAbTFz+FHG5ipR5Huu7F/bBBySlr3VPBzGvEgoYrg01D5Jw6LCfG/
XlSV2ypYNtX8i7gHNZBC4Wl877YOU/Lu3XI0drHkLb7Uts4i3j6x6C9A6F3d2ARowY+uae/H13mT
irBMDU64lL1oDwzbTxz0uunAdd0SFzrL6f+Yi0Lkqy973m2rrj+xwHA1MPfsG6N1JlDhu0OL8l4U
4vZUoei0Tp1nDxUW6WDoG9jfQ/tQ9BMb4/ub1Hwft6DypZrxZUmIknxTM9TwpN+LJHwAx/nroi7r
qc0OPS+uXhwxOF10oOQDHjb/4k5tC/WN4/hTtxBz5V3uKYBrE846BWmK6VONNJMYXbZn3q9LuPX+
2LDiRRlmDDYibAyRcSi1fg1v/nY8I9Ij4cs2gD6i/Q87xEBMUUMTzMVQVZVIF7kUgB+dt+Z+lrQu
++Pf/hHH8r+nKsFrDlPnFcCJfYMPB5IEOdNAnL/IO5PXKy+fOIV+SIOVzXK9HDv/1+7C4f1qJYfv
LvqwuRK2FjDywUR8WUpL9NZT+GR2vtoRwdZusVI9JqLVQ8pGLAaIqQpuhhYz/xAzk138se8SNZ2p
uiyylAJrfs2LHF0k+iDyRyocsL8iJdBpHRLCIyOgboQXUqpy3JtMXT0UPkhevmduXBzjfsMe3aLI
Dw9ppQKMMjPnFVsRT3ZJHbGtPyBqx9RvIe0MY1yKwFI9Xk9zzslOqgCPhcj+iNiMOzDm4icxFWN0
c5fqyKGyPrJPFLgxSg4DPMFYxr7Hu1b8OCWrUAfOqad0f9RMoKfvU+T85QfVMRClGrAb+BAo3Le4
FyyaVvfZj5R1FZ5SGakAYGDmNtTuL4PAIhgWPUf89YGdbl+7ilrkyJPSGNtQ1BE99vOQG59svPcr
iH3o9PG811vMpspmBK1RFVgtniR+axztBE+1baNvKp5lPjKfMPyCPiY5li7tJe28M3WUOzP94Vpk
188iE5gkiwOc5/okNUcNassSbalZ8eMJgaZuntCJUPIHNS8i/ruZxqDuky3oRHO+i9QqzKHDjvCc
HhZJhDza/mdxO8rKAczQNgT1r1sR9baTfMvTcKszo8iw6hQ0yIhAsy0P9BCc5qgb12JD6L95HGRS
dENba6tHy+AAjA3E+uHWUkyQ7XK/TdYCt2G+a0B7c1MBQiTT62hr0JVphKC7Pb9V74MKT+jBPEZp
3Rppv7GqjgtjiCK3jXJIfpR80ifacgL2cZeDRdab9bnIT65TJonsg97ojLgVbZnenkFkZsPe7P3V
OX9DL0LFwl/gDsWLcCJ2ydSLqcOoo3uFEdrxNLs3aLw3jjwDQXwPKfy1PBsfxcbwHjParWA86RZ8
/HilQLrE6OBuQt6+5vnO+ss6PSrn5gUSXydV1UWxjEM8fKmOZQSjqL+7cR0RSXOccwxHEGp0BnFK
kihEvJL55qiEhOljCASBTnwQkHoQBhmdtwLkO22hkiky0mI3NW/jsakfyFE0nysNJHXEMMGNvIfw
KV2RLp8F86B5Q0zKATYGs1FLB8p/FifBWNJ2lbWjE4mIlfnoUSX2tpz2zD8Jvole0fUih60xaBLd
uGY42ToH1PciCKr97Hy4huPjDbVQ4vwx37JPwhBko+v+FqU9DQw9p+oKLrwtQoOpHWM9kXmZAy81
UDrtsa0TCDKRt/XwuTBs8ff5adtN/iCWVnnNgkPca00kD1BAZeQNbrpyLR2r2scGDZtxrnP2pqF6
Ago/Dn/v9X92xctGAoIONE+yJmn5jRmUDVYoHQ6ENPllQQXzVIym0J4W/k4dlhF9fK0LPNEN+ZQF
jVunCiuO1OxTQz7tHruNhAEdFJ0GYEgkMpHPu7RXHk6+UudfJrFRWeCTlnQrd1QbStAGWSy9tPSl
FL5uomr9+13oLmYXm37W1/9JIa9XTm8UH/HhyscOpfK2odcbqh2G1urMHUTdRMlCLr3rzmqILa0f
vydyc0zuAkUV62rSW11cyGyOIcIgjKuT7agfbjd9YP3vJGmTZrVeLrY7seuY7gW9b/7i6TvvJI/7
PusUT4wugdPJYo1gXhF4+g2AYAAxsNOIB61OIDIz/xosmQ5pqmW327BBDQ7bTmxgDRj+Ff6mrBW6
Xerh3LtEOtNKYCIamZ7nSrLlma6i2myNmaVlh20wDU+TqUdO8rrGiOvvqPc0QkKqzv95+rLSFhA2
b/+iJNihSzeDAOTzGRi6bijBp6gv/mMmM/NMH/cxWf49Q1Lgs1BrbHTIRbVNVyu2OLrZnhTUtrxm
xmTTaWXGG+Yv+GUBQVUfFK6mXc7HLU+Zrz6YGUC8cVat0DJ70NHHCh21zfPtQcP+VtMJaR3k+tPC
WkT9Gffp4BBCgLi8urzh0A3mZNNiol0oGQdlRFva8iYV46AHqSZJ1MTVWoHygig8EjKWvoFB0rXS
Op0smVgFIQbQ634wfUP1BnCaS6F/MMPunAmASdaYkELPaWQced6qtoIra3s4GaW3NG6WDCrd43NP
Q/JhOCefnomI8s15HsqgpW8SuJ4NWgNvhKcxoSVBJlNCQxoZWq5h7R7Y2uCsZdDTwfq3qS+lclej
Exn5f8MnIvWDHrzcjmP5Y4k7W/OoILNU5FZ4fdX7Jf/p7+Q+cDv/ieY8DUvyY55rH10nvnkmeOac
S8dD30psPgAQFhgq5tXEONPp8AALk5JMZEkECD47PGojCpnEcvVvo3KJvpBwOKTDLnZXAmyP/u/R
lvdS3qe52ZP0nXi/QyuYNe0NQxgqhjLmONyA3WfnWERQ/HM9NDzR39zEsv6uLJOuvYcfq/31byTR
ft+pg46QjBavgkvsmjwrNZpzrB2jKfCUK7jwN11H3iXrK/gyZVov0jveEcYaCFcSz2CH8Xb3X0J6
GoWucTksabtag6blEMwmE5K9PUfrQ2Wqw8EVyUkPhXo39vLNzuxxN+4lyxjneU1osNbI2lvJ4+pF
ERphp4brbHeEk4KqMUiSUXkXGPzqpuG7Q1mnNXmRpmw1maEpgz7Xrk6guVnphH+owWTGRENm9cyG
RyO3qsuV/xRsGRswnUcfKsSllnvsdOs+xQ1D27qABrPFH8b0lw4+n9Dyy8b85rhAUIUNrGPbBxk8
q6yffAEvhGFNpowM+JdA8C8pUVXlwXnwuJwlAPa13L8NqHspvtkExrMrRq1xAxMT9Qm9P1fFIcAH
rhE4PkJZtog4iHBSG67IgH7gCBV8jQI9kfzSiF/mDYA1lm/Z0G7D36GVh/jqPj80/Tis6JFEZb8Z
gYgzUwzXuieQxkCpDnBoseJNn/iKZMQg2vvwfCg9dAA/TWFEeNUi8K8jIaEjEJuUxVU/xKSfr6QI
bcvsrKaEcYHKvGp1Ph+OXMP8DBBKKhKs3YS9VjZcMOZwZtnQIW95rFiLKsVmwyGBtTdAh7s9y705
NNAPVVcfHxLCQtKFuXvE1qB6HpkWqhl9hmTOgDmczXOwY9ClCLLtLLj6/y3mZVhlaMsFSjkNSBxJ
zZUFX9NNhxNVN1jDdjECbyLf3WJC0maz4rfZXoMPVvjEF33GLbqXd/Fbj9Wqq0e95EMLCfHabR3W
aswGIw83WNnCL1mhj/iwgG4FZeuJdnTgqpoQMcYW24Wa5HWeO3dH93YiwIUgQ41g6VUbBywccRxV
2MOsAb1Ewf3Xl9N9cgRB3341yhjwxTaJu0YFO5QFM5r9nN6M+0AvaQG3R9TBgwx9Ixyhj9jU68U2
nnybkgePwQV2JYNpkbHmOmgJfthn2ot7/wQOyeZNpaXZAdYYBDuk8x18g+KEKVwq0/0wPHkt4b13
Ft7f2tUEuAUhg21jaerw8kK6fMi76cpsCco4+Dntk1nE3/MMnZU4DN9OlRb3lbIjEpMZioavuORn
BEpuriNepYbeZarUTjvdMAttHInGhoMEPMuwW9qCP3ZFIEbCFQ0DJFnpXD4fWucOZ+dev7mOKYn4
IJpPAUxFXV5D5XMVr2vGexypKTjnGLzO/Lo05IkUCRwf0Xminfr11NRXTmnKKGKPT/Sr4rE14xKC
BHNXyjIGPt09wbxISj2+fdHPSfAqdZN+pOKjRiORE2OOgZtkdZEKklubVNbPpFZhsSv7xa1yEl5O
jF0eEDqLA//mmVdjAwlKqHiFF5Kxgdcdu3URTN6Lu0Ql9FeTiBE58O+SxVGL2kVhUW2DCUk6yiKB
CkTlBOdqGv5HFT/XQe5TEfyDUux4BlGNDswElly1pXpeRCzyJ1RpGO1pdkwzGi/tbMU8Q+dkBAH7
Ku0r7i8DHwke3dJ0Q1tGwVBdrvo+ECr61PbeX9tYtMKBBhMTVxpSFTBzIRWFVLIzaCs6fJzYkULP
SEt8Aotx+Y5O0GDjmWfFv4NL3AJhZyxpkUIKD27//JrqCiDq6wRtMmE9K5CpPHsIi95cDNB+9qwM
liYEc725vdllJmgKsdyML2rGnLweEPeUgC73HCgB/TCY6tVmxwkWThCPM7WiTjzBjBU+EizI5AgK
VWjJLYiYBmN3hbNRsWbShuVLlm9gRo4FkB/90rQVJ7tr6sTk6NoTGZJu6p9ZYYqbQMCx3MS6PIWd
2fNSyptfzdEiWpqSOvzTQb3iHTikgxw7Oe3akhGNn4v4IbGkgrpQVxCr5Rn2nlov19at0bprAf7t
8x/l+SmjmDJquuxvZMhgfGLPISwTQAG5NHn9wyBFpBqtel52AezaHMgJjIkxWxAZ17Yp63k0Kmmd
B/le9sDXYly3A9ycqz69ueYM+Qpg6BIbkpttbbgWGEHn/2Azv1sWPO2T7PvyLNlAV8IaqwBDF8sQ
++wbczMgqDVyo7mRq3AdDCvtjhDxZIkjlxKL1FDGqRbwTwNJV5ikfvDl8O2rjw1os9XCs4RPceUF
y/oWVw6Vt3ypf39G299vkOnSRq1mcxza592oMA0rZMeXnhjOLKJJHAaMXg+DMwvAGwQMW6KZTc6s
r7qObFcTYoiAToGD4a14qG8ciQFxTmbZtUeG5j7qyLx2cbTTG7ZklyiYZufPtP0P41+rAz19F7hj
NqewnVwefY+PLX468YoeeBbXGifSiQyfoXeOmGkJZy6e6D9xSz9WQu1Ceo7c7FhsbnLHV1XTMIpR
jDVQ1KIpBecDFNUojaoodBrEFkbnlEjrpmr+V0ngGjRKbLioW8G0RxLyuc0US3Mu/PZ5Zq2UHcwY
lNvY9KUfiN77nx+m36+eTR6h9kQXTmYaqxOC0ILGSFJECMruYAQG/UDPQRmSR5YXZZ0yNxbMBgAB
kJ2hI155zzPfxuiNX+YxoEPOi4H4brcZliq1bSMrUir7ynNI09kTruLCnQ8Lv9Wm+QXtgIh9/QSq
gjDyrySD94Bf8brVL2fenHIlJOoFrgJhYd6azVTLIm2Dm8zVeHpz12EL/6SdI3C8jOp2MqPiiZdP
36jAx0oxnAvtE8bDRn8QvcCQFpjimjdyfCpwXutqDyYk+paI70bpKMoBPLDVM2R93pmwgQo1hK9u
Cv2PDKYAlUZ5ZgC8RDoE9i4WIjJzS3hC7V09cmRBhLrGU6Ae88jmnORG7SOHbyEXSl54klFeno2K
puHzBn+rY24yXDs1gT1/pwfnguZFjNItXyXUOWcdUceq4jkZYw1RCFpYGmkAIp5vSv12s/G9KZfp
nUrWM2RQP2dRpXM6uRUtlapD9nbx99S/1FQ5SdnHNygHZOZua7ZJG6NZ9DdI0K/A0ZaN5Xf5DDkc
YyQOZRn22fDQWqtVgp7XM2gm5vpTBnsXJrqX71EK2en2atTBRG3WuERmXU0zvq0JSaig/oMbcbhQ
l4ZyRUp8EWFLOlIhk3fZ9yVCfBN/vShEHBrXqlAPdipqMIT6GbNcQQPA5ga26k6wHJSg9E0dhs80
hlGmR38Aov56s3dEjT6Bp6hZrHYLDuH6Kz6bKk7nHjHbnfBXiX2Kw3GJIgepilyKED0rXzRMRRkg
FecmhWRC/whYCK1QyLz0nM03U6laKfTfGYINEGDckfRwUsj0VwwdBpfZXUf3ZRhKT2LCTgfbqv3B
UPgFrQOu/oiujXow3WFdVe4SKG3AivpQlppFGdUDnKoRNSPQfBdrG6KWtPQmkCZzH+65m6Y/58v7
/2I0Jp3/8m0/nv7dY9KcjyPAN+GqCgPrkT5GbJvoqrbiM2zCsGvGU+AqmZvQ8Nk2SUFqvDj0xyUn
LiX/CuWcF0l15yv7VfbC2i1M4eUFrIbm+fXMySLN36/66Bch73c0xwTcVJirY0Wc+Ok3XmklR204
r3O1P1OwrSiNf9gIhDDoU+9MbwH1iZm6KSD1SA2ChSrPVR2Ar3v3WISN/gDPEKkVFiHCia31hYQ7
Ix4fRPDlkRJ8jg0yj0BRr3drdpC7I+PINmt+UirS8mhkb1qY9j1SghRpI0p8hEpQG3/AMVZes2HY
AAwX3JuWbJny8RJFcYYnMZkheEOBVrWlqC+Ijf5Yr18p7LJuJdE1YQa1lh6MDr6CoaA35Ky2Jx8L
RRnWHsCHa4Ouv1gVvsyXR2qep9KefcnuI0O3lzZLMm6iTQ6g8XUc8Odg6D3ZA3ggiQwaTZe6TmcW
7yxb13rSWKv3V9tRnZopWxMLnmHwTI74PRoLhayuHfaTX4qp7N7jVWu6aEnocGfpoS8f+8UVoYYL
mTSD4QNKnQPfUXO9hc0wclKJTtFrkJ7WNhiuobN5ZQi5aUKEKHq9dXgXLCk9SYRP+xWWnLiywlvE
dsZkkMPuYm+pD12me8iMOsmYnpTHjsRM51qVflkOYNlKAzmCYUqcGFUiNz1tz2pL1hcGEHaUlZjJ
kfvAFcbNDP8lEgdpJ92sRlK+Ih4hBzOkldkX+U9AjjPRwJo+nHpdngHmEkmiSANP/csRxTu08w03
lka+5xiORE1fi4N0F5sogbGkiq31ZohvU6xe0dBolyb8wsc20Qe+kEHdPqOMUxKFs4GPXK1WC5dE
mhw64N1VFAOmv2eoUN1pDAcTggYFWZimHftGt3PGpf9wM85wqJa47XCMwsxNkmkW5wEgt5+eaoGB
ohpkEqKvuSeho/kLWugPn92cWAipOw8aDaNRTctl+wKngYCQwocvwtb+yMylJPovrxtLmSkGe7eq
Z9qKqUja1lQCN6vBQFnatDPB0UoSW8whTYrIp8VY3dqVl4soRkCNarFgMDWeuFqNG1wdx/jNepn/
I5yBCcNMHdFZza2WzK4pc+dbhyq41zCDuVTMdfbSPWrzQfTMtKfbr++UoQRsjsb6eEjRyjxu2oaa
9xFC/obEwjninnw17PUflxQItXRgmEZfGlWrTEOOh5Z1yBxvsBjftVZipLhx3HTvx+Bvhqwd0cd5
A8oHxXidSqPfDm+FDf9kvDG8ehAEbIMAgrz5pibLSfvNzJ+DbcFwWiYGnkq6R1hzrNNtBaSPnlgG
X2vsdWbZ6Oyya9gfx2CG9VDmxirUmymp2BCbeaEQRwcDxGJZI8q0f+mwF7Mlbsd4vrN5Metnt7+W
2HLlQwYfjhoZU+4xoQUxmUy4qwcLPuext744n6Hpv2h2UoBQsJm+SOKxkB81DBaZHE/hqy9ruWoz
3eiVI7mqQF97rBl5h/yj7UcekTYs9z8jGUCGxjEE+yIzTunqyaO5RIQyAZYiVF9lupFymjGuXLTm
6dFLHAmRVyW/Bg7Pl5Slry0VrWbEyv4v6VBZa6IMb77igyO2l1xUx6Om+mhQrn2r6F6DfHJR6n09
FO7MbMSDWXo4WZI5RBQA053rG0J8Qps+aF06xFj8DSVPsk/p0VdVNtBgRp0YsxoVjSmpuWqGmtHJ
/gHBPOW4qo6L/KSz1N60yhfDzfO5ePjDMTc5VUvSoogdYABVWOCbcaNz59OjN2+WGoaZ/xWo/hOa
n937uYIZo+vHJx9TSYCEm01G8IlxSWnjOGC6fIiMB3+C2kMhZN+WSsijRRXK/dh3USLZeQdjYcZc
L6cEfNIjbtxx8jLOf9kpE4K7Bk1LRswjVg57CKEP29nPCOAzzN9haC5t5t+1paUhwQgciBLS9DlA
TlNykvgCNOmHHwYMjQtgn3Jb3lA4TVdYinOONPnbHSrsw6k/9lbZMHQDWFRm0Qe+vIE2OC8iJj+0
4LFAD45/daSAPrG3xVfRXbYX0GIgmPAD2fXkcy9qHETS9TAezM52NVF6eB8SB94YrGbDgkppPYJj
/xSstllu6MWY1VVQ6gY5ZtPAhzGI+iK/hzckn6Cldn1qLQrUEyhimTOVEpEfVuF150jWAvbpP1Td
3sRaysdHsPU8hvW2ncnKbxZ/0fQMmgo6rsmO3w/SYBE1cd4V+NNduFbHtRhTMPPSIyBZU+KFqzn/
mUMXtCAPaqGmGvMw2pP9/2Zmjbcq5wYt0thtHfymktEdgm+FmK2qrbmmnBCJ16WWhHs4kgJV3N0H
6jFSd5wEisOHAqWORpUy/35J/wYQyP0Aly1DHEMWXfvzVV7Kct0Rb2ohjmU39S6eom12ne04VFIf
6FELSyXX2OzRg6/OZKP3Y/Clg1aXDqfhRvWJ3IBaZmYpv9Q925VXSUi5LswgMN+SNrAuw+ACsmIX
JQ1BXUp3UkttjZgh/pHDg24YLwVLnoq94w7AMZxqw3NkqVzLhcAO6yDy1FbQVeTVMIehPFGq0nu2
nHlW0+eOPoRt15S7iXLYyVPE6m+PQN2tNcqxo6fEwo0FRL8irwtRYH/Iygf0EDe/6BD3oKScpM1r
A7nqDEIWl/2z1cvL3K+wgkejTMPAxrjDR7Q6wGYlBJl+nPNVdR0cxxZ0mg47NBtP4VjM0ZWdpDh4
hnq8tv1Knc1VdmjlaKGfAoDtMffLdkAe3W1fwRb9X+c18uO1BtXIS6t1J4ToGgNudQ5FkDhzxqsH
0gTBNne6xk3La8PI/n1cac95i5JDHRtDZONg9wEvofBP0GrFxo6igkiRCAzlA4d1+rSsZLHnhErJ
ZpRz+GEOnUzF1pIcL/8tC9LT6v+Gxi0ZmvXL5Mj+duznQoh71jeFaS27oT9mTj76j94ZnJb+kzqk
lZq2A7YxkuHzOPBuXT+Kng3EH9bWrYzGp4uTe75dcHnn/nLo2DXnlWX5Qf3te+mVFPDHEhljTYND
iAofbRD2yAdvhX50irFv71ST6W5VITOAth2f/biLY9AE/7qLYkeAtYdiWo/SETpYGm+gmsZeUyPX
EjMioKGaHTgBLWb9j4T0hK9Fh0dQiltDbx24wKktgnZEyi7Vvkq8I5FQHSmG2J6jyztad/JYY9pw
ojQ/wjljWT+WI11yrFpu4uIr1rqgo7wEgY28K9MuuInwUq9dN74cRWyU/fSkj7awkyghTzldrorx
Hj1DAR178Sbz+pkcusYIXusifSO9skf9v2JHABn2QtWSzYZIAA6usx2x1vfwls2qF9RY4+YnFelb
U4ZqqCy96TVzqQM+slee177aHB+7W7aCJDf66OFIRSA6dAGcxYvho/U4NdTW4XMWkEoJAGEidD3P
ccoCUflNW0keUs6/WCDtMh+xneyB5v1iBEeGF8KQFK5FmmhgWMT6YSeL+1sEFQ8X7ysZdr+Yl6th
fp2r3bSuoFosfzzMK4EhI2n9BIgGItZmcX6TIh7G08qhizQHWxj05y7DR1cYIMIgRh3hJ1+6WgN8
SPacoQSLxOaHx94luYfUhJoN3+Pm3rct6/ntUFdJVZGPztZzMojYRaSHc5/ZrClrqzuoo4T+yedu
9VTDUVJtLVqRTxHZuuwYWjia/C/vSD/LDtfrtlrcIfvs57Uyj2e1LjQ80GOksqQtSBI9CjpUS2DY
mbkH/EfQZfx3e9D3s2/aFdu4t5PrHv6hRdoZAQHib1bWA6jiJjAq6OV3JQYjNsUj0flgjXxiL4NZ
maQicFB/CGlSVA4e453MwjP+IqiIlopTbIqPh0MDtvfBbkhgWO+VjLukpc5liMXWh3wyUg6U0PpI
vtZR2Q1CRg6emYWphU00is9S2aSGx/KHtl2CbuGwTNM/Q+2P63jgDl6Np14pW9UoxVzUNG7asH2b
Jscs+9H6SDf4su8D9h5RQ1LUDrNmhT9T8sjmoDcnU6lYoedmm9ZrONbEQK3T98Ymg9Xe2s6zm7J7
I6m7kDj61r/qB52Xp5rfs4nqbaRXLgD2FlEn6MxYSOwsxmfxoVkQitiDQGaQNxyXsHn0wXjiuUvD
i57glvxn4TdoqH1nEt5Q2rE0bH1zLEM9AjzWsYHNZHvqPeK0u44SmTcSKpnYPsMuA5L7JXeMNckp
pkbtrgxIRW2ZXUtRIIkqPDg5hEJPq1fjhEtW0Rbmj9g8EaXNFCREzO2VNGKWxt7E6g5bqHBOpL+Z
Ip80zUwZa4Sq0gdQLi3ZlVtifGSTZ/uWCd2YYjXMw2W64NsBQV4GhGlHtH4ks8V45QH8X3BHMlmp
drsetkK4jE6bz4aFvJvAzgsMYa4d+QQZWjNpC+v7g4Cw2cUZNzAO5zzsWLMRUn2+jEXlUr07z6Lp
9hSxSt4WS6lfN5nV/BO4nr2e8sLAnmGlTKjBvWdnCYBld2BJRveVrzB5dY8lgAGVkn7IIDmxu1xB
G39KT09xCv11mqS0qhYuB6VwUaA487gdOY4pEvXkNSQGy83z/mY5qplAF2ydSgakmi/AsR/xJm09
Visqel6qRkgyVJOU5k4YDJ1KPRe8+GsMy9vhGlcUcIEsQ64IR/JZJHt2Y5bDaqe/wj0C36iPcRtw
ESedGsMmbVYTUOxyDXHG+tjWvYd1vvFoy3DfCYC9111vczwsDHjhyQAYT/xzd0xbrTLfAVL94eGJ
bNn98fdDuwufF+kyVCQxsTEG8F7QVlAL4JxpRpK0PCjMUzVU/Pu5iTzolAYzBkRV9F8QMrNja6sd
XyejgMgq4YA2XY1pAujjAo8Ums2R2txtYFK3qWRk6pX1QDf/xgrvAD/SXyuJtMrHJatwV+eG82bx
aVB1apijobg1CHT2pqMw3biqt2PzyLtTV6iillLOL5IX9bp+/Q/BkQWAJ44BOsp/wfuz3BtgF7NC
TIcqEoS/ilixhck7JqIboDekltI3um7B9+w1lZR49envFzvskB0Z+nKPrfCSRB1m5FogQAmt3xgg
/Ag+sWIEUOly5Sy6e29IoYF24+VUB5mWNEo+TEi4RikBW2+ix36kGoduqC4xYIfWpU0wYM8kcfhS
/IujKhWEsxYZlEppyqm4eHXwrv1QgDVwCg3Xi2/lum5GM1+UpIt2LPtZRpoluHa+RSr5qPHMI9J3
EpbVmu4qCTn9pNyTrQX99M83p87XgymtfwQP3gk8inpsetvRRO6nVjKBOm95YUgkMPrzRZy8IB0z
5nEBGwksoW13BDwJh6dYFbKi7Lmz77e7gCbxuPji8U3lly40k8ONuc1QNCJFUxHPqJY3fb17H9oo
xqGJLwHMHe5ySDFw7h9vDcHqQx+Fvrsb0JZU9nZArn0bcK+k700OeeilwWJUZK+BrmI8DCfPb8vH
cgt4ixJr47c4JwMmc7dgVAbcT2ygbcmu8oGDvNgdR6KTcUxR6j6vKNSSxFaBCBf4OYf7IxKqbsJ8
fCg8M6MQ9IU1TR76C4rtfD1Ou4e46eVUAuDSRz9sxu3thuD180YzAVf3uxxd3RVDRg6HruI60kyE
/JQGHMgi8ZmkuyosfGGDxcSZiHBtdwaiayh4jwG0edj8Uc7G7j1XIuF7Lrn4W4nV2VVM4hEkKBqy
u4W+n39MuPqf4x5jMjdEVJDJMbWLuytHeEo1NaEn8fFFiIVy+voC36FiBDfDz1SFn02iThRUwWgP
shZEbFoE+B801tpT6m7EJq+mtOzTYaJxWuzA6HudrMo+GEPVWHAkR95c5JYSxF3+kPttTRNy0M3u
1u++AgrU+x8ez3v2ZYQ8Q9uGA3KY4U+anLs6bSrjv3H5hZ4R181VKT9Z79DhNHdFvqgX2+pAsHKB
f3dmiYTEc9CYgEAPtRLGYr657KjR3sfx15GTBKT2Uvng2ukHvowUkLCH3qSYfWqBPHc65ey1HDaC
ui9Q6MhdZMOcK1bDm7377u7Q0i8DnFjMxvxhgShc/sbDSNWUIzbcuUq+MAJZUFHZ/F3M9R8C3ADL
pI19b+1T9tUhzr787JuiyaU22nOpjQJDPMXRHJAJVJBvqznbDQqHUULumPpc7REMtr1plhdBcYPQ
X4JbIYqU8sC6FbTJG3zbRz/boe2sqXaCZz0HfiJnjW2PtegROvT9CiogcQAjD4scWzdT4dFROZbV
4EUDzEguugZcqrnu+QoPiavL/ASG92pbhUweiWevSlCK2oh/FzXhBLhNO8EGfT03RaGLaqc5JtHl
sVpM2zpDrwiJh+Kw4KZ0YTxRRIehAF3ERaMypZ7qYNSJswyj3nBmb8sWxSxmEZgPVwU4GAYnhLCT
zyUFTHvX5wIeqk85LA6X77s3AB3VPy8qvXaJUatqWS/+t0UrHm07o1zzR7JPmLZGU7paVlQuWGsw
wgtDqpT4yuQvj3C/9MXmOzZ8WFJr4eRjO0OX/HSi6rrr5oe09xJONN+Xlwoh848K5MD/Or/J1Ujh
LuHc8yGmVNcBsBk+liXGHFNXsX/roAQxUKcfa9jnl6mSvCSd0tRlSyNMQkOdv+m3U+P+d8hFg49X
yljwhPiLklYOinjMd2lPiF8SOvGvLCktnTFxXzBNQFjZg5804Sbb6s+GEi3occIN6aR/DrpGpI0Z
TSqQ5YT8OsfR32/L0pVQFXp1/1MKQV7lZG+fEyMn/VOjfC8dOJ104sAvkAlG3K0/xY52/RFP8RAI
cOwzBKd6uemHN4ZVUi49bGqc8yFEC21YAD23dstf/cESSg6LBq/1dhnBCg3ioUeKM6sBAWIx64U2
nH83uNXmE39tkhSu+huhNujNFz/easiq2cdzYhKJWZNUbxJUQehVNvpYe77L9DWFiSZjhlZfmkQF
cDyyj2U8lgZ/gXrpHJC+vmZtnbZ/vNTzyZsMPYUfw8vl7yy5WRrijUVdG4qger2xJRUZLS1cUI2U
OuuseML912tsCmkZD9MTVhQeG02ufUZCi0AQENGQM+Gt5jJ/HBAeckGzFG4FUySQwx9QzRg7rxSd
QimzPf+8G6jor7BxiRF4LnUwdlj79mFu2eMb5S15T5GU6I4Sg59teGWfNPc92Nqo7u2ixFNTq3VN
2nsJCR9c8sYqjUoD9stVNxd+DKalgFHwy7O7zrnAt6c1h2jWtV3a+As6xwf2qCQ6xlzA2jabJlWr
78N8KTD4h+T+k8FbLpUoKHWvBUhWsIt4XvtbMi5Wu7t6sW9V+X7B6aiYblcQSOxDA+vQtYTz0YpH
8E6WWn4f8NOuaYshAIBUOd8W0lIbcn9IQHn4qhkPYQg471kZtd4dsKeSmiQrd7wBwAROA7qx+yJR
P0+wAk2eb+Bv5XPkTJaA40SFvsCc0ROb0w6zUi7zbX2Rj59vFG5ZuBMgsj4xYP7J6w6tgR1nUrs0
mu7GK3h5d2Q+HMyhQA+7wrt3NLRmNbZwgu1597hubzpt2YVjJdRpcM7MhrmjOiUSqHWoE5+GAXAH
juHAWliPO3uy8lT0/jEiiVfT5b+mcZJaVcHorfFQaibnFE+eyP8QV/p2LoJUMvEZ3Q8PPZf7cxj7
haOEDeyjpz826d4qR3VTUPbFnQqh8TcoYWepCYTHMeBeQpyKfxl3VgkqcOcFZgT5XQvVJ7EnNls8
wHYfVguvfTb6+e17wPiSjrHWcBKab8A6WfPeZIl2IR05LwPzH5d14jQfgb/F6sz6kyEdMfqLDoSz
uZePJ5V5L8ogvC9yy5DZmHU2jkKdP3TgUquCsfJA70VeR2LF/iAEki7Yiq0nvImUciA09GrqCbVN
sL0Zj5AH1qNMrPjofKJP29cMfb0uVODpgozpcjNJWmuEuQvYf6bEHxyK39sYUUB6KX9PuSnpLjpp
BusZdhyBtdVxCydDrrHR+E/jzK8BCqOnEUeY/HVE2WXTveYEB6NOfqZv0vVVixesnaEXtN87RQZC
Qp7Xkq6PU5rsq0TJ92lIZNe3G7f1eLMhv/Yu7MzYmgcHgi/gUb4Je79JxrKdftYjvCzUN8FHyh21
wv0gI0aIjU1ckXfKbtXwQoIuvEOBcDO2hPebyZZgd7Hqv1eQYizfI8ELJg0aeKPfr0d/rWsHSpu7
EPt/Fwlot/XkAWkpYLZldIGhDx/dEA+89hPfOqpeVv5Ef+PMMTHYLCbEq9ErngHDjlKSEzo4OlNs
+GSeE9WX8L3uOocsJxlxmibyydFBQtMwBjodhSoe1cRWgk+yhfJJOg6iesLNyOMJ/+SkmltI5qzp
f5/9htyyUrbJ/yxGYErVCGa3/ZZvsUhCQv8+ocZeOSZaz+68ENuRhC/9EjxHOS5ovEc0FTiS4Hze
/+OxHHsdNXUwFegfq+5S2Qfk7bKRhwIzYWNPibMlXb7fks9lIiGbcNS0ID/pRLIS8CU0HQ2rFGI1
PStTuAahu0zc9XARxJfJU8s88kiQm5QRk0iFrf3jVw0Gp8R0PaJSmJB5D+DoQOer4Lfl0tfzbD9m
dG8746kbWBkq31YUscYfC3f/z8aBOJ0knz6d67V6LwO79ayW3YN0wgrZye81cIPZfDn50BvflP3k
spMfuO6EDbkiE3+5ISgB5S/q8+2qwGo3898C0L+pMGkvHT57Hug2a5r20JEINdIGseNJneRDak/3
aAK8m8fvEMIaiilaDRtGWTPeUfMXpbqhNnl/zycKfPT9wLKBl8V2UfkNWBUfXZqh4LAbueEN8D//
IdmDoRtRruMNid8lXctACEsVyMfOXHlZ7wb/xx0JPvoTJt7CytNaPl9G1+vjSQzEL8fgkmrLHhkV
S4BQFiDcRr2uqGe6pimBv6EVxoP7IffWBAciKtzSp58/c9JJ/z6rYS8O8Kqs2R597tB0jCxGiwIf
nH3X4TeOeo7IhupaKlssi2AnsK8h+YirzpVRyZosEKEP4EjIfwCw+AGqB9hyDjATHpNY9neQL4ZG
CQBv2a5yZaoSZOyIKYuXqoFBQzl+Xxn6UrO9RvR7wf0IdiymTexqvSX9M63Uujbql1G281bZTH7N
rYNneAGL+KcyppmBA0y4w1dJEjyEdy/tgfhfN0CEkLL9lVLBfRiyDRFrT4z2s+UTC4dDUdQVpijV
q4648tNfH2g0VdQjQg1oOPj7q+7R3AsKM3h+RFYCI1fSP81mtAbdRFoTOd9vvBAI+dMiYx3rLWza
H3h1scZvES2Trt8jLRB++4B5/HVQ4U9Piu5+c53br5enCAH4Pg1Uy508+O1Juz3psJH1e7ndFoAB
rrqTP3eduSuwDYIti5xZF+/l/KS8HSwbKojh2bjyW0wE/9o7ry3nAjmFgbkZ3lwKVX8A0T5UFd3P
EqcGgo+hPEeyuBa8mND1eO40r/p5j6bPiUNWmPQpTveHwX62ThDmd0e7bCRxN7X//39h6WawKEzr
s0ShN/Q/+aqh7Z8AqZo0kDx0CXKynJpyO4ooGkcgmVWub512M8U9gGf4+9853/NkHHNB4q6JzUwY
L4arO3wJC+60pLsMUdVZSfQrJ8mqQHu9EICxpJTY0/h+D3Ji98JMJDKYJFzqYWse4peyKWJMowwq
OncU6DhN7brstEq57v8X0LGjV0kLA/hIKVd1SOJS6Y/oQ5iuEFdSbQXj/Vd13IUjfjVfmzZk+13+
1u4H0wpJndFAmuDOcwEyeUXXaFXlEg9N9P0G+yLnM8+//kN1QuLUBP7wa8G2KYs5Y13fLcJvueQo
gfF/QceHK5drfI3Xbnw2zaHwC5qLLBRDcJVU/yXhdUI5m71hpSF68SY+/muGA2mgfCCV4tNxiEit
Yy3w2trgsIpXzo4kgfyN6KBtotX7cfd7HufHM2qoBPsZbi5F1n4mRRrHavzbmgXpcGaJd3GKMbqU
37RXoQHx5GoH3MzwwROlOREgAKmI8+2E9e9xVZTq0PdC9dVuAeoghZ2hXtvs3qQreiiQTRjfWICQ
TzrLAflzG4widDgipKSmoSOEt+MFPAxNZigO4+satKL9t5dOYTn8xWcp8hyH7nUEBVtrbrgW3lzn
iOrteMOb/a2dsmocVX5f9c5Qq+qNyGP8nZOduhzqGKlTXJI13IaWXGENtJAj0xk6yCAAO7nOF4Bg
q4f3seHhx3rda6uhFMUtjSztbP4bUdToY1yClzITySOsRJM4K+mhiPypOf6alN2/6WO1M+T4Jlxh
uC8J3GKGx9nZDAn2reDqLntrCyPqfP+iAeDKk4W7adHAHoXsTZwy8KHniQDYsI3eTU0WyNhiAu5P
vdP+9hndZowD5VOgmmaBWmEVH1HIl2sWio/PUfKW/102m81/VjiBel/m3D7KUcXqRRV0MCzqJN5S
6TEsfKfWoCD1onLFvdVbsqzgUGOgEgD++fNK+GSHuXK7TCyS+TlwKaZ7RSinA7h7NBeJiB6EwcOV
8FO5dtu5AASUY/jJ33cqa90cjfjf3hFSKf27mEUWi+6wG7TY0gxVlaJTHaMNad/ep5KYzMUEhSg8
fTFN5eY1P7Lkm96bbGpEPLpUrkoiQ+TT0HIFBMPLrbL3nlkzJcpKK7niKoBK8H46JjgEohnzr13B
O0wjzBIYhXQr4AT/g3bexIMJqnb9VKFfL5f94ZhTO1/sOUbCDPxESylnBabd8l/gy4gCqxiyKJ5A
8rMdE02KO/uU/pmLB4aUp6vwjrGU5tyW564+w9utIL5IyxdwJIrj+kPIqoFBQBsXwoYvzvz9d06n
OkRAfyRMwO1jCM8Qc84icuXlZmEnc2V441cld+B8pZxAWU8hrjVPZzK1vyvMdpC1RcTpvv19ESfX
iYIgHtdsOz4TXvQOXtezpPmcCFY+Fug4Bf3yzj/yFoh+W+Ij1njF+lNbcVMiPUdq2YM1TH1i353i
rTjdoyPn6pbpNSboosRw92C9V1FdK+qaRulRtgB+mKVuuqStbrpwWMq2lbGi2o5oM7HLmANNo0WG
fKJ4m9X1Ow5hrUsQSmPrzA3FHtWsvZ+YT98z73xhY8OElzhLwXC0cnhIiii6m7Bl2gakx8mXa4fi
WjIrsTsNbkQsDXqF3LRCVB+czOGbqcbfgZWyLyv/LB/XvsFnQHweGttHIvAbZbUPPQ1zJ3oTn+JI
lXS1erUxw69VaYB9aOmcZghTSkCe8ye+9XI676Ys23fgB3Eat1MVzJR/u/60GWgLCbcNLrDCi6jI
BUKfNP2L1EL5Yc3LDgTXQwHuvQHqVOGFOIWUdD4dEU2bez9a6zXMfwsn1731RyXt1+fFUJzj8sZw
sKAbzA+NCEwGK4zmIkFiZS7zY5nqE2R6EL7B0PvR9z+2M/75GhE1Tfhk9q0qP8C5kcqxR61MCK03
8t4cVNOKhOJBXx+o8UG0I/WX5eOtX2kG3P8a1yV2ErcUwXRG2/zvFTd1z0NO8jQG+8W4R8xZPyo7
oAhfr6tE/ERS/Mm6LKKjmVgdOX5x+07NjDRlEWDpXsVrSPFYLQ9G58NQhxTKa9qYApB52QVH3VSL
goXGg2znTv0DPAdzRp5KxpPVasweKnE6imiODnrmN0gAI3OPJuk3VKrzUPytzH677BIacYx62uaA
NnU7vOKPmBVLiyNScFQpYm4F5O7b/Q55rbhFGZI5fAzGNQnoMO8QxvH0/akImtuRZp1rBMd11oYG
3R9SjlvbC6O/gM0szUvc9XYL5WO33YRT59QO5QAmXVybQhsfjyfctQoEacM81zeKb5scOYlYbBGG
6EZUxzkLRKfZeB8MwQ1aHayx8SDzd+Zly8JtHhiLMvmx9n/kk97mZkidqPWlgFyPGrkFAE69140/
OCcSG1YaiqXyyOdGUX7zvYceOlJDysxbwy8SEE3Lz/x5ZwgbEVy0l4kgvkgFkQ++eoQPGoRw1NsX
Ec55mAm00lHaIPA5noL7mUMSqzYnmjhdYv8jbOl+L9GxnJxXpV2H5Mi5LA9EZW1FchXKyCcOJuPP
ZTZ9sO3VoTu2by8LJtvcSO6yffUlASfL5Gwzy4HtVWWpFMRHXurtlQMhBMn2LTiRtT3ZgIpI2XNW
ZVx06mPiXcvgQdEtBE9yKtkcrkL7tEeFo5lsh2jDm2UDMamCK6FSd4cxNYYhVH/iJEvWjwIWAJbD
x02Y1LR7tZVLgiIwjLVA0gbV4WuYe0BcVqtmrZikQfbmsSiJeKSCvRt+U6IZpgiLYk0QKk1j9DKI
D7aNPz4cqRrXduEs+/dFZ53hFfpcSi1J4RCJqcAwOIpfBW37D/8DOp7Jb7kqcHiG5S9pjgv2n0aD
5rCDDWt5as0wQ8qZSMyBQMinuziNu55gHLoa3bw5oYTvSsWT1YdqS5bQvZINrWnzpgxoebv1bZ4+
R46SdUmAEexztOwBvmBGklYz0yQfmV8F/U9DVcnV2DqCQ6wku8HerlYf+uw7PCiUgILDrxcRWspY
ftqQdCOWoyReS4uD+2noXXLpyXqPx0cpyVWSR0E+T/HmTXwEVOJd04zxeotCOgZp31nFY091ZGTa
Iax2yZpUrxPwliiajLaZBJ7XAyrkY3zqeJnfb3bDYpXWLo3p/VRJkNGd49dzb/4Jg8Z2xIbn6dus
CUU0hSmYgd+ehxnmaIo74JLB/ipXqboRQVzbgERu+XfzU6t4Hb2pJReb9Y7VUQX5YBICtwGtF9S9
u0tEApVxRp9n9vUboQrcWnud155lgJg9PHQkxXc0rm0X+F6x2e6gdnI4/pyXQZIH5dS8GslqeB6J
UglkTf02A0WZbVvjTD+3YVmoOGDL4ybqGnVLKXx+oEDg3LsqRb9cskXdEphN6wCRffk8xs13Btlc
9vPxqmK8eJOkUffUa1bRgdJtk9valpiqooI7I0jr3i5akb07QdT5UhdsaBxK06sjSq+CBo0yKTWs
QU2J26P4N/d4jIRjwVC+2zO8rRTBUwB1BPmK8+QB333Y9fE7PmpG3NATAXWNUYK+YXjIzh3uoR4B
xTuuPiyIlqi2+zDVxvv6YrOQsnXro9vasrTtPCu/NlQGROH8/TfZn611CiERmc+uOsurP2+6rJme
3gBw1LsgDxHivldi1z6EeWm+cw91vXl+4PtGZqnYLshc+sMjFhNGe8rT++tVN82KBCHAo9mc6b8Y
NMs5WvkUkElFkMxZFdcyLrzYR4XaW9Ew4XW+dYDMJ3up9jugd6+0irpyF+FiWCy4Rg4io7oIlxPg
ouqMoz1f+PalEqQZGGBX6eDAudHa7QkeDSGsY+XRgRYjJVzxKpVoBNVqBPsOuU0vizNy5dkXGHkL
SDgTyI3bAbElJC2kdUt/E1dkFG25mmQAT7I07kQebAcm+cpxf6F0XYiLC5LN3NBCu9cUqyAAe2kT
ccYcjpsWebxxuCzH805EbHz1MW3diJQV2cFQeztdI/AUBZX/bN7RAcgszF2SKNNe6Jfg1i/vxz8O
Vn1BcRuxY54YE3E1E/PWZBwjr4oD6V4o7N1DttdzgyqvGT8ZZndBPdEMc6eO1g/lO2Lno8kHTLjK
oDdXMssMsKpVaDwu04px0oVc40Cf6HYnYCzvcUx/Q28An0IhPHAXPAlJDoFR+s5crgBRM6Ka2rlj
1B5O+dK0i3NmaRLtqDAXNVgPm7ilei1ANSwcVaEr5p1gWyWB/GFPNvpH8FVcV0HgTmDilNByuAP3
vGHqwxgeLIa3lhAyO4p7P4aDSlgMuLnuy+pbKM+Q+UXSvkcGyd5TC4MfcsbyXUAG1qqtob23q0kA
2vbaGnHhZJVqMr2qova/zFbcc7KmI6RhtR/EWUoVizAaI5YVwzlzCJsvDxqv7znKxM0q2nt/ethX
oLJlYVgQgeFU7I35dY4G2GItUW3e/rlWaxf98yOmpu+UbHdVvMdlhTTGbh2fj1gWcXBEcQCJw1IF
f8PivVU++nhWX7S8pOCD3Vqio2wwq40hSJh8y0Ht4FyFudEPQ9qVQx152wAIbKvanMaynVyCA/CE
CTXl8yPkrMJInrjSoVxG4JAa+viEGSrDrpghNUIlAXhKVGSmHgyDD/2nIVZn+/+WJXWTSmiGDjEF
sDOV6aaXcDSHKniAIXYp2bSXwD/b31yKaqmNTCI0P1uD8BJyGuelD6qkxj8fzm/s4r3P0FXudjeY
Jcdk+Wg1CcgpEt65eQIfLO2+ld4+M6BndxI2ft0t+1giVJ9+9EguasILFoV+7Wn2u78UYDlSY51W
2tvzAB2IZP1XAa9hBwK/7E3kgip3MuuKRcABuMsP1qkz6nPMDmqP/m1gStcnbU6B1VNuopx+eEJ4
1sb6NZDxOXpYewlF6eBUFL3v/NwZjmdfXbRsSSRD+siwqmHcXCaUV18QJyZt+MYgKB/Q/4wslIYO
Syk2m2AUv4n1Pqa/gZSfb5/9OkYNct4L66PMYa+zI4fAlvteZwLDqANXj8B9Po/dh3nSkZQ3lhmR
zm5/0Q82Pq6Vx/JJ1z8/D9EhjN5LvMzb6EniM+15qkCagO0qjMwJBCNG+D9e6ODJ7qF2U07Kz2xJ
KgwnYthAJHrqmFe1gtsWkZdD9qc5lg9Hw4EYIE2RkvTqit1PwLLL1WNC2kKE4OCbaY3XbD1HPzXz
e0RCz7WCLe5tgYj8XUUhTLaP/YxrBeQTTv0CrRtBok1PZhgjrvhutF+Kfwoc6WnRDyv7m3+P8nnw
dF7ZQIS6M/kUwlTJyujH8xibTzC7nmJrmkCeo4LNR6dqhJtQb6HQl7Cs3eZf2YRy7VKiLHH9bdJD
LbW6IObg7i8LAz0gdxHCXLAyqlQFbPFMGTKqFVReeWoNywUb9tevIf2OW6+skclIND8u9gO2cCuq
DkAueDpsZNflBKpWntGANTAA6bz0QZFIK/EPEw26d3p15pdTgIdg/VMYLux6hxDH1PXvJJehlmA4
xD26DVxFEAz1X4NwiXingPKMwSlKchAMX0mLz3fcvjnMnYRHf25qoSW5i2+EnSt/lt75lVeg5WUD
9jn+k7CCtwBhBxAA5BpiikjFONbOW3fpTtR0W6EEkZAmtbmVzkLHIrvcqSYBCZhTueQJMJvAruYi
YshMsukQoHfACfSfiGzRcMgY6Voz10DNCL53hT2IwpNN6Wda0q9lajxz7k6buX7yK62ErUv0LuBB
c0BbYtQtkLClpaRHkeqgTefCm5OsRTL/IqGDlSO/zxSxCuBxk0QAUy0Umt9385TBbxLnVI0IGFRi
1QXzS2IMrDSSarJemqn5s+NeAsEOExPpCEobPx+uUhGNZd8HitU9thcocuOWH23EqQRESHRBiktU
mIvCTmXHr9HGtKKmKiTnAQmUBbPV/LGTzmxI74ORbXgctz90gnsTf/cntp0mLjGo8xfyds574eDa
vvHyL95dBwYPwwXoLxkXke8NRp2DaBdiagPjtJjSer3uQeFtn5SFXPIE3axsVINvkxr2vX4tzV4V
TBIiQolDWW2/x4yzDz5oB+WEtQMy+kf8EF1tEAwrn9c6wm1KZtvxS2uMzcpzflBOr+3eFqPIhjCf
y0c/BdN4pzKA8jblPogepOkVn7lSv16CcV5u8CSYqRoOQRalBUMIr2UYqpGPUZ4qhF18SqD4d46a
ACusj6cgaCrescVmvgcfJHIVDYEoVO3viKBO4rmLq1SPBNbG5pRAORTqjAd6470hbFc7AViPX6Yw
HCII8K8P/TxQk6mxTzfzGfb+zvi7Gm2CV8yeUJGr7ieXfkLkLSc9L6Bs9utSVWMHSzzVOIyd4fZu
RMr5oto6H63nA+/0RjEnOZljrUZrutDqe2mIC4q/YN1hNqJq+3WyICWh7fQbP1PG1LpBi8TvEOPw
nvA5Y8gULXIlPMwuepA0ENu1V2XdftiSiFe0svMN7mjkUSo8Ukb8V59mdfz2vzh6rZgCOWlYdPBx
AO1SbfqTNJ9qChpIzdRvlBI2VS6CAH/tD8xyuWkImVfNlNsMKKapXcHoZdjZw4ZHuQqXYSJAJcps
uv+/etZppFoaIhZVTFu1hriduryoiIAsS7kghYWZfKp8TkQ/At1SRFlOPVj8c3gF0lAgkP7+08CG
NYc9w8A3xBuqsEgsGtiTzUlxYnu+Zy0oGbKBUir6bsg94USIeU3r7M2eGK3QHFegpOIZJOuXxOit
XVi3LGeG4/EEmm0OegW/wJg4XVk4HItbDx3097XHLTE5VUNIgRiPj1CyBcJNzmJH4usStKOQ4V5O
q+EKPEYdS35XKT2u+R4hpWvm2a3Cx3NLxSHpVS0tWnz6SBWck8sd5WNlYTv19gs/tSEh1n7uWrXI
Ndf7Jc3P7ISNlKaE5Yr4n+Q1l6xW4FN05mf0JQlL+fGcp1GmI1nxPaL6E2YESBHX93Bd2aPkE8PH
EzaIDjAGFLoKYHAW8lDJIR9qDD+MfM74mJHyZWLOG6CfuxJGxtZryyzDfjnokUyYTVHO0ymbw3Wm
eDY20rUsvoro3vZAzo9L4f+HmkIt6PErZYa40+XjrUTppavFW4+iFcMz1zxD7hexf4jnSSnX9Syy
Wm72wTfmurRFzAD/kstcEtREgZ9UMTtROz39UQzn2Zbmdkhkz6p4RW/orVO1kZAeHA3S1eKz4sOu
E27/l/49MCM6W8BqQLHJtx7kuEmjMyVIbyOHsL7xrvtbhHB3MeECbbFJWzUGa45ZqEfapnmLNa49
E1S0CnAPwQ/H/cE11buVgZSzAaZjlIh8OymsZl2xoJ64fIqyZmiv0J3QchDOBR20Okp8dojeVpic
NMGAk6JAyqUCaFpe50KoeJxJkuQB5fpKKxKQWFZbOdK+MzcDCEqZXf2xntqbcRcFIouA35nHh/UM
to+/SEvrLRYhdevQrI2dxuJR0KEPSJvCaZSE0V02FPv/ZvYA0bbBX8r/kf1birjKqSD+z7rd98wP
YNN6jeZ0a2psxlG1dX+VY/2/y+RDEGZQEDRNb32VjvDOyKrRbc93tXrxKk3Ms5El+UjE8YPQwUMI
yq8b755pbk96XrYPUGqH5MTFkrMl3hWiYcFXOzJOHPTdMtsmM0rhCtkToh43BeBRV4fVAWWfvtNe
uwLZuz4i+udyyG2eTyA3YzUaxGEZsCDmOmM7smdwf7muReztBM2G7cTz9irvpalRzgneu7wGB/o9
VSNRI3/DbB/PtwHPipjKK8RA90JwaHPqUwET6xAVfCmV5urf7YuhjG6eTdEn72RA+O02VfNX5hSQ
1kSprDC+rLdVT2GAq8Nt597JBlRDljkA8jaeoLIzZeDy4tcG92itJpmxXBk0LqpdTwatoi+SKyu+
KnMWM8qVqct6ctdpApyzjjD2arqb+9vZ05rUHbV7FmkzdAV17eFstojPTZUMpihCVdZWF376YXK4
KuIMREirRyaDThayRfrT3KTIwfyau0dXgd8VQSzTEHPRQXlqf35evfpe6+kowqcSXt6zIVv91pHc
ws8Xa6TWdA2Fmo/BZ+DJqbcBTwxuPtqHG44/i2Qnm5KWHDaLTfjiV/nRgDbNazSeHIhAWfKRHCeN
vXFB/Eaat7i8n14UBWNZMaOeCWRprvaO+AtqU8QWo7LuZh6HmL3k/0y4iRLScSNntSCQOrm9J6er
eQNn20YjDunspdmG8Cr9C7l+JS1yw4BNb0PvN6plXjw31V8elQfV4uGjQCMkJ8BDTb4zZwKP6/Xa
F1ikkEuyo+bopzZ8Vy3imCi/Ynfe08Go1T1yKzM/NO0PVyZyhibP/U5iEQ/DOlEPAblZF1mlFPrj
h4tNbq6nN2GagqGeOK6yw4q8aRJYWHMHf1OLkh82CbWpZN8vXkeDCyYIfbwkXn2LuAZM1BsUDVhU
KMQ0WKgBes+YE2sFSccmTIOJM5ULL+JZBcSsTQKdHddWqkui1t7d49HX/gXydY9/eubnCKFTSknL
ARb9XcCtt+hX9NZJtYimmafxtV+NxwUvoRWzmtXHoU9tylFq6pMoODYHSSYJPVXyzofJtwSd+nbK
yFs+8PZEqWZz0EaAK/k0eiwfNEhEJWCYhm+VEEDmTA+FfLKYVPabKd4hZZmIobgsYN0geUtr6PRx
IoGiO/74nj1OWc3JxKazZPKIRVhZN91Wvcju8a71dqXv5v0dg2Ryzj8u6yIqAJdFXdWOTfmNTq4e
vqVINFmjk6itmR05bnmO68xnLeY4nMI2/ZN57YWG0TLnSjmfgnFLvYYxHzyrELxFS34u5o+dznBw
dhmwaGbJKSUQqClmgv4L9zsVc/CAHwaolHP/kp6GtcIk5GXpJyhB33eT1ua+PZ2/c6P8Wg5AwNLR
owZTJuki+RKWIY5tgOuAFWmEbLBsB+c/6Zs09mMzW9qQayZZFXtA+hipNXb1JMMeABhrHTB3h+js
3uci3o447qYwXZO+dx2Cw7RjcMTJ8nmIZhaxybUQ6efvZXRUmrLel6omi0kqLIm+werdZDzMChdJ
EQ7eCMbl5iW2+pGbeXR42xjLLm0ySBI0pROcjqTG1Bnk4LzPw56Ki/f/r/Ir/Fcm5SDNFLg98trf
hBoDSNVwbVIe4LU2f18frK1ruyrMV8zeUYJUtNH5G2FoL5ESYA4tAKaiTQQdZkmDPVJ5dyOzRHHj
qfxnZXcmADvXNwduDtfQ6hN1A4qK+O7kS34mT3oRgA78l8Rg7vsYR98XeL7wYLG8wkuaXdImMBos
kDKz+re87BL47F5j65zunQoZVX1wQfPuk6YDCzsq50fnQcfjV8B3jxrrBmTjuMbAaWxiAJRrNpfv
9yLTuMbY/86ldePL1rXZsQMXgKio+z0x5UAPC9/JaMYJP/TI80HweZnAdiW9Na2PxMKVz1zNj4LF
x098ar5QNGFDa7naRiup1c9lWQ7UpIhEamXHFlZYkjKMqZlEbmcdUxV3i3Xp3cP4+3L5+Y7mUZI+
/RRWNetosDXfh7WrkopJ3HX04SwT4qEaxYO8bsr1WGTCore6VHL4XDxvmXKf7TTol19XrN198yeI
8pzmo22GVNvGwC+WLZf1X+afP+wkVvgNQZraHRsfzcwN+zIeBrKDFS3z0+vshSieTD9NZkxh8AEf
rvb2axiLwGIu4hk0am9J9m0ZC6uSHLPTAAMfKhhjQDTL0QjBxQVb6Ufh8e+jbljr0XLQO/X0k541
60Bwm8+6gx1ScFIgmFHjiRwfxKgxSX3HsHuKGEKCNDR4EWhbZPTojU02t2xG8+7uPlCT3WgrfDNt
1xUpZrQCsoHeuEEW5vMizrkvSXcSxvoPAZyB1lDSt3oqPPIH/jK6bbvf9+reefdigMJOCkFzO7+M
hh4NakN4/fZMIrMDBkAKKryB9IGG4aZMXoPOQbDpEi3OgYJuPb/Q7K5FlUjdtSvKj/dN3XbZWK/g
PLc7dx0p2bGoIie9bpncq/Vip50nLB2tieZztvJSKqhTlyHfuxcl/ezEiZX9qgAzhxJKzx9dlQvO
ri1ydDMlOexUKa/5VD7U/gKxh+DTGZryJvBGqGgNoYEh0Rpv0bsmf18TG15FYiolDF++B8/bU1jF
puv+sd8y8j4ZRHYqD4e+2TKfLokG48hZqkFdUgwjMXU7agOvdNamyUV6MhuAVVRJGJ7goHSh/rBc
wbtGWTtwUvS0UGq0VTZf2B9MewJcnX1ONorHZ6sizrECbTPBDoqItiXeF/LNd+jJ4r3WmYwYWXxo
YJTxsRpMigesHAqizyYFe7E8emHwyEeFjNQyDJWJ5UKyzzQ5EYU5C1/+volcsmqqNZGr1Lr8yh5L
/hmvX+HM5fzD4ouZ35bcgK0G9jVpeFlr+MKGHhhN38yAWCj5iHDIrZ9pjsIyq3kr4MfIrsmantXD
zjhoXtrCuwOZWZczknJr9AXJE8PPZfzTKIGkG4Bwlx3C5PbLsNIzOKC5FoIygFNd5BwEVdNO4+jg
jnrZ2eRwoex/9vuuPwWKzhUMC0XlO8EylSJaDjyubaDJsBBrSeLcSGJ4cYD8MuHfb10dRiQotb/q
TruEU9ocgBhfubb+qSrx6tLAVIgdHitK7q8udc5rrkaGS7f0am4QW/MJQmWwv/5zrPBmY5VrILTH
7dAoEpYbU7OSnsD01p/kaYFYqeoQmc37a2BdVQxjG0Ea6KmsKKGK9hgoWwYpKS2pgdzxqOobOvLi
Zerfk2Dsx80F1cMq/IX4wL3f1plJq0GHBiZADaS5DtgUxnv4ue8MrBaTTaY5D86ng1ERxojKLzzt
aLMJah8bXwkkmLxUy+Ayw2Wy73z7kzvzGcNtxqxDeSDSy4ub0M9cUItV9uid2Whc8cdED63kMUjS
5OYviLAPtxTvPqLREIRrhWEDLMqtz79m1dQeVHbeE3d0EjC5l9AAGLKr/VCx/4qRjzLcSveNgRDv
jniyHSt3GX4v25cvhZLt95CHx+v3Z5cBz91/da7OYKNkw9XYVThsDrDPDpw6hNOS0i2UK5IVcEiR
nrdqdfbOWF+QGSbJv/MzzvhUghrrtW2YDPGDa2iNGFuFSqljs8U74kGp4MOI4hFRZIaQMdO5+44t
sKBd6IAsxExF6ArOUa1IrsomCZc2V773sqF/HxwOq1gb/Re//kiOODlSDvpMztscCfF9b62flc+c
t9x0OAEs3vJWPH+jkaai1PKLe0jLeR/IYFmafnKEjyN9BtGeRfL0Zhe8J6W04Mw9FjLmCeY+bhda
bDYZ1YGRwEfkKw656Lb31jr3En3FR0FODNIWurhHx91Bzwou7tz/kN4kIrd+FjFG2mxSCT4jp0sz
bltR78VjznqdqC6INidUVdm9Tg2XF6N3qWWYe+I8zxfAB80+defru1ZpgGenPMqxxGuFdt3wldVy
FbYrnUlsCqWTBYBtvHNV4jFjeW+kKyRRJEYuEFiYKCurtdv4WG1JTxJaUs96w0xQTecUsaoltPw9
wgQwo9o31UTE+9KUWh7frmay99KwnIiaqQB/S/f0occkQ7kbke809kThSEaVanUoqo+uGxiZbhJx
+xwbCupq/468GgFbdCTRn1N/ME66VwQRX3jlVogen89z5iiLpIDYf1M0UO/sUSpJ/5I/9yjSjJJ5
P/Wm0GsRnBWlMBN1CTWcHo5xnrqSXaBiIRVh/CDrjDsQMXVH7REiQ1K8j3APj1gQ2Qp13/qq1lr0
NJx+g4ciqYKYqK6ctfkkL0SfU3urQ9eE0eFeReuTGtdJC95F+5EFMPdFLvdGtMCjkaWchpfrc0FW
NU2kC7V2mJ9J387z7OMU0ZhjjTqJsEHTgg73PsJa9s5OF3Q3Pqif04wn99sXj5ZdPRf0x7XVy2G+
w/zrfIMW54TGQlsse0WIBX18LUMNqqQs/ve2UUqEMvXXUdD8rdwWiTIe2boorp+vJhn60c1yKMEP
SwE+2eMAaWAx3xIDiUqnHElVH8RftdVr279XpgS3dVFafOKf+FvxbXnUU9mryMnmeGEyjTko/BKC
l9QkE4klcLrAoywaSHm+IYF8u1KllqkRSatvBTPrfAdcmtqvTfrsLzDyCrlxFAeg4mVm+dfV9aMv
D3sTwDBrCIX1bBkHkA1f0H7e/2DSrTEwzdNEJEP+ZhCrJaWOTTPNbf851wj9QALNWAg1y2sgdQdH
QINzFY3QVe9oB4ytww+wEWQDwCD5BoyZMrb31lQNGjP9KbTYUSNwPCk9yY0GIjRoiKwIXDY20aAm
Yb9lL5N6PGkJvk2gZOGFOrBHiwhcrZoNlab3NmQ6FrUA/v+6sS3uYnXRdil+z/P4Pi67bismVSu2
8xexTQB+ORUcSe0cs+tczrmENJq7Ka0RnXqfcpD6An35fYBx8pRODrt+ujFqc4lef4TIEk/2h2IL
wjYDvDf5ea9MPoybJPdAdQm5HvIRai3IXIkFxjGZhf5yRNaKwl2z9PFh2vepdKvwb09cxzJqxC4w
aRHK5922/xQOkZ9cMo3b/sBqa4kb4hVzR09WJqmEMxLLZR8imSD5dDc1VPdwtyqYpKlf9cWan8ze
FIiQ6vTZ9x2Y0n8qMiVDqebr/U+UhsxqekGA/z+rcNTUqpG8TBlIHc9Gud40YNgvUf70aqZmrDNw
H495IVwTs28tWj4lzOm5VOnj5usiLwCi/VdGEYxfRkAiKUDiL8Ng1ZCiryrMWxtGs00EMY8QBUuF
yPXmQYmw4oa7uJrv5G6SzywJHbl1u38M5hxCw7Bp+2qHwKfnOj2Xu4PI0GJiEXPfvpwQqsoyrnCh
3O6a4SUu1JZ0mRd2yGI3kuVo32nYUu3TKxrq7Q0xxbgkJBKyM000wazT1AAKaoi9UKWcdGl+9Zx8
nImXFWJ+AxPPKxnzOA4Tyu7ONIQmdww3Gkua4tJIAPF8jHtpfzPkc1J71rdyNOa/dROn0QwGVimJ
vhRJUZLx29wr/Z8PAfDMPegddKhU0drScR3y+dSijrAsnjZkmFfwdYQNkGyOHc1hZHM0BZ/8VKlu
UbTU/9B9D1kz5M/ILgN1Bre49oaRwTzBnODsOGLbrbbZ8t9ds13wHVTJ73+2lV/RauGROlATH+jo
wqIdIZVe90W2Uj9TFSw/JWXLgQcAz/DulpnJEs9WKSQjCUBIi3EJJ1C2w/j0IWUcuoodu+p4NtU8
7Qt0dirUySyjOVHQuQ6wSkUDxUYLMOGabYBSpt0kLpNg0OGfPzDNojjHA0M/hpvZ90MO7kecja+6
JSao014Aq3YRmi6Sagn7knAYhRzjlEQhpOF2xeZ3TtafHRGnMzVpJ7KWFFTVyBaf0OrAkF0Ht4Hc
PKWd1abbAZc0BwKJs1YEEvTLMKSAJBuASjC4dBvhehu9dk1mQvmqb2kS3FdYc6f2vEUaIZg+bKA9
SVzQ7/x7QlappIg+apnN6WwjOiuBCRRQrMGGWUnos4QvWxg7QvYixCPO0UMIy9Ws8/GeBh37VCVu
zn+kyyo7p2Qw+wk37M36tp7vs2NyumU0c/9ksdH65qPtKOEdXAn/nYEaAS9KeFAryAkEcshTiJ+a
vf0Gu/VXt4qw5I6+IVBg/Bz331726Kws5U6I+vt6ZGPa7QrH2ZX6lBM6q5h5Z5IaVBz08D26QDlw
Mzq9bnjJA5n449APBnB3T2Jo3kc4+gKUITiA4YFYxmmJz7WKB1K2Xow6wzZS5/uVbScRbF0mbsuR
NPhl0tAL6Q4ZINozcGsQgxsl9QXFs33poIuHYVe/yuBkdmk58PTJgWtNc0/C1qUubkuVMySJYI6T
w/WEm6OkdKQf4P5PCKST2NWufyeXfnmb66F5kKgUkbO399Svl0VbwK/7WsVzXldw+N2Bxs46Cmar
22VvTTcWE7kBDEWJ95puyXcadgwyik4aTMClXaHSBbthIT6a5oxdIp0CaPvjh9wIc2hwwOaliSG9
UMeqXtxLwrCx5kAwKY927KEqiPXIlhf2srJODPtkG94vcnoi+R+6hWA90GE5jKdyU/5LUcpZaXkI
iIBusLX3bLKFwilOderb+Wbta7xsnZuD/aQ+hKoIegDp7owimladsNw8rvfmbiLVowLVSuXZiOcI
7wqw61B4HvhBWNhXYHdCAyqudDmQS/tt4J0TKDyUuwQnXFIB6D+efJie6IymyD0Syjq80BZGWnmg
BYg4LFpVMCxTJ61LYMBQ0bpw5dXCn7nGTdbrHPptCGkuJ01kp1LjL4SMFe0SdC6s7K4X5f58sGtZ
DdFJ+qkpRyoRgmAEU0YevYBfOmPdXBIgCp9h19/ywH9ZOPCWPbqyfPkQfx/6mOkkNGoR3Pc5bg3a
44POy0HN4jz6CZEY67HeHjBU+eunNfv7Mif6oxMTu0ck7UceCMUJBDexe6C7F7+EhCCB52QY8mIe
dB42RQTnD9V7sWUYJnmU4l/+rTL3dKy2QsEWLDqLZIJlBUntfzeRDQymLEfM1aKo7IwKOrIL7LKN
uCPt3gpTq0EYHzyO/z+lPh/9quMyAF5yHRWo+mCz2IC8TqAs24ttpthikgw7gTfLmlBn+bwGAaPb
aOtGD8dxdFJ7RsuQqvb01qd1UoBI1voMgC0Yxrgkg5+RROYRlKdw1zX1+DKi2YW/VQGgCUlazHCt
GtbPmdGyX1RM6WnME0a03idVIxDNlY6lW+OjtDJFQGJ4KOYP5yoewET5xg2uiyzialkV0EQTQ+Bl
hoQaoSFjMUusMkuJHHn+fzTvEE7cv+SpBYe2e9tFq8cjFf+3w7tvCl2UC44rXNSEv1B7/SMTXsGQ
/HCoFklexJ0DRn0P/bxmk0ZmbR/xwBdjfaC2yGXWcZEO++YjGCNvPNjKXoz5DsVYwP6arURefGyl
Yo2zai9GQAMf8bMmkoMW9+gSQzxu00sRQlh+sK9TCTk31P/KwcxZIlbURxRYZd42jSbo2EBAMc//
lRiW/juV9VHsBrj6znI27M9RSqns3nfWjKmu0lBP2wrRQIcrN7qSw/hAJ4GydfMpaFP6U35+iUfa
ThO/6Nyrx3vktKpzy65essiPUOY4A6aB2SkaW6wWfbAH5xw68XnvRjfCp16yGSA9/5vIyD7SJGZR
jxMvS0MDsBZTKB3cVtatPM/TbS56VXZraHEEuGNxnDwLq+XO5V11FFrvkkG9cFs67Rm0t6kJmqnA
qzSfUIGyQcMLgJGZsR7aMKgGMhDzsNO1NcHI/lkn1+I+RBu+DUDcJuZ6v33tYp9a8RxlxJT/D7kn
WCDPF71Cq25VnNQKL8ARcr3056E/MVuUVOK9jI2e5lrRuzEpPmng8x9iU/z00lf1ZB0vu1hkib7R
B4bidtqqt0t3sJ/zIkPypuh9B44FvXLqzLc99lEPkiSQGmxiI/2goNrptcItog2f71/7LrFOfYT6
YHkHC5osWdu8BqESb+sCnfha1y8EbTu47Ul454kvW5eGe9QLzOv0y11PIfoDApiOx2QAE0uKIn0n
Y7L/D4bg+uJ19Ue6VlqsX6MhD6lJrgBvxAIMgTNvuIMpXl0tmlAGxmDhpiuBAD3/TzE9LDy7EIUF
1Wt2e1/K/JAwcZBfL4+mcOEsmbzeAlohnM44v0EaUgCAr8qAc5KRJ5V6NL7GWFU++iJTRNnpVWJ6
Sx6pFgsDokPaNy8NXCbwVwhK74/Z+Z363th/Z6dBdYweZnMP5bWJymwK/3SEk78kNW3JWodzzHLV
knQch4/sBy6OIVMD+GAO7ua20XaEBFw8kU9ZWVpMXgrcxu8I0IpGk/9qN3VCf5hFsMI0XjpuDnbw
CeNWbMMQbJwg9nJFneruL/hlnbgFyb8Sq0pfRRMXxB4ZtGK8E4ok85/J0tcQVcoUdWk071DCInlY
q0MHkzLzNaalbaipiUlB+7cTs5GRQxNRYKX4xvUHWe47XZmUMqEUP23xZtc1EegJg3vT8aMyMDb3
06WxfX2+JY7vpRLAWdoPTmKB6vkvPZnBO0LImRyk2p42YXtMOq8/W+6zNndpPqNCoj+/H6+KN0jW
2v0e+vcoUZqWEYbBTiPZWCe00Q+UTkVEu0kbNJjjtHm3FhwKQ54WPpixilMW1bgaNTc8Kq0+1gJi
GRWHokNEwio6uxkv0cUFDufYvhLZl3ibvl425IHRIxrTjk1Bj6vkP2LWFkr/gDhtdSs8Zw8pJrp6
v89l3RsoIwRwyWKIoCCCy1w+ayg5cWjJkI86Svj2X5KagFN5DyKv+rWN15rXJ4mFTvhn3uutskkK
CLPfNNAzKV+ArxpGhmGyNbaiiZTdAa/pwmL0Syf629bgkDPKpJEZW8Qmt638fMbPYGMVlkJvpD4E
LuNJJAVfPRphzkr/3owYGrOpkW4oO828TpaEyJeGbmTy4quQ2fSTp7yoAd3YCZPqHA53PP84SnOp
a2e3OwnK6oOlRnFtnjBnskT3fnivFaZId5zy0rI9JYKSJAta5nH40kDCkuEJCuK+4m2rL/Rwj1G0
zS76ORvMvSOVdC+ufbIxGpJ+dE83cL0396Y05a90F2SORlNzkSzgKbyEytVaBFx3X5ARLd5DU92M
wNO1N8QewuVq61v5TUB9rGXsBIMZ8kO9+xpyVT2+a/E6vPK4tdzZBTv6AYrU6jzL/UMJy0gcvPhD
OUE/LTCkG3uNBsdv4PkbpGBCpzZNyDriVUrImQVXCXNNBNix+ZoBFxfXfLZCj9JKNN7JFkzenYxs
fbhoUFjHzUGkzVnT82P0EKrSJYO8HJUb7F0SVjKFw9NscXydhsxpz0WXi/6NWmgpsHuTuivIcNsd
zkxnXq1WOWvZaj0lNPjNfUtVv0F+NzK9pzV5cy1cUtuHDnT5UGuMFqK4QfHnCId9sQ1BS5Tp1chG
UiSDszaqufpRyTKUnRFsxxp0Wa2gmpVgS8sIYUnHw6rWDpo+VzrUe558Oft8eDWzPRJwjIhg4sMt
us3w+Xx9XfdB0ZYl1Gdd7/NGP5MgiNHnZeZE3Bu0QAOFaeR6eMhkSgFRZgMCAm3ZH5wK9tyl8tA2
6W0Gs38xLBH4sjCokGG1OXV298n1fQEFFzZ2n3e71grX1djvaB2WV+7+vzcBJQtEH8cK+9BxLpwU
BCNMZ5sK68BMLA8c2W1Px3UAHR8CUhUlKac1qTyd+lQsZlse+HgML1HwhRLWW1WNHtV3yHLhaVwM
JLz1G4gONtLhdcCNiD5rfA+JXCaIgyFb1o+ilcQUcd7yBOx4VeByJPjpOPxamc5DmC/3SIsbyXVY
WTNWWiy25tPbYfboikgf+vHlO9XXM8YyV2pdDFuLm3F4I+ma4wEWrPZbLz4QgyZOeBynw2RVYBfX
KBvyTWIK6+o2gpv9bz5kGTOZugF+JNx9u4BpE3uXchhhotfojoqT3HMXwDK09GIbOAs1hdBAwYoO
YdRG5tVQvjq/d2glVs8bhgSVaOBEp4VBGS1uJSZUhu3rEc68S+cefodE9rH7LGhOmojH9VCIr9g7
zGFV/GTWDOoEKRJ+hEQE1gtXMvIxisasV/FtkrnmFM7SYdG4MmgUoJ7ShRTeOK9MqEuAd2RF+Xfa
bFJxhBTufBK4FGWJX83NOjjRMYI0xyNvJ/14ScwT/DLH5qaNTgfsHPeVCElsiy7LbYPEAJYgJ+9p
MQHEnG7GUJ3nuxNGFNKQbcgev5GD2YVchDXQhKT46OxNzJ+FRt6mfidll4P3d2S6KYyZz2yWM9Pa
ziFhIRMTRhAQ8N+2y004JURrQ0/F1h0RIq430C8cybRVrH5CrX09KZ5PfzKjLHCH+SjDPI4Lr6qu
LeGL6HGC7og2AFkBYlfx3ZaDu163WR0LfCpZk6qYB8gpwM0uanx96ygSxGlzOdSbm3NwNXsCo/fH
AwD67F9Sz7OUr0zF95P++QXSPGJj7jy+awxWQXKV2WpqjvlS7/SSBI9toF0ZjwGq48u+wn2pmhAD
fGKUcPw54u2AxWrADQd8CWWbGbSzQCoudN8DcRg2qdmrA0MKQvNgEZqGR5gDHyY9g27Yr9YXQwZv
jgNU2JKd7HFyq+IwnueDmw7VmvYy8ecUjXv8nANRRbEtSJnCos+IEEoFjhlP6pgMjgFXEn4bH0qA
pYfFhTwyfVpE6i3fshs2uukjOUD3uBScSPgAN2aWj9lq01A0oDOucsRUZSYyccYr5H4c68Qo/caJ
JiKk+497HOte+ZEPs7gEEv/0b0o6is/dNryvpNHRmbIoZlbEyRzOdliOMDgNiAQlLAZ61yMfVxKs
Z0xRLO5GRm2bJU/NUkTX0VmNwxYRWYpdjoljsbwOld/04k7gsWNR09JTd0fYZ564IefPNOpjZyrm
YW3eVLt0IuLd+89Dv6ZHIZitvPQdr2zMpaiDtC/sNMriXmALPmr7pr5kESURaq7sarGocb5R1eFv
8B3DV3UsXIS/AJ6SzL4Wk5BlEKdgmYSQ7Q2mKSuaExkAl1HaH8yuk56iMiTgif8C9TquWCp3iI3J
diGcBlm158+e/hCm+esYsT6OCzT8/QNEgwuOKTwZ8gdDMS/r/reE6Dva0WvHojio8wnzw+5IyQ45
mxGWyqS84dCnzLEOypEfbYcYcJJnm+MlrAzvE9hH96PIbSSmAY5uGVlZ1klf2PorUEECpTmv8NCU
FL6CU18x2MV4ELnqDa5+ZC383cP7+51ZPQDLvNSm+v3hCGK+fSvli2CASDODTGKUUqPGDmyZLJeq
YOZs+/Tsxc8WbY6lBhDUeRu0UvBSC9IL+krfaCKqIsPriMEc9hdeNPMeCjUFx6LQTxS3GMWWHxV0
dULJ9tJHZr1JpQ2VwR5din/fmLYSgdzx9gUa60RkoC9pSYjCeqMbQ82u+ry9y3nK3DHQuuGibWnw
AAmreyF9RMqOdTdcCzSxTbadTmGkiAW1zFX7b24oYk98ojHFguMlh0AKPZrmMZK7+suN/cSbEdD/
QlCkYzNqKRNJidjxccFuBYn+DMQlLwYuatIL5jJkBChGpeMKmwaaWIXmcf8ila2IxOhUCiUozAEl
WeIKnmEB+7BpUz5P5hOLPRpO6a0SbUdgs1Re8EeHWwmzKUYHTW6pwZnQvtoVz9kRgnOnoIXuj9dl
QVKh8yNyoLItTlxCQ8pX+0bWCNQZHJEieFArKOWHNqXme/E39hAQ9NsVgDREcrgff92oDeMkXuco
gkoRwkEz93cIlZKp5VefZmGv5/YC6FypNIJvHN5B1zgnVRVQI1iFX9M4l6gSGiO6z+F74P44tt0N
6exqtSIEGxNXWsz0odc8aC+xOokPomyAl2edqhOEJlE3+9ogIdOz+A2wzsWQSJ/ORZCVYtGfSV88
CV+P2Y8Bm4Jb5V9OyyHCnO3BXT39efNK64+GDFNw6m54oTJtCzwuS1vwNHRsN5KrH6vZ7j1Cme5M
UzjvNujLGvBPJejeowcCSJHd7FcrMIX/nYOY7Gia5wgpNsFee33avZuJpRCN8meDGwt3hugzxBQR
kD2IFmpZszqyB+bxPkHnnX2AKB/WearAcuhkjZafdBMVrIkwlO9aSLpD/XJc1HF1+jTl0eUjnK9K
Hsy6hg1Mzba1+heEe31Bhvwii2oXmSGgFuZCxPALrF6xKJEJysfwIfzZ957ZkbGLUXnLj+Za4fFh
RM/pE4mX1MAV1Ym7WuMdUAoav0SL9w9uHjEPEI9wPM4p77AsZtpTTAeECUcn/no/AytAXkGkKFad
T3u5IG6pFoxziojxQ0DL6QGIKPfq0EEaVHDxSkOPPp4zzDRQneEJX9L65oob8JBVymX+nBLZwejb
4oMr3tLjMYWINW2hvb+G/GjaIOqYjRhv7MjQXtK6ebsa1//scCyVv+WLuLDOhQtCQ1nI7L9inQ8y
+cKtoHhzFiPSEXi88I4bDOlpPekv2f5/jsbz5XOaZgr4uV+sTU6RUAj0iIopBcDYFjZNSWSVYo/s
12rA8com0WkYyWVRITFavMT9Es5gnMZlOgpijpl8MmD2yd5N+SPcx2Q5surLEMEPrt4jPPLctogA
8M7Q9yc2i91GQiYPXq39MpQD1O7b+fSGVKakNWsa8RwP7AZ/7xiMaGnXrn+yVAS3WhkdISA+4Np8
sCQDOpCbfqARlRfobqIlQG9FLYjYSogdUrfafh89vMZnAIPOEujnob9XWu/qwtnzWx2Y5TxB3tQ/
eQj74qmrxglEbBVwc1ZsMBOniEEJwli6fo21AOSIDCbkPB3D25xB74XUlcr8vuyEDYLDLkP1LmHj
LWz/zntStko2d2zbSWBwt/GVV/03nmb//ZVVbo/rS7vKj8FB5uJFrvfb0SAf0dkrztFonfKuVGWd
eQ0mM346TzPQ28J77nqALoFjCLBZ+QZs8H+uLvtJkaws1bBjsN1G3nKhxHb16EQ5i/EnEdy3zowV
TZBPaXgUb8OD5xcBObU7rqYLnp5aahpHDr3uwsj9aJjpFOlpLf/ITST+YJ3TRV7oxO60dM4eX9Uz
zA4Hy0X+mWn+xIU6M9oj+REthAoLTE6yhIHPvCUbnPoXD5HRQ2RSCALu/dfDFwySFoObaNRp+X3H
uyD6PrhKrEuX9VlfY4uWq9lm6JzXpEKG+pmiFstb6dsjRjuvgAlbCBtiZhTCiDlVP+pYKLRO5voe
CMF8bVKgEZnYKCNaXcgnHnG0cpy7c74FoPnnei4+wp7UxAfO/kFdq6Lm+TmQtRST3yULKc1rzY3U
FLaEdZBWidQ8J4GU3JOe3CTTEwTyCcjZTI0XefCEz5agi1HY4mWeD3xVDXg1/WDSTe2gcWPpHEf1
PTMWLbiUhqY3Kfn1kpZGzQDkHHnARZ16yeFSbKK/vIKGdmE6QhM5TKlAieR1/fXHJUR3MX97OYIM
aiwNk7lhunVJRofXqBuQf2f4TSrqI4JmJfpcv/R2LpBR7/wRmq6E98BURzWoIK12e79MxAb64en6
iX/7bQ5tRIcFdkzQSo7F5PIPeMNtpvnyz8V+FuvVh2vcVR0JM6soMu1FuYDbYw9tSPjvvArCZdTs
ZZ8uFmLXDYnhjj4f14pQfMjFADUejq/55tJ9y2BwnEwgtyT3x+L4ZLtX5sPBSVoWptuMy3Lv1+zX
nqJ2H7emAEmKWm4rDa7VP7YUenA2ebwsptJz15mtMjdjovgeoNwjee0h/7BynW9NIP41UVUJs2FB
MiM3U8qPLVuoc0rlUVGS0g7D1Tn84zOHA5CTKIPSSfleG4x6YqLZGShSrFQ3xGh/1zqMsUlRJ+uj
fDnf4bADYKsCuIpgKPUM7kCG9v6HO3uQpq9CUsrutsuI5sBEjY4mkmyboxEnICcAfx3En4EzxY0Z
zqiEslVoYINIk4jhhJL7SqvTKlMJo2UCMfAlo/MKyRftez+f3WmVE+jPGUuIynwRU30uAZeCXqN3
DFReTqFEDWF9AYZmB4AVo9v9gUardizQuyhtR45Iu90ss2wNxF9FoUUpkM/H1LJJCTyIE+QU6lp3
FyZHeSneiN6zAkJthg4kFrEq6bbQAn0Edche417yf7ODNoeE/BsA9scLeodXiAhV8AWFrOyAwKms
A1imAr7CX5yvEi6g3QOilJ3cQuzbqCiRmALh3w1D/9MJwNh1lZvXOyLgGIrNT1mQffumIE8EM3dM
dVsfTPfiyKgEPCKKT3S9eOZh9tmvALJPYkkn0PLDpuihDl0S+zKn1hm+AkOB7O969mzrX0/znP4Q
yymLXaLPNoAMnMjbFywlDvmJM3HnbVCrrtmmOMRbC3Xm5wiFYN3LNloSdSmyj+j3r5MK9EXHylyf
Jbtmvxv/6P0N2chOqdaKaqAhhCJ9b20QXIuAy4MdnHfIx0YaiHWx5xceBK3AYGDOrQwQCVVPLkf7
5Tn7ZO/8SxvS+pX6X9mRd2b255iTYRVeLjymCcNHwVNUbewH13hHgoTQA13J3GutEZ1KR7/0JSEo
7P3q6j5Y/6+QUyNkwvaYdJe8CyI/xuZ09AbOcWqVtJmTQy2zT11BV5WIdy5QFfpWRlCw2frNBsee
qAWi2lwLfTeHP1BGtAPZlzlnCA43JEQ8MDjrNwyOSKneHAemOBwOCyh1OEwKYBzVE8UnqYjm06CE
tiff0cmtUPPO/IRs+sKlZQhhGyz15sT+9ncic3uQI20wRwlxPjNKNiVFz4AyylGX0FP1tp/T9Oon
oUQp6v/YJ7DBo0Z2ZYRgD+87HEKMgYCIaeISse+z6bZCLUuB/amrc65Az0wAXToMApUNKhmLB/Hu
QJzASpyeMjGfB3Zl3aAqVSGSglXQdY4HokgdBYHvGNeRaEOxG0HHRIRKwf/g7wuKC2DZJF+IcclE
VIb0vK3OgkRXod1r788RohagOL6GR+z/sd4Flrs/9ei4mIYfTu0hkbz7qESIhZVsd3d6qhRiPTqt
Nh1MPPNFWn5OvkXON3VAoKVbQwDyfxmipD0rpxIXTU+2n8HCn2xueQhPcmFkeSTyerAy55hEvAD0
fuVDATkVzBNT5x2mjH3L0Zcvt86BnkEGKiCHdtvffwHhqxY681K96sNTmzAEv70ajCvaR7dX5B9r
F0M9S1AyCO1yAtaMgDDXosqSoMFuTIi/2VX4cKmIPy9H3w4T3+z2e+IDGZNV+nYMXyesKPrZ5kb+
FzX5/zx5Iiiq436hRlq9Xb41NdsrnarL7QVGxhDpK3/ApEr9Zo36UOdzFt7tGBApaatkmqBvyAks
9xuIlynOe+RTOuaS4mcWr8xvsezEiWkvPbP3Idr2f2Q7PbZ/IPEdjLsimNRvQCReFfM8cgmujwTx
JbscTZuh8BAVF83yBmRjCQ+b2Qu+vage2HmbsVwYXmgh+FnwKmlNtnQneqKheWmxzg1uleguokIp
Z68Z3iPH6shTGgnr1H7ln3wfWMIJELqR5gHAN0aqbpEdGbDajXGlfk/JqJfhCamPvvyZsTSP0hnp
eCpPQXXYgP5CxpBZMAxjtdhO5IGwR1jnimLt9FdbJufVMJfSOZexATdUbot0LjCSsvdPibUwIRet
qeuRPueCVYJuKzq0ACia6P+bA75rurMYBYp98zwmaPnPLeNONVPx7g51oL2X0TJZjQanouXc0QJd
FuRSioG45DAgiXUtzFY1Nkfs5aUzto4C+ZXWooL2UEpocnyx58xlTXP1bWEE3aK5Lst7fMM+Jkew
5wCvXBSZo5+1DhYqxXeY76M8/SC4wq+xy4i0MNucSLuqilNcf8kqUWECWJiwXCswklZnXtbNTuKF
j/ceYHIDbdAPKPYf5vS8Gl5n/Oo3580T7Q2kL1GmzL5blZf9pxGXQLOFi7/6y9tA1eMnwEZyOvOc
mNndjZXMLdIrezs3kYgr8AXBlvFWeQU9jKczI7EQviT/QcQt/8Zqlna+s5dEFywhVyJtvJJxoVfm
GhIt634NQzrxtNsBaAH2eXztnsUaymxjwxAPKTYqt04zDH3Wl3N+t/2awmUqS+CVdI5L/MzO8q1N
YtbUogtYEqvIkRP5mi9Ei2nya1+D24b+sm4vgZjj9njjraoEmJygE2Gi8I5Xi4BY0nX/uKANzmpc
sy2Aa9IkSl8RXdlnoQOQYLwc7RjwUM2FqraNYMDm77/Xa1w5Avr5ShIWfLyPmEtH8BEvyNs24AY5
KO16MYR5vaZ3gSohouNchpKKcPQBsmtP8UmWVn+0hR/ARJ72mD8dqulZGEBwKVZQ0Qzjo5kBtHUP
T8K2iPJmLv+oDM1HD6LJFShHf9BOreS+lIb5kQYD5Y4rTIE0K7paLpq+48dCloKrYo5s36T0L9NM
CiFaFQZ7Zxx/FaYRCOH9QewIxmYxoWevymHw+USRD+P3e+2iTQWI3ICxZv3l29y51XuqfRSQttQF
/X+THyAdsHOC+m/ABrqpN2gckD2jnvMaOnXbLQYB+pYJDnRkjU2EHdA4JwgVOtQfH01k1dBOozxY
7gbWQp8Ul+kvbMYqKNCp1R9ahPUXXFPxP625SiH27fj4wyDSgfjSkRpxKW97IKDw+XOXaGdVRCq6
iHw16UFyxSddAJ2hFTgbP79426GkSD9Kk+uO0Nlm5mhriEP2VSeZMs134eUTm6t5Dy3XqPmo+7ke
KUEILteqQ8qF8awSx+Fx2Z/qfpoAyD3MJuSmhyQVgN8M6VeBPCjrf1yFSBbfHvNxVABs2LoUZ5SQ
WbnkdqNHQ3yDoDVjNiTuY7DqpuKCXyI9Va2LIrpM2778VL+MBbFeEvleX+cGY9ozr5VbSiJYghpZ
rJv1iCcZuJnAEWcgNuATIUkbOrvqOZ+ZBdrjlEse9Y7lkcIuBOaDx2dFEjaYqhB1w+7dGeMGeHfi
rzcAyE+sZJ+5yl0J67Op7gMjFH096GqA4uhHKMNVxZMbkkXuMIw+WaMrRIxs8JO1BuCPk0nZGMo8
LZ2krKTjNDMIpy5EKQVdgoDXZuQ9j5Om2g3kPmoUMTRSoM7sVsTO5S+O53V4dwfj8KR/fn1ZMj5U
47feBOBJOZX2yPp4h8r1A477ldAqmynO/rYuQyTH9/eyq6stu01voy9a2NDaEd6zyVUFzW/RzDKH
K8+dtYhuzJGXhSW8YidTjSVIFjeb5D1B/8OU6jMrC11iywGA3E0hkNop8BhZjmAJ00e0JkI0Rt8U
ZD5wRgjo5+aDjkx5wtiCxUYOtuiu4KjFpUZqf5Eyvh+9v2q0EZwoeFYV2+lwswOGa2eM1XSwvkzx
gC0rPxlHz50HJ5F2L1q7isou5s11W6uomOARNoXA4tk+c5tEwOBCVWVjansDbLyltopOAW0CLfEN
oVZGB+13ETJF5+13eX52YPs4RZWLP/w7nhw8p0YuwWUV2VHqNNHdeKmw+Y+w9Lf0SZgAq63qH5cK
uBJHeuNSHsdy9xyLWI3SYw/ba1+JhWkMFSLr5EELFD/TPAazg50cORMiwe468HvAT2HNolQX6iwx
xKsKHRMLoKSjTcQILOUtRzWPErjIqpq8llCHudVkSorjkllw4+kupMqSdSORx8z4WiHFK0wGbT4O
jQtzETRHbBAehUtBI17C5XnZKmd6kEbhkoC0x1zc61ygx+N+a2ifdUJmF2yH8LhEa6BzQfTeZ7go
9TXtkqygHNWNe0WvSP7H7IL93rNxY+QRaNkn/+W6SkxPWUpmuaV4TPsXSa0kYtIBDLotPC9zdEVK
GYR5ZaqTpYQK5Vcu6MhQPJ2ln7/2f96gedLjW0JI3tRe6Ja4UkHoDNXxg8rj4j1a10zChg1L4BZr
IATQEbGr/sQkOnWyVuE8Y1BNpFoleg3W0E+LO61CQAa/0RquP8O58kz4KSeQ3XOGLen3cD1sbexR
4CEpufuCxKCujTCEPe8Y+uYxRU9OgwM5AwpnAr8WKL1a1npm3/3Dpgvt8Dgsl3ydM7/+8eAc89Td
KyLnQcgWa8q5jQfdF+GtnfIRRrY0hfz4UWkEfaePhiW+E3uYhuzEaezhNaAL7QjInZjDKMGuesZc
chu33MTcg5PHQSi22V4YQRl36AES4SshxmMJzBesce2h50j/cs6lMYhsIhQ481vEMTC7CAOIRXAl
swDvy5BWgvT06LZBC479sdyWJjZVW4c6r55nbLeuXri+zBFznaQtGL+aaUCyKyaEIksxz2tLp7Gr
4XhMhrpqX4o3ZK/qkVH14Ee9BF12TeSViwLSUVETV+iFwgioQ3tXwiqmgvBNlBy4COlaIMGjuDEX
iL1S4qdVGQDfcPw5Om6LR0I2WL3j07KdVKWfwK5ZuXeOayH9q3a5C9L+fjBuWODcqZ2PONJwqROP
p86JmziDBr926W9bNWCFgEPLpzu55+QnSvotV/3/R5Yi5MN+mQHqgO2KXspIpX0TVDSbkozt3FXC
ZJA1/beZ1acuiuV0c33A/TNBKo9DcZR591IgbR3tUYQl4w2AC0gcSLQ+mhYNu7O9YqAK4Zg13ZTA
AEmHNLLt5cn/7yIC02gzX7zoxx5sWAWBcfFIT7foucUGTBwMi/TvHTQ7XwAqYqX5aJPbjn33fKhe
ChZKnaGvkNE7IN9ygJH8anYIwM6i7R14//eenpfiWMOnmTVNUFtj6uQlfVBV35YzXARHORm+nDhZ
eDpDg/ptQywJA7rqpDQadmMOgL7QL7Slt3PEIPFUE+moqBzs1UPazvvCJ6SRHuXoHkdKB7EsXj5K
+l2jQbPshSi6nEku48rh3APW3GsdZKA2RppLxsSplmFmrxfqvIvHXqzOTEUvZ3Y1smq7IXn8Umxx
1073NB3JDXYOWMcTVnGQzayMOwRPArTenrIJrwtxRaOKUDfS2+RxrMB6YwNG7LREg/fKrARYvvoa
3SBk3hUvs31qGG7bg06IddABIgC5cvAVBb3HzQ/F/xe9R3e1MVGWwXTu5O89qBF5eQ90pRLaAB23
hHLmBd6J9monVmR+0IEIMfzLFkJwDr7cskg6bt85rs3uoU32HpOesjh6eH8nv3DAkDJEC+RE/grK
7NEWM/cTacqL9SP9XIF9+7chg5SYTJRiVvbvX66OgRJ5rbWZ4q3zUs6aOWUAe8K9ZVJ1PBzpCAT6
wSfxTtDRUsbgmpEjzErVYMRXRO4KWIOfvyWvg056thgfgXHKX8UJiepRgmEcPzgpZPxqd73MKNXo
6nud0V9SGbL6sBfwc+cQMcxO26CRMsUMYri0uYOGEaoptAMH/1iOkF0wYeooLLYezb/9IY09Ty6c
sqhqDTHVtZSKDhz5+6D6YwRmW3Uh1XUmupCZtvkIzvOz/fETQ8vSwV/6nk/ZCTWl8kKC0dKYYZ8a
hP0VXDTZDUZ+xL+D50xZPCRJpuAFm9hvo9aTHXpeLAfyt8HwMnPEFY/OXHEPdqEBVGX8tTd/ClXN
5RoRUYB2my9ElswBHjf+5grrouRXyIHpYdvxeUhdsKhxO4M8gz3oKZohbvWwUIJi7N7rXXh9WWKq
yXzFAXyuMOMRbieoGjjvuBI1xs2uATmSdULSlNvyFC6rlpl4r3n/PDI0nTVEV77G+6lg0rBliVJb
W5UTqEk+jdoPzMlXcyMd/imWPaUirDTf/wB1fRMdgCalSR2wu66R2u7F71izrNRmMuBnj/4XKd+j
MFCHRiGAv4iD4BT052jfYufl5eVT/Q8vEc/2SubCUwk+k1hz+5Z4QWVD92OaUE8/DbV6OkWjltpK
uRkGxEV/lxVMrQrzxAWuFtUsWDlXDZByB8rf/mbM00rA/NPdh30hcsRAVKse51ZqXv1vflMqo14Q
SLnM24bmJXHmMDsrjhuuQWz2K2XTHQw4T8MpwUAat1FuYJBFw+BTRVXM6cEvRPtLBO32vTRDx2fM
pV0WZiNwO0lzs/XMAzTXZjPIFH68p7NJ/BNJggcbMw4lo2XYHJVRen2WIftn2r6gtk0FSfxmIi47
V2Tq4v0qQKmKnzxFaJnLFWC6tWIL5cJaZ9C8zguNUUsIOMMQUIrm8CWy4eSPtyszcjNkXg/dr+yI
Kcpw8de+MUlC+2t/NeGaY84wlZN1Zq/Y3Nd2kq0vDF0eWVPG6fqKqtEgokfaztAofdqFxSZAdceC
4sPuh0SRgHxOvyx4nIDiVA+m8JV/u2WoLqBkdlrXcOscugB9H5lg8M85obg9sbxTNnggqfigEEF7
ygx6ZqN7KvW4Y8bPINw1XFeY9WSKoP7fg/iGYJoOXL3Pd2n0eJpemA3hn5GH+qzfpsg/o5M6LyNM
S5MU8Cp1djtto001BQSyYntfw9ElS0Y8FaSV3DrPyvGeTUZdH/cBuHel/2oAhiI5bejV8VYVgLsp
Y197JgaV8EjDB4S3lFWtYoY/4Fj1eYB90UJiXNymamj5uqDkjWaV1f4KnJGIMGKrgPKxYOEwjInG
LpSH4lA6QSRTFqiSa8IU1LcuvSAnvb52GVqB3jbCGm4esKwJov8Z5j9Bq0Vza6TJInkXQi6M0DBu
Zwe6SeskwkWwDd176ErKs45/xamaMXBVwzABY0cD0c1CTR9Bp6af5mVN8wMyT7Ekohvk4J25w6Rd
agbEHhxLV0kV5nWSROHcuwjKR+BY6SyLDbGFd/kNzg4DHV3z3LOUP5mVKaoSeJD9S0QfLRC98yFz
01xaiyGuIYxqEcfNcPdQraHOR6Or6eGoiNf629j4PvCOwsE98EJHiElqnOrxl9TUanwWc20MYBFB
Sew492WfMDQnHcGbCzzb6364Bn0uWDK0fayZ4FhLvqeReNzjc3xeli6WwG/F8kf9Jo/cZrXkwjgv
6ZvxvaIMuUw9JYAQNDWTYSiB+TyZVQO7NlEenjWW3J6NNUy8woc3qnh1wDTtIY0B+RwpmMMD5ILb
rlfKhc7d6PY7NDnX7jHj2TZqzSZ1+srCX4yux6VGNjTq9WqruuAhkH/07ryK9tgHclAmxQd5q1M6
3p6lFRP7SFRViI8eXiUF3l8AuJ6l26Pt9C6z4lE55na5jAZ4EE1Y1DfGekHX6o2znOKCCVDS0MkM
ifGQBD1ZmbcsI1QUxhrnCJADElMDDZ+7ie32LPnm+4iWhxEElq7JwsXueQFC2nae8ynWOsW+2ZSK
DlSEPeKfUpWcDihV9kgm4aAMHHQ1u6nVxvvTexP1mJ1ZbzcVNyoeRaYcug/XxivBt34nXlWwgLd/
RJeMwAm9GT0E5qXY0SMT2zQJf4ZGJ7S/gqlCINJDjgVFZvzppIQFcbaqpRQ0j6o0AKj0dJyurJGm
TnvI78tQ4Wsi5E/Y2UktrQmaB26ntSFMa5t+bU/cKK05XDN2noLWE7bJm3U9+Q7EnSr0XcJcryZj
kNgW92uOAtnwlwRBJ6mAW755RnlEj+a/hLt6WL5TLQemsBeH9QvO2wVwLUrHTKbdEplRP8v7AZ2X
jFbloD9DLTTxjIv3K6m/Xg3ZxDNh6gfKZ7sFakBRkn/QDiO3OZ4PSa+aVgjIEJ47mMKmPc5Df3v8
jK46jzUn+J/vm7P9vqppej25AMCo44pLhMK/bhjufsb91vjJrbE3j5Bql3LRk0tQwNNYBksSaxOh
3sqJLdYddwKqp5hCgx1y+hwVS2VojieIkq4cCyWmj069a93X0gUIUog5Dp5aucpVAm+BcS+PvxcG
J6WLBg7Lq80R1Dd9z6M7zRSXVu00oid3nBPrXadnQvs3q0i1lY4eFm5MG3c4RbvCQ4W17GjVPCFt
3eiQ/ECk1oNAdLzO5s71dPSt8ckeYtmb+EqHdlrbagZQ0w2c3MsWJVoRoK1Les5b8fkcjjTp67wz
2R+9nisf+Be/m3w+/rTNtnf5E67yBdGCUCwwL/RuAC4NuVWLY/In88s1pODcZboyMdLacN/vZVK0
LAZnvhXIXEDPt8eQedPuZ6HuyOmZ7aKfOX0rZSoDxC0hVMUYxw4inkGCIvCus02ldRVJ8obVZrrI
0a34ecqlFEa1HntfWy1jWl0eBPUG+wbHPg+xLDS3uYvcw0Fn7+99Xy1Lp+qkdkXiDutI092azkST
ovwhVsKJa4+SifN2MeQZ1C9wVYtO4cJ0eaHnAihlbSpRpvbvEp8DzkcV2ClhXd2D9qDxkHtSgG6/
42dz/uw/YJIcXryExKGB9NgORsY+VKg1LBZQJdfvgEHaFvgoMx7skcMbd7eX3rw+ryyK7CfDUbNf
w8HOA2cJdlschigUWgOS7rUK3h3u9DNkfY/8iZKTKtHC+nd33yR0YdhB3mi8CMJLohm+01vBsSlW
6CGc45yTMHYZ4VSLToKbcVFd5GyrlnWpsq46/f+XIe8+8BvgcuL2SgWSV8tZ9yj0Hsh2LdMnzGgo
VOfZQGPIm+Op8lO1Al+87qT/sjLPPeIjmlaRJJz4FnmSCXJ7eAOweF/mjND1GLNij4hqhqrDHbmg
vXQ2iNu7S4erz8GYJVQ0dMMYOOL6nK4izROAEIHGfAJWqx0HifUSOt77LhBbIa/o7j+cu0xWoK7G
5+SAsQpXQWnPe+tU0ff00g2dTvXaRh9NKMmnl8Sq7FjNEBWItQ7K2BUEUF35MqDAvqn/v820ZlFj
ICKtwkeSrGjkzX9JrWA9x3BAApuPH19fq46DZOSoOlsyEwh+/0T7rSzV5OfYfFJeGNBMtkBeTF6X
oZAC+TptO6H3w9s31rOvXc3adHDtkIA7z6Qo2fkzqCVln0yNTkklw9BgOA2PHAph5DX/h9vJIpH8
tcg0/DGLlvpnnJSIDaa90O1rkujuPdr/sa3f3WGKEkgOUEF7gBgRD2ThwBXZMHGyQfqvc8cGS2Kf
ICa7JANicon9+0+bM2Fm+F0LPVI5CMaZQMPx9FSx5xK5bL24fDOqrAC+sKe9i2h7IV7B2PNlQO+d
SqI/2DmWzky3taaAcvicQGpw4jIE7UBu4ydbuzDBTN3R/IgikGTlK9toyfD9LBGWmtuiMA9KeqUj
MsO85+Lix0rDsmW8NQD7pKWBJQ1pAl2ekrPd97QI6cHgp7kCFg2ijRv0oFuIyexx9hRZWMd4jny6
Bc4hOc+lER7tAAjmowA7+MKhqfBUiaP9uCs6voFSxAje0ZKvkhY/VMCAjDXriGp5fswTOu8U9ybH
az6ilzu+c1zT957il2cbDsQrpmqCtIH9viVAwIwwvc3tyd7tBcM5dhKBlElh5UuzIRJOt/XF3una
zv1FaNAZ7kWB+E7zxN7isj2QEQY8aKx3hAxyfrTtCE1L/djCA6bz1gar5fQmr62xrPdAey5TTmiB
j2YACGcAJmEoZWhZeBlEAh52nGiCF3uKhKxDuMvKDR2rnlLIHnUTIuvUgveoz3Pu+yCKFy/BVKS2
2R5MEtrqvb2tkMidRe7LeLsju57qVeZ6hR8dZzLqB3z1PySFAxS2aRxQyOd0O5osI+7QjogknYK/
0uaU3PatPFr1DzRto2sXAGJWmtXiQiYREz2WIgC8zB6STJCQGCQGZNU7HgLFAi3Zh5/UgfrTfhV/
Nv1dqVSdwU6i5lV2bSac8lLC5vjL0xA4YVl7RQNzfnAIab0F77l/4ofPpAec23WdWtEjyQev62Kx
sJS+Ah29l4eNEuA5leTAMWz3zQ+LqUHkqfP4KBuiPrJGeds4IJKD3qItD6qfV9xYLPjg1Dn6tV93
x5eJSJO74TpasbYda4SOOOYlviQ9k1YeDnh6FM9bn7h07TH3GfspyiDL+MZOIe7yY+XA/uLkpf20
fjk+BFzaIzpLcmnobrXCDFlqQtZd5ZMaF6UkbgjV5OqocP7JrdzDQLbOxRyHXZH8xrz1/MV3NOYw
pMAgxauKO8hrJMytGwtSo/OIjsF5dclT4Dx0YTGuM5xIme77nORo9GVjYcldJK/w4z+h8pK5FvFf
dKT4SRCJw8DWhjSLwwv1ILmNHy6e7bY3MYIPr4p35OKq8Y1EK2w6ui+CNd/H+5FWoYOpYOZY+ss1
PA6cyXQlOQxe4N54jWu3qSvAl574hOQprAis4xL993lOJHxo/B+ZI5nKZgDDh9e2SVlRyX+wYdlL
sJBq73pW3MT4s+mkzCJLHP7QyQuEVwCUcgzw4qIX9K9yvQW09mEar/FOAvp9dcmHmKROH6OeMKEs
lWlsJ05pYjE/EWVvolc9ZM8L4DqnWKgVN3M6OKV6/4P+ynUnw7FNZQJz5GRT1vykgOR5prfoDYiG
22XbjVHfi+naA+6JkchKfibiQVWUjv5xA9YB3T522TjoqMo+lU1WOlZ7Lqv5wYhdUZKIryfFeko9
b2Rm8s1JrbCDXv8l1kv+VBtvO6WmMTplhjMSgpnrcebd9PIAIiQVUydl+PYhYkx3Fp7w3R0IFLtj
CT4FGMgTAUsDON2XpbxPoBxTgMox/DiTBA/SloNQQk4/gGmMSm34lrhL2UNhihEegceACzXvkOEw
CVJ88S0E2DTTA0043l0fR6vrJoy6Lp8Lr7IMVbnPidfKsvE4JzOXtkSFtC14koNI0ryyzKZVlPP7
YEqywh7xcOZfiQYOVCXjFAO/ynO+459wIf1QsPu30UeAdVOURe6737HbIGZK3t/dXo9o93Lw8MMY
RhyAUJ0ql8wrO+f934gEpuawLpYL2g32QYLPy4cgzHLgx7TCp6Iet4YaSsx5DEbBsqIZw0FLNpRq
TzNSu5yMeLFYSAeAcuolh8fHxwMMIpPiTr4tSIRFnp/GjUTZbl6HVnGxsEfmrSbahvyODn//QbDW
h3e2w++BMWyPJkCVIGnY4hzyOAFkm9MQN1eakediM6tBYuowcAeYjWilJzhOKgVVvBVPR9RsRenL
b4zcfT/suX5YD8nfHE3UasV/2NN1p/hZ1p1I4vUo57l9652R4bQkGbYH99Kt0LIwf04z56XPU/ZG
eqXnCZhxZ9LGt+2op+smHZiXtkY7uwRB/NssvQYLKKLZoOzRLfqEnfCeD0eOBoISD7tz+o2D/ez+
WJdyYOhh6wwOhhyOoXRUHRXEQ8EKskMIAzV0HsvQ4c3qGZPOSUwos2NEggBsTYVhTT5VijV8cUM7
ahsBp3Kse1PAu/dT/E0hRcHq2nNibU8tjpQ/hid706G9ed7X/Dt6Ar0/r2JZ+bR22HFwHRZibviR
KACUd/bAAFL8aNbbl8kcXYb1i1yx2B3w76MQrHT2MnrauR2l5jJNpOAh9SaQ4HVToGYQKZAV962i
NeAyR0J0Z5WnJfAVWH27aGHbQcbqevkCfiqBe6PS+eYvPPdrpHG/s9SLaAc6eUWRy3LvX5j5OGuv
8UikZTQYnn0DWxgaWn+Jp55jKAA2oL95f8FsVpLYNQRO940TqUAh/ExEbMsb0EbsDOJLLqlzY5BD
mrsfwginqge+jWP/p+XxzXtT66JtkIJ7YOt3FLXLo/ncT1NGfS/EofypYeuS3FcmzGuAdcJunngb
XSrbtPfER4iyfwZYHwUT88TpNfGRNwmZ7GNobwhYMKo+pAgXu9B0d5Pin5dI1OtDTqGyy4itwKFi
6vufC6Be1VDf5siwIEK5aHQcqeMUctuMTIXN8+gWHHXFNLVjC0au6XpFkk5IqUOvnFslt0qIuMqZ
5V5E/bhVyO7PbyAOzK5cvzeov5od/fw0DgUsUYwf9H78a2fAZ4++kbJnNVLFnSxFJ/9F1CedRUyj
dXnWjbmPG2e3P36UBhZnOSjMIsSEf6MPKeeEXMjm69fuG1jWoC1Wlq/oSmRIe+PxZW6u/jyMWIqg
xCW/hNsdjehLdAG7jUngdKSoPmlwFDNo/ux+rShr6m0FOpnEu2ZRvh6fOVZvbtBQ8SJf2bmwU4jO
F1Wr7HzKKns5rqaZTNb0HfQjRX44wf/49r3wt0/dUooo4Ak1pWLSW3FT5eVI/nkMCkEeCV3ROdiK
otG6Odb/yfpk0IgoDeixMUAEALH28gqUIfXFvWKZXj85o50qwIHAFXf153zz/RewiAT0Qa/RLpYe
XiG8/viEvN07nxDbYYhVxlB6WPE9kg2SAL4NcFhk+/+XwTxsG/oxBtcw8Sdv3guSW4xF96CJENYm
tW9W1fL83S87mWZ0YfDyF6X23KhDkFal6yHLDlE6ex9Ny9Rw5Ai17/4Oa6qSjm2KcYFiCmx6YZZf
9+WH6qPo9FI8Y6lNvQJrQuBTOoIoUIN0Ae4pgnkbl+AaHmyl8gSt60RPf7rO9wKrOdKNp3yUHLRn
U0HzzX5Ylp1IEtxsNjdeLexIpGKlziXPjIf4U2Ir2brjDmlssEe/HpZB3MroGsY2Gr4EorbsISNY
5JqM8P3s8Ehn/zT3Gg+XMp4diPDYtxq4IME/iZjS+lTqy4HBspyg9z6XBOj79384dJpDpZr2Jj+c
coGbRayTpwKjBfRqUReZPLcy3LXh3LgsSVBo7mhsKAo0RcGN5Juwbr62i+xbLRNW5V3q+yaNGOex
zwGWW2xamYeYKb5C7UuNAyBW79U0dk39ME4YqWpRSV9MDkeLQrdP5K67IVxzsqb2BJUWs30iWel/
1OLrRLEtAfRnS9l3PeCcJFrBLHci82GKBt1TOESWiTcbafTOBWTYJ1QPIfdE3yoU6pKX0XXGw7JK
rTLrJmP78286c5Vv/B3oGPbOyfpLNrLlia/J+gm0pRD+oi3kDnXbyQk5vH2Bp+TElyRteCymi7rr
aEbA6/ftlu/WHGRmaAIe0bAPUQ/PKABMqjMkk69+rkUEQqeCviZ3seuD2tZlNUQwq9dmK51hQLHZ
jh9oDFL9hMv2JgLlEcrWKcWXYkQnSIqV2a1TmbvUf6WuaIR7Io/Kd+d+Pcctkv+Q/E1BDKtpzAlU
4Gr3TDbGqOpSzZXWbcJ4MpQLn3gj4jMrDxSYHi2yNMRZ7oPCvW3ENERTfzsLOuOfC2bRj8zjWzcp
ZCbijAHoHB3WIMV+oQTEuFHddp2dOD4kJS/2jAuR0j/c/CwSfKyhARyVX8yIAp4cWys2j2pz9Mw6
8rGk4ADPel8KA5SU46b385agrK/0PheIOwaR0S0FABtrMZAZ4LPa9hSRW3atK+JMJoVuLEH2F/CG
LUQ2ev3yUsv8b4jwDHmOv46gkpSFpjdnWXFWCl9nsey+JVI1yFCv43pScsnmWSiBB7VBBBCUBDuD
L4BOYUGu/GryziXvf3WV10ZXKmRUOIDUukfmhDUugs0BUVr7OFRNyVY7FKulVE9JIeCpcePt510I
o8iI/Pj0hJoEQuAndYyTFNfCtERDtLAJj3sAZPK+Wtu5BCbnfVbMU3d0PnRC8v0bf7IxTDSZrnU1
D5HsNRPWWZe6dcBxS0VWMdQFlypoxpJrcuRCnidkb0nnPpauyTGopf1zX9xZIGfCpKzCaGLhE5PA
6T942BJ5UQep5TGKa9i9JxCxfXuSWGXBWJ7+fV7mYdWTf5KeWxekuaXA1samlTI6YkcO/qHKRfiL
m75SuHMnKaBr3GQfatx7F+fD5AK/Bke78mTwxky0vOQbOXGiLyz5Gay7yne+CBt/6vBWy3ETB1fW
dSQ9Su5ysOYEGL/LBLiRAqwRAfF+v1lnvaNDkeGKoPO+vh0Ae4GxyFvOPb2zO/1JTq0I9SIr2M3U
+OAFNaJxPrtCPfHTO4ixYcIcdLypZ2Bei0sCiUCJkf26pxKEm+m5F+o6HXouN798uyiSDiniKgCR
M122cNN9azNe+AkryM2+11jeWDJ/XEAZZo72JH4XINhhm1PGa3C+M/jpQrsYKRD2HAtnyNq52qaw
NCmC4rRF4Fvtr1VCGV8QdLg7CWum8JsG/0iXA/r2jAd8isyxUsyhBVjMRmEw1EprTdlouA2LYOUC
rV/8m5UifDp5zTuWK77MnOpQvByourQoEaMsfnoC/XQkhd2NzLALC2MODz0fPtCIA4PJi47ciTGp
A3clFCjnPEVJ1wo5Ec/NpFw5YefjYou7mtQJa8ZvShcbwb/Wl0jqSQiTg99Wb2d/COfc+WbUgACM
GMel4cvxTmJlyeVWq3k3f3msUO2YeLelHwYsonD6kiN0MFmeVgGa2yEIAYzh/90pigvzT392EHzc
5nyTcwNiLrTosAOB0r47f0D6M0CzeL5jkeOXRPVkyccsOQIHD/mJ7eMOcc8UoOA181GXq+2twcih
A/dzaTCdRmx6GbDlA2slZajC7bFhvGZly9rVIOmYuDrXHaQ18R/RppayVUflHKJpkRrWAnOq8wTw
8QdYfSlMs2dHS8nKXf2+pv0V9NbYA5+EgHbzako3hDPPOAO73LLkeptvyIetxozTTkuQmRlBxKhF
1P4OROjFZ3XEs9T/P9jrGLImQHgbxS7M+bD6XWMHnWdmsZ6DO1cJPA6jKZCjsBF263w8KaU9uacf
w1Jtwb745a0Fy4Hd/l2Ws9mROx3mOiNKomFg2DIMpfB3fXfH8QWrUVMcNFXl3zvZEXkWqz4zJVxz
gx3HB8sUEsssg1LY3LZDPEeGl6AwPNSOX6ay/oq1Z+WjMJIc+6AHYVlPcE7q4MkADAGlA36s+pZ5
7ZqXuGqHyWpU5xEVkr4+JoPaJns/90PU4AJOrViyY7kp7aAS0MaXWhuVK/b0S2OBJt8ta+LMRGfO
NURsk/H0Q12E2cRcq+xdqFamPfC3Bndc4PSETJvLZ37DeqsJl4vAbcTy3VZYoo9R2MKzZAPRd7xN
Zbs/+ZjWTf1Bp/gHcyhaBkHSaBBcFGMS/1RiH4baPHU2Boo+OEDPJo9SGJKAirtzqm6l3QI2o9As
XPBtpagILmkx3UNPzTUuiez0LzTnzAq/NG2b2jivjK0vfJLbIMlVAgfsUXtWLctWHiDDlTajN/aZ
QuAedRF26XZXrNc72Y7nek7XO6HgmLe6p/tM2B/Pnagua21pY8dXRWI54RyBYRyIW8kkz3Ekaap2
jmyBbYuZ9oTMf6vHCb09ngAbogMM9V9NLNuI3TiXbaM7vrqNYApDdZFYp67TYsfwOuZZ0rRiN5j7
W/8xmdnfaNmIuD70Ndv0WwRGYdMGu1Mne8DHJkPe/fLIYPglX7xMEySqfY4C/0LZdmTFanOg14n3
c/ysRGtHPYgipOh1/XdTyrtOqcOuuz5ACPut6DasqL3tY6rmyJazZ6y0EN/T6E8h7TrZoavAU2qi
hpLwolZqNxf1huYrzAdNwbz67y6UMree7UxfqGbZj0q0woEKLn7FcGTthajcAIabLVQPIzskAGbi
YIDxxRePwg8LqgeI5ABF4bn5EvKxASfLNzwsEgW5TVY7OSKbUG6qgpdwHbYyi5u3zwCPeynszAf8
CnRI2Y9x4QCBVQHjF2o9rnBy+hOrWjR9aPhPMIkwmQy+3iThKOIwKof6wPXhVMfbp+SSntj5i9pT
f2n7UYDfetpSTtKi3pi1okvC3KcasRVe2nj4bJ/CJyZapteYtMxkMNVrDOZaUO+kM2DTsDllM6ZA
kv1GBozYTHrdU1g/jSsFBKM9W/Boc4dPcaF72jd/UgBMxD3hMsogyB4Ne2xB3+xwN9+hfH2QnprP
YoHKEWNQ9vPFfIByQNtSNbOhLVjaJqK2A3ER6DhDtmzH7lDLGu5WtodKiNsaPeoYuAKtm98zwnl6
E1Kj440XCL2cphxTPngaDQRBmgbNxGcqZqRJ555cwvIFXGTJehD1y61izpXCT/Rk8tZ6dG8jb2Rx
nZhc2YrCdNpl6mWRnbT9rH8TE8mK7hVAxuqRoNN+vpzFqVyEjO/1kiMNGc8McWS15J18X1cxZEnt
NsxTegkSD9gD3pacxoBPFQZ46BJtVOIBFCGfhph7In4w7vJP6Z9eNcfYQLH0k7Om/H8xkgOcxl0x
Dz4w17wSJCJgD0O/yM9m946Lh/NaR3sZ3nxbbryUaxBX+9LTHmPLwDhQpIibAPk8V1uj71l1+vg2
SBJlBT95E336Y4/pVi45W+7eO6I2OefcvGVnEJoE2XwiJ0C+IrO/yCOUoCu1eOEdUTZg8JeZN3FQ
DfA81bbVMOZLyHFFB/4kYzxo5thrz7/4cliv+VAWQM8MbNOqhFRUrru8GF9pM1Nbkb4Q4OMfUEBB
cewIyUKiBdJD5d3rFrOe4XhC3QNkC0c6rP2oAW8Tp5rXSkw7onFYBNuBFn7W1l5aX5swY5cMK+gK
KSQn/rr+a3+HEmmj9Lwiih6NlYFzuYqNIMlWp+Hlp+BYERWNLD6BpnCuWwSUrKpdm8GE2c+yC012
atdYfGZZlyLc1ND3ivV0fiQ8BhnS6NJZJX1GLLbylGk2o3941yDkTPD34eoFjodHJ7ymNO0c6Xvl
ZFCsCzgSkRqkR3OECii06BQSIeIskun3NNGC+SF/cSiAJTEoOzwLNzmWRlM6kbO9HQ4BjE4nZwkm
RUUuCWjDP63nXXdp4zDq82aHil6aoZxyH5MyCXM488DRldcTyKDtjbua3CNBWqw78+MFd4CGmUk3
kGQH/0NcS0OwteuOhNYXEJxjO+fTfn0VblBVY606birYP6bu56SeId4dFSh1EvorzaCjw/tRnIGl
hj/KgVDrqOJIuDOidBcsr1QsmonMBbwtfoD3cEqmbTK7X/a82O08IJKapcMpNvN5sMd4C6RCcYHs
4YEHL9BvEsZ/Sw09w+BdSBAbpk8c0JppM+sSuvrKzJVM6aDaJ0T0FC69aU3j207KVeQsV1eGxGz/
T4mCEZb2qaztDULrxwuM25y7bntuKqt/tyylc3804O/I6eZGBIG34N4fQZMM0iARuJ3sitVRNCEn
72+MBWJWyN2PhhN9ZI3yM/u8rp7vXmVBupJj5UKrmyWq0PWYTP36sQ5AlBgxtLju4LjB1qBOZt6y
l8zj9Max6gHN22iKEa78OJzkm4GrgnGNvgucL58DjONGUUYXdZORmpAKK9rSCmXWPT+95xiJRbrK
5RHhwuChnu+kfyB4aaNTWlIxlK+esuhpoGvyDYQCMEtSqoPMqbSlWJgvXN5VVysdRZd0GZ7TPS5e
iUZ0ymLg9pZUIrr8QLi8aSZVM3euFngrznS5OxfZfItibJmo6QdV+VwDzWuiooLRdciz98WIQ1Fx
cN1Poiu4O3PdtBn97DJnIEOHbtqNdmXmB0GOU2tH2peXicvsuSIaA+3JydU3sbPT/VSSSDfMId1y
S5epyAGSclqSOBV3nKYQfUoXOiIU6/DfxR1v9ShZ0btCvzbVdFGvQOfc3F7oJu3di9JgyscGxRq0
Q2Y2rj32CmgKDCUBUfHkAsVO1r4l+VpY0NYfRFqg/qgMnirJXOf5qcQM14eGmZcH8mxL+HbJFzl3
vf0U0i/IHcSOSkCXvXqfK751t+/8tNW6PsDbu24F2cKIOlbpYqvcJvppBtKtL54tz0vx060Z/p/L
45k+9707phz1+BBSYzppVJNQByDxp5giPHEKXQ7A7FIy2GW1E7+uOHSZFQJ4Y98kW4tPM837Cb6O
pZY2x0uh2SBnAXMjS2NcKOpjmnVvIRFQWNl4VxUFPpK1NG5qc+XAnCndhVhWrOJ1EDF6AcqoSvCN
w9miRj3NoYSXwo8NOwHH4/UlOeGK7tyQ7zkYpDrdMjlRiCybXlYJ5vg2iON7bQrFvIPUyc611qqE
cFCprvsao+yMl/62R+3mmApD0BKVywn3gSWFcPEm5YrYSbJNvIqvvQoqzkk1zguDG6r1qvDSDGQ0
FZYPaz64qPPp5Iub7aKZkbIKBT4QRFMFifk1DqJUTOYJV7CM89O41lCwkbrHjL5atsWu1Eu+T643
MhcRiUSL/KmP3O69Yq6Ux4horXBgZMIWsjcS2Qm4rwPNKJZpUOG7zoOyNi35xKdxbabK9JferWqp
QrVm6DHTluFyW9iDrmK0vnRvR4NyOlpYLuwvqHM2WrL2QzGlwr3H3tkiKQfemhglvMuzDWaEOYxV
UyJzbDoNViX7yTKEC9Wx0165QYXGX7I1o7u39fv1OpSuSATWmZf7c6DbR1SMJvu0erwO+09h71Fj
pl5xnyTUkUz2NKmhrWwbN+OMcFbZbp11eTv4NSRZBWpxobbWvqU7yG66Y4+12Tvfj5agKeW0NLLD
MHYHkSYLO+VxMdH1Y9C8vcnV35+0v1gvnCN3Fgb9/uXki4+FLEvHYs172p5B02KoW3nSLig+w2UA
tpGA+oOp5WMvCsH8Yhl7VTwrKEbXvlb/oUFVNDtmme33U3pgdvGb+Qq9Y1BpjwbzcnQSNyEUJYlo
vWArsrT+IeRxY8E4dI6xSgqXO5DTbSlqcAgA4k3ycCpPLfLPCLxgk7DRI623HLCyavvnCaqrPQjV
81y5jPBqZtiJrlKIB4PMRXmEajzbHgzD96BL+Mq2Yl9TfCchs+dvbzy3i0Uvqfr4KZHkOF9oxIF3
mVO8w+rVq+1YDr5Stziu2GSr2tJEy4NFA+hI7P4bukMrKy7muMiT2iyj+h2LNfgAGyHFipXuMAXQ
l9hvZlaKtSqVyaoowButasq0VjiNaL0uyuUnX8dGxAoCTwubLdJ87w7eQF/5x/+3hbSG3eoO5+5U
MlD+Nq1ndvquG+N2Ge/YXo1jIx5wPd2o+CJec5BsOMgHTjEbHqKjT7MS6ASZvY7pIS/ZoA8Vd7l5
xQY6c7wtwxAQv5FBAfcuA9OtT+O2umzGMEFytboiduqE1bJA0Hfu5CnipgONzIKup9APEiJl2uXh
9/f203EhxVOhnHXtbmfjGSmexSC3gJohC6lUIiQwafVLMlv8kc3KwZZM/1g0woORPlWZoeAUAsxE
VjrMiZtP1bYSw8pO9J6ux12mrNaUtQ8IFH0OpJBx/SQ1uFIucwcmUPusAzZ76Z60QdeknxB5LEew
e5HGuJzFaUwxC3BIPoBQUexGuSF1BtzOZ3xuxEUbsyDrbKMQUZg0RHZnpOkDh1swcIatxppH3YyB
KVBogjwl+mWgk+DAibb/b4Bspfrbtw3V5POd7mNx1eg/IGEvfpyrxU579PBQIAw4Y3Q271aEusgv
penp52CQoZCrDEBCYCthYSeZ3IvpfFqRgRgVqqjOCyAIHY/ScWfprMiXEY6e/uRksTz8MeKFxFvz
s0L1oVt4DK96QymB30LHMjay7mADnvQPFnbCo2DDELF5GEromjmMFEQ1hduTLHOJqyPpTeCdPPFe
jbBGzBAVykHHP1fI2r4U134vgV6Vb5fi6y9aXbtVANdBKvgpVsZuPcRbtaLLISBhMEBHaijm54d1
gV/KkbNaQ74rw6zuBfB1GQkPcftt3pstsufanaYwl90ME7P0W87k/OTa1vnRUm1BTj1rHbPMDusd
S40TKUqFbirncHYC7Veay8b+E5rJjQP6NqWtRiKxu6Y3B8smRSgKFPxmK50fR6A1p+IO8bNYCY6u
pQ73oHPKN9LXrbPi4qIco/RRZia+Kylm/0g00j6s+IfM/rr2rc38WEgzZNZ8OtwaewHBoOQ3pG26
icCm+2Rz5e72crJbKem6CUntQvKInKGWfcg9qYV+7Us2Ie5KClyKgPKuqXfvbtGJp+FqwgfNNGmK
sQ8fOO8Cg2e8Bwkx6jTuQQ+eVVUfNubjMU21RPpSINZukzWL5JSPM6m6PZJqItg9WOuLbhZ/nXCW
iF3iFW5NIaBUBk+QWyhEsji7f1KvLaawhBYfHLgBtjTPzFXG/w1huHEFT6AukX+WEvfkoL/2qE8W
UpURudAjdGYdVnmdRQ+z5hVbsga9Yt/HD5TJVX5H7HzRkxLbpLW+YMpnfZsH1cYgMemGhGaz7BaP
2lxAuxKlfGxzcaU50H7iTaES9UKGw6q3CM2xtjcP2UmP2LUIvDoaKuAqfAsH6LatCXIUg1GoPvpI
OjAN060fExNYYf/5hg2Jw1tJT4SLWTgQ0M8WylBCLSLliNH6Akw6RDThTBPL6Pt6gKoIaYEDveTU
ojnWckjLWbZR4uv3nsS+jetaaOBTHj0nRm636eFae5GZtqljahx7aitYXDq1OYQ3Sg6ovoLZYz9y
EGliiYdENf4dNe7/7XUzDsWUineKtNz6hzvWP+fRt+q1aW6U/Zh5zm+9OMKVMssAR3L8fzYATcUh
sd5HnI1o9alaYZ07dtp29hfhdr9pV+bfbMv3IZcgmnLYcaHaS/s51O30zCKc/PTl4XgrcACrZS8I
arHWjNzYvgQa+g+kpElVWVOITIn9FSsYT1PhrhfhCouS7/841yueue9JasUevX8wVd95bqlLGCxn
EIiplaZvBlNPep+xykIEitp3lBeUvT3kg5JjCOthGRHhKbT4l/wiu67KjspcOnw4UiqUI61zdY6P
i9xBfEYAWV/rL/TaU4pqSzWrsGHb/0BKErDbC/9lavwZPdv5yLxyshsKPdVXh3Hl8W87R3KzenUP
8Pg5q+BzksHxDP59I07JY8Ocs3FleWH5dhnHbY7TxAXRjUA0BkVzu7eKN9cBNNMG9TK8vxgc2/01
4iJzbl4paLj8paXhHU6Qz93epyYnCyna10AaGVd/cNdu8bgQmxtFP0BpOQv3vD0V5DlWkn4u+3YV
tox21Ux1ZYLt+IzxKg/bBiE6MoZjZHwoJvKK/5A6bKGJJpKUa1Ig/Xm/WmlyIPUxYEruhoGO0cxK
aNgqyerxFhUBfOObZ3SWraBnjzpHqMuWYNjZcOGDWGgnG5VwyY8ijHomK2M8eOjLplZXLoNYcfTq
YRhAAAes7NGfMHoszETxUUs8rLhmhIyGZRm/7Sp6tn3cEKNfrFYtaXvACFZSHfc7KYvEVsrHc+f5
nCLtzGFoR5xJy85twMpQpC9eska1ID5aM7LWFPeFTmVSxyaClSblV7GR1os/kA8FWgtNEaiffXMI
oQwf4p1RpM8DHd8SgS/qrDB9n4Lr3h/kxhttOhx5MXouWPNFqUp73oTKtN42cnxeUsW2kFRrVw/S
A02JuZsbf5f4/mdK50JudACRnGL4UVwr3QI6sdKqFriDuEH5dva9MIxayZ7ac5dfplOcwGiVgw95
QvqscEKA9DAYmSF6bQYPEkraKVFCbNlpHteh0+a4oX4o9fCyF2s/YMEcYLrFe3LycE/d683jUVs8
XLZOiz2KnWqG2rIq60FYgrncgTLLJwas3cBwoK92lvPCGVz71MkEExKZKMepjvtHr0Tgl8brhmP3
AmK6kxSYs1ppimgB3dpPvtSomdw8a+UvHfAf2/BKaekm5QHEzB2DEsFqse1PquhQ4+Gq1BbsaSMo
SxP0PIHDtA8LV3rQwQejWUp5SZWpJekuFNfiR2LEtvUpyeApGg7SHqfsv99+8Q0aIVNkqXPSJyeA
mpDBR8N2rbvBUHOST6Be0thzA0CjnmIuns5KGQXk31wjDyJPmloTjg4MgTjL8X8Utn0/TS0gh6Fd
eQRIJxvKrJdg84jhRfJSoefQhSRs1vXg0y0fYdzT/MKZ+HbuH5ZtEUiX1FUVRqN1HPDTjohtMYBR
HF12vGuj3H3EUTHEWV0S0/3O1ZOKggXwVISUXvvjy1bAqsoNycgTBgxjNQv4RH0WnKRqAGKVQJFM
f/EKB6w/GGgrQnFNVZpZMv3KtUTHaHCgqihsUX1cf1ihjyZELiQ1MkOFXrBm433/7r+fiExDxT4a
ZT6bcGI+TNBxpO8vToLmwWvO5rs0061lTCMRE5m0pZPAYRXWPb182ArJSeWrGOsUtuxRnFVWWy99
+MlfNmSJEsrmyY9Q9ju/0gOlin2Ag0z/nVkny6Ss5ZqLvZpyY6IzUvq67at1VuVUgGrcJzyg+fCU
ToM3JhOyQQ0t9GA8OGJ+aT+ud3Hd8HrO3jKfyxYIx0V8c2eY9DziREuVA+bLMPeaWeciLR5uJYCT
elPkIwRVMVBsVSLQjok9pIOPDgyyeNTFv/Wl8B+P/w9V0LonGKGn10oNCIdGl44nLWU5of5hTq0D
f5oCNrtL9OAN2BalCHp+sWqEouoYdZ/fzma1mUdFF9rMlhjCoyzzlx8PdAO0yt0KRh+11p79IFQL
xnvxPI9/1mGKzk2QxlRoo2UmpMCWDemO4xeH2F7sKASlrYKd0V95Zsgf3qGobrFhClIVVLNEu/tL
b7ojSHA6n0FL1vUW6BQSfe64Wn9pxoELuV+qX+3OOtiP0WSZ+pamghpiOtSbS7QHwyUFGpjigloj
qCgXIKDKmibeBEXDzdh/7wnnHBUctB4uPGDauJn+jqys7++puZXsK62ulZFBhMxEp5++tULlI80Q
W2Z4hiapv5J66qKT/ejcKkZWAJvMBdINiQBCS5nA2RDhCEe352TSFAhwVmPsxmXoYqtO0hDeNFaX
SgkwYMwCHTJLEsIdZckFRE3D6FBOJzQkUI9Y9eL4x8HGCMjZpmLpYRuLBnXOapHdr6ypioMKf87O
+9anpTXEqN9g8fQcI9gj/l2snJCrww5S2zNMcyTI5wQvfzIthe7Pu1D/tQrOPRUx7Fo+ooxQ9yAm
v79mlVt3YXiAlAP2Aav9Ic9pY4Uw9kvqN8tIzpYd8D4F9SnZfV/+KkKPoHHnSfH7YBxVq4xlYqQg
H3Kn9TsHOYM2UgDDvCpvh/UqdZNHB5filnPMZICuEjMgBN04QRt+/HMLhVZ3xzpInRqrWczacAYd
UDosNFyljafVl36tAZHVdXpAvoEGpZbe2JfHzjjSAbFzGfTMAqA4KHvhV1yU4/fuFa7IyhH8ij2P
N5YwWbZV0dFJzvncTO6T+ADKAjkJ6qRvS50/hTMkuvNtf2Y6454mRTX5BOATyqzuSgR01htPPUQa
1Fcuv7/HGKxUFQUgLLNf2WwJ7mDU3VVfF7gyrte7xYkI7I8y92jqWkNdTJX0BAZVJ5Bq8OSgfXZR
gm31ug5y9q4Jf0B8ws5t9sUafHiWqLe9sKKHaLC3ubMTPep2TwGh9OI7VUtGwVlL//TNfAk4zCDs
JTO5ehqY3Io3lnKElcByVQlmI7WI0SvlpWoM0zFjd3Tp2SfZN87zLL8Up3dgCnrRnlIq0ba71fF3
Q0ZvJGtiHFSSuaWbYB/p831RJJnOYme4qClFGfJNtNSYICPFLh1fu7eq/jW3uvAYLZnnlUw4kYmI
lAuySKRkNNTkY73/6I/YvKZ++uQP0poits5Oa2P0ExDp9kwTtglghWa0wjPruFcmGbg4LFmgypkT
uRjggjEw+y4mzuSskEm2zf6zUh21bSg/1Rhxw3cbosCbmmpbWJYX8wiCVP1/QObfKwc29FIRTxYR
crTPwoSaNtNmvg6w78NkxRrSOPMH8nwy21nRRoiwyE/NfQQAO8sbMyxpWH5AmUlCHP+B3FXMu9FC
tlJE6t/9tKUSURkRDAfHtdxCtYX1OgXye5n2b9Ay5kRyMuzyWBo4XK1woz86M5eNHCVQLJDIUEze
cORtPFbv16D11WlOYwIHsjYV1tWiVbPMwy2L+haJBNEzdOZNyqoc2Qf8EV9k1HbSdrrgxeoHJMOx
fQ6zCj0LrEygHc//r8+pj7+WLQr3kcRwwSJ+WJOmQHucK6sZHC6+kKctJSHZKICEb7O+KAg95wsi
hIeYWy9pabG7v5HGeR3Vc9fXs329kSKCCByOO4AQ86yl+XNzMCdxcqEa5/qiGvlerSJPANveUdMK
TNNxe9XEKLVSS9fo9FkwKhG8xSHYfQQO+y5MzO1dPCibE3/Q8eCX9soJAi5cRPL1HikXg/Azlm+W
tzpJYimAOQqsnr/gFrF4+7o/Y394ES5SwNvN5vlA/1cnS97LSdvwt20mDAYQrFJLAz/HmLPTru/X
cwU32A+rbl6Tk73aRedH8NOb1g1pfujx3KBpukEXL07gVP1OwllmgIgw5/L3Mb/0A8+IFgb7Ni73
2YvNtuyqwH8mk2+haDaPP352vZMp2Hqw/hEwG6SZeGba0u8IV7TWqqd4PSWqOVbacCGlIk5E2Jka
OvZbCdLizeJCrkbgxUjBhk7Luy+u7LjGGTj/JibQdEaEod/l2KBeSMHFHXxoTzakh1zh2b0f9Gvc
9dVonMWODA0ipbhvf4AhlNd8uCvTlHtQgu8A4JfGJhcUSL5oWlqBh8atv5VjMzNQt8+rFt91itp8
70x7FSmagwL2RGfEet+R0TAWxj7rKOWrhCdt8/RmmfInjXZ25sSCfKvDVU2/aHbzzRTBxmq8c1xb
HotN/gsXQ/IMLeaLYvbhqdOMAulXGpYEZoUbNMBDt/14KbHE+c0DtN0TTF1rpxGE8KfeTteFfnhJ
L/2SgwcpXA723PwjnlV1++KswzdwWRg9kWWhsHKnqMx1wRF/WiZ0Q6cLLBhSio7k9GMCe0YniKiv
EEkk565iMUkezclZWXDaSOMejNPkIcHH8GTj8XNkh9f3pxG0ViaMwNXrFGS/GyxjidyqHKLyqVe6
//p004zAt0JW11yXMSEQtUgy3vA31bSdxOdbPE3NtMA95KmXdLQrcdiErssaEZo7rxgsgtqIZbu+
DY5ksOUFDKf5Rfz1o5kOhqDfeETJGKCUrkU3VEZaVG96mSoNHCZNOY53hCSsK3YW6awylQ8aIs4m
H5dwdzVp3sHRNaDCjmHrMdexDYVUPxDXaQp4yAYCf50JsysCorpuzK3B6/7DXfm7S/YSBB60fj2A
IgMiFdy7tJNIKItD1gvj/Z7SoeHQhvsaUmLbfk7iJThPoUUA+k+YJVVreAhAbqylyHyx4sbgXoWC
BKcBJyqlWTUPb/zXzpQ8kU6LJNIc0emKUpH5C2NU9YkWqR42NyUmP3yUOq9Otk4ij86dWt6pAlVA
5i4QMi/kdzWSrEUfr1cDTgCujfd/hsBxlhv6UgZj/OwkKL3DGApk0MX6lf0oRIPWz+mwX8F/vyb7
yKZdYSXxnTgqlbSR/3/4okdHuGlzYwDigL69GQSFfhmD9hEgtVnz5JK5eLZYEPvSCZxdT890K4fA
P4Wsp3nthfVLRd20z9J1Zx9fswjHrIzEMaxJ9wDGDl84MHHknNZdUHATZOT4GdtDXw1ta3KaEQUu
pwTuPNjDPbos2x7hL/OBtpthtSiMKWazJyQdr/cMb/A0S1eBB3heCDssPbUo2kOJmVvKc9kNcjRD
3ewzBueqNaS5vZvSjrhVll4yzTgg7s3/N2uTjXO/7Pty4TgqwZTeKN0aW0A197VhB1Qc8e1WtwYP
gd6tds0hM2eiOux19my/gXTpK3NqXOrPoKP4Dp3gz/fk7h+mZCkOROX3okH+x0a+U4mT+l/oRCgv
mHW4fRRKVBvMJZJGu2PPuEV7RMv/+tFo/nSE8uj+bsedm4HHkxaF71B+E/HX1eqVSIBGOwOVw9tB
Cd/azVTgpcRtvq3/6TLiX3IzdTz4VZM7gPNsr6ZbwDmcL3tp04yB2QsVYnc22depfsBLp1qeavAE
0Hu+Fh4WExs+93o9wCv/iLjUQ10GSLwAL9SFpbMYhekV1//f+mMPQOSle5kFSJkjy2KX9ghD47Rl
Hgyl7IHxln73iOWTbLv0MArPCJlz/ZHOPtiysaqub0K5FZJMXg6X2KFqbyobUn6901olz4J6f+fe
x7LKfxezy1pUXwFmGW6O277vCAFLWc/Hsd9a2WfSsDSp/tSdbgNt985K6tDw0Crmak+1FI0UdZ0r
jumriAi41WlF4F5CYsRaXjSKFGzcH3ZZdbI5qUUk/W+6/x/MVkGK4/yx9m5QwQPcwcXnO40YuQ5M
uq1fi3nme589RsY4eHyv4Edj6VNCQ9NMCmFqpC0Y0RtnK6YfwXt4VWSswUDZUiCawmoDl6af3ioF
rXjrc2fh8uKgvwqDNs8w7TZ4nsM0wveY32AokUGOEVKRJlgkokylEr8gqHYgCA8FBJE/GQCRnbW+
D9BIdhrP+bV5KxM5BUm3BWH1vHq4fgnlkdBCUEtg2ap0gTY4iWZJVlb2Y2lfxpptQmQOo7OaDCdZ
VgCDIPL1c5M4FLX6n49tpkmoVjnBd4Yvh2wKfv4KNgRJsaIYcyBVSdHGHEcXVj58g890Egit0iMo
YVrDsE2IGRrR8sGDrwV4J9D827UKxQMFODQc1OSqhpVIgxqkzz5lYyc8a/JZOt2bkMk5cS9tCkW1
Dk08mKRZ65yhSueW8u0qwb5bZyeWSUApkWrK8q0Jh+k25Pwyr8fveCo9/KGlfFlcM1JscPbCBnxv
X1UlmJwTPUYuLlNltghL0YmGixpmJe43RUvx45dg8MveEisB6xZsCMSzY/XtO/+YR0OyWmccSEm/
O4/aIxIoogBbNEMRORbSIp0SwfPl5KShua8x2B2mh8BtOhzEVSe3KGUTX9ugL6ZUkC8DSkREpQxX
JxU+YgGZUV0KzyGkdOAW5DD6lg4JEHzQkwBrIgxOI2NTCODpxWd2yC9PaDXUBmGNXaK81tJAhA0j
i5bUKNirY1spuLJ2D5CuuPqo75XsU/a0muSbk+9b1o75r4y6bRXAlwh8De6I67RwILejOMWSuUpD
ZBbOdztGBxlcuzdYXjzaB//K680Pufixr9RDy793VIK3WrXe0RLT/awwJ8uWE2K2xiOLRjU3y8NX
OrgnNNls0umbYQtxKckYa/cwAKBR/uLg/lmDrHLDGo9hYURua5KREH1GviWW4/mYPKAi11nJH0cf
odeK4N1+prycAeIGDeiygqxAj4bWjqkVxCQHEzmF0tPPHXUmor4TC8X0megE61maUqVqjyjETm/U
/OsYQM9NryhFYo7r0A9job1CDmxH/AXOM1+ZaFHvpZuVu2CkZaYqdM8wHKIjDOZWtgLrkT95+/sN
uGBNfOodTo5i1e9IAvFPO8eH6VTY7Bw9mjOk4B7UvhXzuGCtF07h47BzNpJsrVlKk9ICa7jqJwUN
zmgJxzR9+mGoKhrVfRrhUamhT9QR2F06+D7e1qiOTZwjmc/ZFC/74u4u428AA6UwYggCn7UmxjTV
BE85Fy2D1oX/yItCDWTdHJKELd3et2LCzGLHy+6jPuUBTJlp0Rj6xUMjuj5NrrCh6SHYlmTLpLSZ
4yHCBxeNmTj/n6IZ96Tp31bekxUndS7XNqlHR7VEDtuTE8y0MOSySPDRMrYrr6+TsWg5CQB+YpbJ
ZAaI1/VNBmXxxNvp2UMyYJWNSG5WjShkp1aGJov6jExdVPUkTyLYWvUZIkOMeCZDygmdKOjiXjRK
Sknq0eyuAhURsztv3JLacL3/7C/U0f+RxSDurfAwqBc6lRO//JCluajgrT8LznE6HE7qhAgtm8ga
JY6SKcI/pykZpzmyxO80dRyRax69Q5snAVnUBD3ZYKyNqSK/d+uQYTAMGy8/qYUUMWH/z/b71puP
IpWIpt9rn2X7Z6oLu97hrICJ3e6W2t4zJOKa6uMVm3I6DSqnTtjwtlFZvXoM/+6KyHQy2pQj0N4g
4uy6W4JRBSYi/NleL1QEQYC+SFsn4McsqbT2kTq2LKN9078UXPQdN3mDBNGvCmXlViQ138kgKFTD
ARHhZYsI/lBDKsvCQo6/7QKj+Y1veao92v7pK27uTaqot/S7/e6/2QDyzw6u+K1FgodVYleRXWL/
Kz++1LLRx7nstVAukoJ1jQxJ9IdmHTDrWIv5P07Bl+LG2j+n0pdSBeOVt3F/eRqTesh4+CmuppBS
MqlyeUj12R2aX+RQqF+uPdcr0EJaoWVZ0lhIB8zu1z/gbBH3xJUi0lTnIqd15OoKD/N8gGno30Po
CgqrK2iMiTBAJaBXdQ8FHtPTNxLUDGHZSubH4L5HMHastTbI9kLCAmXyokhiEnM2+xMhmWEtxazS
UPcze7+VCaxCMn2490+H4Ls+sRd/PqRmLINt8qZqcr0k9Fr3JnKHfOp9OyGHizv6LI0vlHJa6mQt
GZ8hCAxgqWdM2z4bi/rQjVrjACL5EoO3MMACjPFcAZLPUAzH9ZlibVrDpz0vQvYMDD+8JjqplLZ1
7xZy100Mw7uVQsW8Xr9qyrBGptpaLD06sPZBqUeGcJi2RCi6pYyN16TNxF7fmWAfj1lc6JjBhcDh
IqsBAu1X2hAi4EzEu9n2IqSpGfM5awtNqSJgAaBDx4R8Qy1vqwlCKxz3CAz7SE+s2KiiKaLyotx5
NsiyLuoo/H5GIxYx9IlzZxZrI9fHPOnkTrAKbp3nDADsv07cWwP96121pgLHiIq8jB7HsxQeLnTw
/L7+oZskBD/XOxXp995cnspBypWxa5r/klgwaCZhoYrrg3hdtFhGkCLxwNTw9OGHPhmzcUCuv8mM
T4KWoWJ0BQsNky4l2z4dQeJtZs0pDeBDbJR00mnm5hsoEt1eoNrH2DvDSCb9jt18lmE/SjP4hrTO
2HkaWN8fxljuJph7QPm3XHhopoUaBQl9Fo6+Xt5kxoJK2Ttds1U9uxipJJWK1chewSU4lSZfX6zv
wYueluTLZnXemOBloyFOFvT1npLQ5D3HO41CkPDU/jwl2EOBHEZBFlJyru45QHOv4YO2r7r98Qxv
K1WBT1xXrVkLZWbff7u6hkjEN0XP9X1zhwRsdUEeDISCKrBBkBiqrM70K3FseQ0SD5n1x5RfVqA4
XWLHM1rYsC412wI2+PaYJKiqgLxA4J9MM2mQ5O0ouaYGOsUGInF1adl8bR3ffNc31PoNELhEp51D
IvjZqJDm66jiZStvWH5zaTCfCNA6ZQtKNIl+LwrWnbLc4YVEIAskwueRdyiF6GklHO62Pdi6hNkp
UKAC7uMDSsizhj2i1PLJkRKmH6+knOdrEi15NkarbdDlqrcSZjtUZ7Am0otIlY1BewJRnk12De70
bj7DXf21u2PRm/2eafA4M+3XZZLve8miZHdAVZ4N+Gb5uPA6VV67JeBya272DSQ1KRuszD2BJ/cR
dFFLPo1BmdSeYeeCwBV0ZDJsq/zCPQ70YzFkXuzBItntykpkGBaXeLJwC+4+SwVwfLfX0Sv7zblf
Fh0QzEPzw6mtH1lbaeZFabf24iaUK9fFF6/u3yCEMKiX5JYiTkbuUJgBWwtt/tnzCrZBHtyd0sJu
GPGhQAMsv5DXZr433fYHtUYAYFCa83HTeNunWB7EIJHFiN3MB7uH2emzDKZG7Hr68roH7MDhOqce
ips7S9mkqrLSDV7e5plPgxLOlzlPgnUB7ienzwe/X3WgnSBAmglE5zLlmdTUtv1dviwsqqv1UZkh
omDSahD/UPD8xvpt/MX/DwIHVz630NiTKxeQLTfC3VqcAvgzkuf2reWXZ6x1K2egwidYoW0TAEcg
Wy/h5IaWfiRrXXxVzIkcFQSbGsOd/Tt4VnMDipcX8UrciJ6W1+Q1jUjSRkf0mocwrUbP5vpjfK67
1RxQ0pTPFfsXXm7KF49/+3TALvnjOZBcqoXYnD0ti9t5eMAt4QkYkY8VrDh9+CD0XJq6hxfm507D
/F9JVQsk7GvtrSspwdIRznrznAPLaiSw1SyV3kNPObA8/4n36EyvUNg/j8sRtjurD6wa3Vs36F2F
uExBbRVVoJiuCNgh3w32Z/ReB5pqKG8oR+XyXb76s1ccmDlwC4R6uSb/i2BHFRkGOVw8uUPpKmc9
M/9neVZwgY/B/LxF7Fn9G1dxber32+oyPrna6nMf5p2WJB4D6/S6ffXRAqJmWH0982N+5cM/uvn7
+Wm6THa+4sjuRG/D4hwewX94Zw+AWVqtmp2HaBCyrwGoVf78JpTqdw50Cj344F6CxzihGOtijyxx
oHZVxK3qkpm4MZNOl2QAIXlxOgEt4002ta4uI0c4aiV5Iy/xAvWXfE7j7OjxfqD2HApNSY8//ezT
8bI9cQfCxSq7AcQDwrWjlDe9+PT/hMDwwgZZwcKEXcgD6HxaxX6xJH857gydy1lltoa5CfLhslaF
d/hr23Qm2UGCfnVJ+BXWgoWdmWm/VLiflkHG67qGM+JORAMMJgzc0Yw5xoLp2day0AKZPogB+oXs
rUILbqZbSPEvmPPNFCAiidHY9hf6x0zXrzr0D9ZVDtD+dB7opAY4J4clXHWd/HZtQOrM0tSNDm6e
OpAG9Px3W/sFSpCprRD43/Td0MZucnW2i7f2wrnwxh4MxuOmenr71Uj6tobgCQOEivP54bqFBkrD
nw/2fAK7Z//9BxSpq3VbjK5Yt4ebelBX1tZRri2nITvd+SN12LIoV1zaEHLtI36I4BDLBTUxaVKU
Btc2NvbbO9YhRV293dLIBR5HIjF2g3uqiSunVGesLXmL5+boJh7sqi/PvfzvzqwnUguSyZpWkxWV
F0u+an8ONlbDDqqjd5RIeXAKceVdVE8TrrKgSZj4r222M0fKEH4k9zDbKHS5rTztZgNyKMnKQOHN
eFwF7anzKuDcTSSK8nBlpPB8mBHwVDraVcxwYuSX3SZ3XID86dZdmjVqBFoZYca5skNJ+SnfXoVn
9jHFBfkYx92Nucv5DXaDPktfUZsM9CG54Tlya+2NJ+7BBSjdixdWrbqKKGBnOn6pJDvU9TW4cMcG
gZfeIZBsKrQiVO/0FLjmdDpoV9AOCXjiUiZUtIQUPRSnqq1lnmIueWTpZr5yy2s3+bl98PHgFs+8
pMVqW+yAwai156WEnhc4VsVBPcVx+i1Q5621bjs2WOYK7qp6PuXXeFsHLLe1+9Km10AP8HhFesSZ
M/I1kl0NSVe22TIkYvTRtPHoEMWeclmexa7z8ET1i3pnNCtq4quog2m4NDE+sBaJXkzu5Oj41lt8
cdcJ7EQCzvssVLYo7wV9BNPWru0zeJOEjb8s1Vb8XebiJZ6gLUpYf2XRLs3dNf/2P399JhfXfj5J
Nyxs2iCPHIEn3XCU2UkuTXHz65vpXZ4hIUn/zkLBK2hzxKsgVZDM3V+RLWJEhtY/B7k/Y/t54kmd
IBpoLRa6QDWxI3iRhx3AH8kAWk3fAR3djxpPOdgTe4Yz2K/pASYdv47fg2SoLQ58uqzkrMNYx6B/
VHJOD2dfHr6GYPr+glKS/zQDEwsaUMCuX2jS3/swBe2hpyVePMQ3N0IlGzQ0D3BHZIpRxsCyeKsv
jgYVw5+cgYLME20heILRnQMSlWBtMXrG9lvG8yJrrZckLPE14g8PqZj7PP/0QKIXCccHXBv+t//Y
nkbIqv/nOA4cPNJV+o++GWqJL0Qp4/XjAAt5EZ13Q5a0HZDbH94Gq+BG2jayPnhgErre3aT976xA
zWzloVrksoa0WHzI9gfCrLz9WqLmvdl2dL9wD92Tmtkq3EBdtZ9epGQDbkh4NaY5kkkqts0XCOy0
pisS7HcgAuJ0nqolta0uVilyWza/PazJU07aK86W5tJnEO6gMWbR+RoIHZsG38v44hgo1nVQEC/v
3w3kGYOwiB9JVLLAJtbV4hpMk2uXpkBDrndqgXiOU/RhXfo9TscxoDV1scTapzb07eXSEE/nH6h1
G8kTszgvB88IeTJaVZHIDzUrr54e1ZxcGg1ZwkAWbab/ljSeqweJUpi4jEhnrD9f9bczbI+fhgxo
aijCDwhsNCbybAQtDGhhv+KS8pY5KprtH/Jdl+Tfg8N1IqcW/TF/N/EhRJja2brd1QjA83GjkoJw
dXoCRmsTDiyAG6XjHEsqeQtHX7VGddEntRqQMo3eZgHaRCCQ1q9qf5OLr3aEYbQdCx4ydt9LTadi
hXu5FVQ6kwuxBf9ij6Zs/p+ImE0P89uq5ReuMzds29ifYtIsXkVZXaDMgz5Ybm7B9/RhK41JkaAk
arQZLbAiYJDRBpyRsh+qtV8jFFd3tfkmMktq1Of2z/l9/hBCSVx3C2DDfHH5RRkFQc2Lu7pTKQq0
tvuxx5w/lqv1GAF4wD8Xz2z0I25nfcMsbiueviStsLxPPk4T0hdpRnR4gRgPsNrkMUCFsVmX2SLR
e+ePbb8CU5NloVTD6FKPJE2loQ4dQIGO3KV2iquUf93dPDF7b22SZwyhuwLuNJrYmEUNB9Spe5nU
WBxENLCi99bvXLam20X3cOQpjcfylRvYtjTNDXS1STvp3ex37sXzWI9d6/kYp3413kcyNpBPbF1K
TUCpSpV1TSSWzLy4kYaM8F/4Qxfx7NLaFq1BVj4TLwioZM22Jkut9KUDscY3muz4gTQASjSXs3V+
jt5Sie9xWYJZTSwow/xJCqYCdCfK5oMpymJW3ht3bBTHEhGyKyqCsHNt8jEQygdpmClNXtwtBjNR
mP/+UXrC2ACAtG6htdhDAkzF0eXMN9ZTjxVU9Sm8XFzvWdAip5mqKtIT5CpgUGJPrtVB0X+zrh9N
wM1VMAP5ZAj6ZUOp0aJoWGhGsH13OincBbg0sgFhPLecTyN3qZNTl7DycgEzu2AThGz5/exBP1Z6
oy5YXPfbfo8zlbWolKfU0Hk3o7KiWpA0FnWzeOB4hzghaI6m5FET6TF12bK4r5Auu9cUqYBJAgLr
rRTRZGcDhLadKpc53IKl4IAg08x7ylBFLQ8KVjgv71wijgD2u178+VmwcieL0suw86g4XJoFJMml
Ss6a73Ss/e/AL5J4r9t4NLmbh8oTAZmmYn04FItE3nli4ym28dY/Q96A0WZEs/NGe97G9CFQYpDo
TcoCYvvQfNP/1UtXBlhtmExXyuE95q2iOk3UAljjQOhMAQ2rCBnY0mUrWLThBcwwl2CQYkpU08Bj
rKa9OvLgl3koare1+NWBKzMQnyCTcE/6yOgUBC9j0wqsrh3pMrW/KHYLf1Vc/NKtWaIEgrV+o3dJ
ceIyTzagrfLCC0PmqFyBba0kzqHRmLMx4LpJe7ZiCudZN6c+HDVEsLN8glZnghJecd0gmDCjc3Na
ij93l3dqDRDfaCkBTQfpq6r58MDdUoDK5BLeK4qk2AMvwD9q61x8f3UwmzdgsKo1QldUI3RBzAsl
7Y+HiuSpuiUiBrJ9/zyIVWjpHeRkrij+D70TV029/oQa1VaLTMVaTOOe/2Y+kqr2MyKvpq3x2j3D
hHLdBLOLGi/cteL4upthEzDwbVO9ilCrJ5P0/taVxZOwsVkQR2H/slIJSbwxdsRnff7F87QBEF+3
+HNkxEtLtAPRUoM1wzgqK6aup9+sMH7wlpVmu7bhkD6nZ+ePHBSox6yBH8x9G1/SbwRsnKrFUHWq
jPx0ZKvOFfkRn1Y6DstgZOObLmB+HCRXWo/xZtEP5xL4dmmuFkoMjZqhWaqFR5KBXYxusLB5b1tt
hy3W2EJrEsoAK+8ObCXNrWSUzXXLiUknjSh3BYqNRlOw6fLOWGRn6YSFJ8LC5yxp3cuFdDbL3AED
3vbkt9yMXiy57oCvM7OxIQMVJKHnEj6nHlMlAlZMsJSK/xh5lXZy7cFdGjG4IQDC4G6iQbaKx2Xd
XrYj15y/h+kT7OprzDNG+tJ3PaWKS7ne118o0YfeETbSvuOUKtkW5QxsxUdkejUKb1IMUnBbdzd0
0d1FCm7Vtg3fg4cX0ewxZZmgxIZTLPUUkWT9y7yAeQIIcNn83+8si8ZE88n0IztGi0yDt0UCtlel
8OHQDyOhmL5jFaDh2MZsIz1hEVbL/Jh8vVPFpBpaOAdFF/borhOs/Na+WaLTNGwccgK6qR1j/Wi9
1cgRml3iF2esX7v6ay9TOEuqxwFQ11uUtKsrTQg6z7dX9ws6aiYCOC1HZQDXUcA6OKLumpjJvWFm
EDH4GBRTcqzASlfdxH8jb1tDc6qaanDqKS31YQqIVxl647YGvTtYv7yWpAdVx8/+USEp8RSpoz2Q
q/qZUTfM836lDOzUuT//ib6I3gpsXM3dGoZs6gM8HrnvIlEYkFpDL0ED5aG/PgoZOFC2VvgKbAo/
evUruThpMqivU7HHL7VTXtgKX+6lOSlYyaegg0Vdf3a1VKhP0nVcMFO7UlAyVo0iOEq2UhByGt4y
4j8lc6QsgJLmZiqrHQ7XSG7hPU0DkNkvwWxu2T55X+9TLhQ+1VMHc6hd0tiRxWIzj/xkwkfft5Tm
pOdzbySliwBsC+qJ7CSxj25K5E81EvEyg4OUEpUAgtQKq3hmq6G7Nty+UjZrZLFhe7myKGz1J5hh
BjjKuMUuCe5IQ21+ZPcvx6AP01dZdMAVVN0mZ/2Wzt9HHxIZKt8GXoPFk4wHm9OJqbbxjuPX6LGn
JpDKL1iQlKBBHJLsb/gFWrG3puhfAbiRP55C6oj3I/CKkooAjG6urZUzw+KVOACH60jlDfRuPY87
7QntMiqhtmz9DfZ8MXrNSWL+yEQLO3xRiiZYM/oJlsPpaSjtSEvGnrQIL+UhLDPl1HvHA0gBFLvl
4fr7ZgWFB6BP2JLYZYSyknc7eyV2khaPrE2oGvDceeo0TdSODWJpT5VOgK8m5yqWQiyB1fh25GXQ
IigzuQZ9dXfmNeaS9l6fTj9Dzm+bX3WZF5bFSBR8MaLmnWJcld0N7a6v4jxSitOV7BBhTu8HFPkU
hFR+cnIl2FHDXHlLGwaCwjQDMxmOoRLACtjibQwmPnK0YDiKslv1oeuMtSI5ds1alKbiB+PAFlGM
33FHpawZ8ZBkMjCTFWgJiUcOvb+WBqlG8oVbcTkmDCzMB/xCL3GyDZ+bEsmmUGn25K4eTgTFV7Y0
8M3zr+N1KKnMXASUPIIaxrswwzTWRsJrGI5NTRuAYXoMln6ozyRnB+FsRwH8QiGEvKNwpRgLMt+s
xyOwZWmSxV1wWvmYIWF7D2hyBmV1eeSR38fVcXmV+f/tVQn2FGqghPUJNkEnm60417HS4DPPeFdu
rAlJK/eIosa9i/QuA3yomf2tC4FOIKloeT8WpLo66GwHFHxMGhBJYgmDspMzFw7/zdIGj07+bFVR
dCaeUw0EqcQ5WavRKMbrimfzs0fG5tZs9dI8dB7KolsQl0xvW+ty+OySibQtvYZQgkwVkGWjaGUS
N/Ne1Ar8nij/H1ox2k9E4r8uvDeJxHSLjshHciM192jRlhsJ5XSCbNe4aTSzUlnpBq5N2Z0tUcHf
0UgaRUlqM1y3JVWEauzhAGFGO80UwG9DGNSkxZ2YAquY/ZQeOQxh3nvOdynVw7L5ZydQsFFg+2Zy
bmjl44QeHGHP6ZDJlU3GB+HzLmsp6bp9BzB6lDZRMBKTGV40m/Fk4G/d/g0pfh+MLs8PsOd1M1Na
697OfPH2+wPflmPKUyWVipMX9MzWcMfOjuIcefA8+7R0Z5PRZJIzK//Q/XE6UB2QywWbd76oPbU8
PW5INWKVQnt1nMXTiW2GszHRDNRKDo9KJOAfF1kIjUMyy8hMyrx/k0+U253MnlEuoEdQDYtHaRKj
Kk3Ke8UQnCSrDY8Kd0gWSPL52H9ar2Ej+jUoyqeH7UkwqalC0HQmR5WCR3txhy419tP9NWpWgK1h
2e1p3ZX4ULGbTtV/YJBvxzkJRWD9pwOO4ld37/fXIcixwxhOl5oCUrK3lH9E8U1moBQhBWIpsHTC
xH2jLtOPPUglKVWCbF0Ofh/f6X8K7NV/bw5F7lb1oECihazsPMFiQ+FD7zIlod6VHIXdxMN8LwwP
L2rhZqmL6+NQ9Z8gaFDVxnhQUUpiK/yuU2WPDHWdGEjQoZUp8bbq/OZF7MLFGSw176Uhc6npTYEq
+eyhJqlOHIbaE2kMmPmyTuToWnkv32CdlBe9mqFqoqQkbpPFuncZ0NG0vtLL+D3LZgKZ1ynAkbNp
mF5YxWJXpzlyM3/gWVyTUnWqDDsNHXmxo1kI3coAuMvx9+qa2AgHK9pBfUBiwOZPhD2JCh7bVhbZ
2urGoGAJ4Q05fUWp+MUYSmIUGRN7hHue7AsbUxfHl1PAfFjLnsGTkduboYajHzkKj3s8RRTPPjfp
rEGR048yRjRTlp1fy1wk2imXC9g3c0RfehLKN7LrOZ1dwZ7yb1vr+ijOrnKWBHdwF9kxC8UxYyP2
qqRcObhB/PJf1Rnq9fLi5uzGqzwHh0RQ/b7kCZfsnBQGvneH1JBeZOnNDIzgO6Iy2kGSr6wWXlmS
u5ZDeFFBqk8Bix/dbegARdYlH1F2ZOEwFSuM+Ou4wzqYLpLpBhx/IDi7mTSBRIIrdh9jMFfAYnkT
HFeceX1GBRKR7Po484G9hu9+jCcA2biLDOXwdErM8YJIJOywMzppptYjHskgdV3lKMJhhh1+7XcF
y/9QIo510TDIP4j5U/4V1QV1sTJdmnYMz8+XRajL8+Y4veZVoZZE/xrEzDEcoDwo4664J23Glg0L
R/xy/SHAk9vtx0+1ei0zkNbdGkZJoaI2grBIy+nXtJ1E2Q+bxcPoizHsdavcZPLPe8WVfYC8Buun
EGBgw8cY6xJp9AukIDu0Dt1KQRkJ3ocCVXo3JxbxTqXorSJKpo20AkUjLnpla9rDOuWpTUJPBnu5
RD1Kj/sYTbK47g+IBA+dDdgPObesLmbc0Pl2iQozlUmBt5Y/bN5HU03xFjzpm1Tjy6xloKjDWoAg
jtgvCa8MhkT+fpP2wPpxS8JyfgFt8kU9Fxqzq16x+cepf9Z9rHYSXI/xsKxsbAqugBtZdCVYlN7v
R18NN/pvJPBBdwa1mwM4U7vsb+Ad1ug69AdCKpOyXEkQ8+FyeOn02oWQN+Z9GPZKdlRMbAnlXnQC
eLqEzS9KSZq4UCRFH5yHdIcjvY6mE5XKwsOLv96pfKDedY41AYBDCHur0xStTH0laFTCkuW1dWAE
SfxwtPRFiYG0QOgyCkfETcaOJKD6JPEA63VD/k0JpTGflwfzT/ZoAfgSqaBDKZWjLISYq3ZoTdG/
j8uYwMXaIemRgcvYmE9FgiYtCxL6UCOAB2xj9Kcg1K38jQ2GYBK3TIuf1xWK9FtnaxhyNo5NnJUi
oeZ7kDiWJpwLUUE4cpNtt9hoO/uj9G14s0w9J5glKmb6tZz81oY5W/flY7eu1je9JbbUFQELKI7V
3TfH0BfHNEYKabPXArtV7Cpr8IoZj5VUJaRQTKPV/9/ADmmb0eWeyQ7nGPE4wf56if2piofS5jVf
aPvFK6qnkVS6SLkyUgTI+0h6DkltLxl3AeMpeQhrd7PnNcm9gYVWDq7tVmhbFzmcYPtZcYkPUG/y
N13pk746p7CUW7ZxWs7mwadH5Jje3+Ifv81gzcdfRJotVioseFUf+VwmwYoaui+uH1zRh9lhJI/l
jjiRA1GyiMhyG757ilTJDHroqlld+oOvER0bsFM5Ib3Z6gM549Uh3AGMCmCiIuSpJDBVTaOe3BK6
IJnD2UZBhFJXlwRngLZv5qfzyjwf23ILI70ibOxod4tFYLyxwWzs0rA1Fle7xqhv7mVUoBsN8lkT
tvZRrm8Yf4M79sFk/lWk9CddjNMcrcEOZ14n9tF9FVL4fc+h+a3OalAskVocVSUC45/r8W/upqLi
KxQ/+9cXxZWkhX8oMw7jKoqnsPGkEEDUqUQ0DVvAnKIuTyYoX9fiuWlM+EEexsTvrQvj2W0BvQGh
E19TGtsrGbsX+0oneHaXHVFfYMxvk0RtE+TfzvfRe11UrQ3llukzURhfKm5X116W3UWn0L2k6jtW
Qv0F3qQ/IEyv79TXXkappYRz8cAxk2QJMp82Vzmp3wPqg86Hr12n1gFJD5KJK9og3xagy3BjKglf
NanZtjXs2RqetEh2q13WAzSx6x/A0xhXYuaK+yAU1QH2Nd8i2Wc1MB2OvFA8o755ox+eyll2U9xp
gv0CsM3yCZ4jPx7QyMo3RE3CKLAG0P+lU1rAWaXLDikQmIJyRxxy3et2JEe/8BrC3EEwGoO8BLVY
v6wB2nDgwashF3Wx8S3FDB47VR1NTkIXkyvJ4Zey53QRpaa8jQhO7khNCi6KiGhapC0NfO5akmkS
65Qzfz/hmU4JHmHu2yypX4ReDca0XdgxJuwzNxagA7x8NVscLGUhJ29A0EpT+acbi7bvheIPWcH4
OGXKhdemrYAxdjdZnMFCYZ059rpIqeb2Qt5DfPSOKSSJYojxP/h/6pJqxz98rLmgTyk4XZCl8q2Y
z6D3mhbIC49tdFXm5iJ1wn7Ylp3yEsXwUt2VyojxvWLimFv1vSwqm2p7u1A7os1ugeAEuwpim8ZY
PWxRUO4obJ29Lgq7oGqQElHZGzgcCz3gdxNCY0kGkoYXPsp8UAWwcb446CNLLDz49o/3ZVkAzum3
14tDTyGBBmiMDNvQ5CrI0VYCgnVhhYomv9k+/4bwtSqL66nFZ4R44sVLHJsoY7cE7EN1m7Uw/oJB
j8+OFz+PhFM6jZk80JxSo1NV4HRXUv+lYgVLXrx6sci/QMGsqpStQd4HA1ymgU9QjAFq+r4NG9+s
W0VDu2iBK00zwv95m1LOpTOApKL0E3pI2+ecla1qftOVvFpZMu1gVEpPxCM8/RhciFQwsluCUEyy
sZ5T+gC5G07KIUs4MZSY8BbqTmuQLuSa+xCRtSlOfWmYDzlfSoOINa/Thx3mcn4gTn9Xi+kMih1d
GG44ZM2lLp7+tE9DneZWt/jRoSxstrRbQW1xdOOmE10GkVCX8UYSQV2x+l8EC21ZHdwBZnrEIwyL
MmiNU0gJNMDpNAMjjSCpVtspdDtVfoAeozB/aAoovSZe9mvwRAUsD/1IQjHXW2Vr6eB13Xzm1lrs
sdlIeHNSlzGjnsJ+Fh2jHocEBrcNbr3XWBSmWzxMVSIzgxkc7iYZ24CKwBawb0qtAcGspFEhTgUq
0TinBVMzynekM1PNJ4byyhhSyZEsA8VkFbGo4Edf8g0c6gXMviio/RrBDJHEKRBBVzft/d//EZGn
FEkhtEEg7DG37q9Xn/biU5KW07ghEANEnt76/4hJIE33N5453Cnvr9uk8yeF3MNJ3858Ga10WXtt
F67V1NF1NV/9eeypda3XNPtPcFlKZD5sRq8hDclrDdKuado4p/YqBVXsUM0gCmO1CDEWp1/t2dK5
wq+pGsmRjNHZKbpz7llJb0u+ygLqy5j4T9CcZouPYnnGD7++L5L3TkLYOf/SM9O2rGprck35OUL1
dF3Xh7EqbUUIKTVo27bWyjT7E1qx7RI//+Ku4DRtU7c+B9cs3LsPRq8dn+8c6cYTcSK7z4v3mh3F
ouTI9u1usoWo59iyT183bxKkgM2nYO69z6pYIKzaeyKnRiKBMl9NkR6O19Ujv+pkf7F8kVKkUYO5
7ALkQ/0SFc2JT7bGLQB7DyWm/jQTHhSAUC42vVOL63A+Av50R7iIamF5w5JYnPhnc9n8bri4a9+Y
+oVR9c61h+CzZqvXxTmrMXDUVcYGjVQ+EzhHYDPtxmyVJApaesyZNr37k3750hE8r4w+oNnL84Q/
2R3n5CWOK/evJWXTjBPQ+BfeIGofV7f/TBFl2F/NiqhpQJ/fWxijwkJguZQl0/6XoLDu09AYCeNX
dnEhjFEYs52KkA1hTlhDg/zDNBan1Wujyr68RbzgpcWoLmA9S1yviqljZKIu97s2MzM9+PZDN5Z3
mqETYnYqvCkxf1gtjD6BRdZgTV81Yn9Rvhb6kMyZUHfkHRJ5Vvkl4AsoC6KwWudV5TUEb9po6jt1
16QgHMlYoW8O661dack0G0cIH6g94rDE69TpndFkvrOldUDWzK2NokqlI2XJT3bGs+jFc8949PRw
EMqL5FxtL81+I9x+/FCFJpJDC+mCglK4Z2A5g1YwNK67772rcG5KB4T/WT8Lpe1Ik/QVDVsBgkm2
XDMX9sVrHxLCYHLsyBHStqZC/8/kCupCr1c3Tnmk0l02EI7OhceXNt4PfReKiPcdL7000CN8fUW5
3z9DbaYy+rkNs3tHPm0q5N89UzDr8KMYTW2UbLpvIG1WkfywH8sIEnS8PBmFWrmGbV4Xcq6ygCQs
PpS8Zwr9umhSVCuNRwmOQpZEQtS6vr73y0t4gJwuriqjBKEzIKhfyvW+aIv8cGURuCa+FOOtTM5t
T+Yo51Ie1lDQBb0tlzgixiaaEHOONTLlGGzOryBv6H1GiSykRL0VAjSrgasNKZtf2f3dD2u4Jb/y
7Z7Wj2azLLhavOoeh9CbMr2AM08bzEHYouV1crx6sxJSYAimXox6ZWQZvHsfQTy2jNjZ31k4bgOD
VQmLJ5ssdh3b/YbyavVlBLVMDPDL/GddEJQ7ZXgOKaTIK6NNfb4OtQrq4YvfqkQSbAZhq3qU4NcO
gB2qn04j1z6p+l1iyBmfuQxUYmCEScblpg/8izELHxYWAYFhwqalFX55H91djf6MtLvHeqtLkWHc
bYYGsQAd2yRwmhE4zxQTLxnlhOoM2nw1X5s6qpy5/Va99ka5fmf8EaafLUjaUT5smaiKr68p5B0N
UVFauCZnj7yIPWQBWCxDeSnS43Y1nuiXWUmG8QRKHAXXcd4yEdtyjiVb05VlNF9yznvdhqxm3c0C
jW9uAGXDaU9FzNwREETBWmdApoWuQJVLXYfb4rhS1u8S2ZIFML//ifFaVHc9Rm1opDoKqBvMnmBX
/abPOxT/u/GwKSLqWcG1heKmrQ6Uh63avHNeatySNWtlWnJjulfBtTx8VA4gM0sl+cMSfLQS8Smi
eVltzxUY6XjClaIuct8GwycPk2d6Hc77EfuTAy+YQESR/ALeOxzMgfnYg8XlMXUfg5zJWb/tqT2v
c2iDNTBCxKLbrz3ru56F4D1SyljYzMiliXl1I9qwyOWGb7Mc6F9yvhUxnmUZL+YBc6pOyNd3gxw3
TzWt09Yup8IsXL4/J5h5CtAeG6J9FIp2eUsQFxx6INAflxYpLMnrhq1x8olAREPVE+q6HXraW/gf
ann8PXPaW6ehkF4DMC4jOHMIksoh5bMFZDophTpvAxcYx6vloDphgNTWrIzPQItQFIlSkzXr9e3z
UZT6TED3hcKmvjmQHBFxwsFSabiA5CtygnDulQsFybHjY3tYSVP+P+hiKv20LPDjlSFIco3tMoC1
7+lXhv7nMevVMBtbUYA5DoinlLGivNH+hUPsT0lUqUuVw1JzzMMBTKa6Oecu6xufYXT2760+K6ja
P76oao6oyIsu+U7DTFtwgwvEtP2UuJNDOW0IBCwAf/cv4JllJumIQXMWTr65HDdYmekyWtfJ2cGA
KhJHuuw8g+OUa4wl+EniiHNPOS/OTsxOkCwiPduifljDP/bkv29X6XUtTVXLEtEhjbjLbziNIicS
tWKHzOzJnUZBjTdg7+WWQpe1Kl+Eqh1x90cbXqzAr/GFMwEW2yJ4zU0vvbOQKEALkyAwg6pnegoA
3TZU4jpgICTZRFjvsLD//pFXmpuUWDouByTUcksUzQGt1JslR4kddPLOAS1+nSRccUn9QXvfLn+P
eCM4kI/7kzf4DAReOb7Yp5Qt2lFHP5kYaqTe5Sml9gzzZ/G8w6XZyzUHcDMCBEHUSjMDL7jxmWCb
6tXtmaeBnL9GhhspN1Xfm9BlI416++XtUbhF+VpIgfOa8BVBirjF0EtWoOkwPAyQtPIgTEiVV+t3
Jl0GRpeSphxy+4pHak5FL+ploB4RZ3dwM1IqkuZgVyQIblbQUa77JgQoO2om6zh31XK9ro9kTDJu
QWshV20S7EsqWdYSuQjbmhZlYg5dYn1NNGZvWY6zLcXoMzrVqTf49H1nKYR8TuJ78vrkmIycFbwp
TQIf9M0Sy6DzU6AXqM8b4EbWiprjnNvblEqboWXoXHIT9RTKObjWd5ZET9cr6nKiLvqcTX6boNn/
mbZPpCe/f5tj46/Ro8fODuF0l8cmYn+djOpFovpA4gPb7pgK/Mb+PJKY3nwntY+iFWEiBKPKR41E
/NFa/plqIYa3WnFA4ZFN4fuRFRclpiZ0rIo/l9q9mo2NZRX5Op5Ik3JyaLk0aGJdSoFYOj/gWc0M
uYYrFBbtvFX1+y8r7pR+Z//Ggr0gbxKbwhZGP2VwQ5HYcz5IzPbkYOT20Db9X7Cn01YovBDTEjEI
nF9jzgTrZoNhJvEvKSv1eP+4bdM75yFVu8A5HCSJZtmtRY3V8IiJWBOA6Ob41hdEDgo4pxumVLXV
mzeDl9URyqQYFwYCYyWMi30DzK8yk5dlmGwdWyTjiB/zT5BtU8N9p1jzLSMkMw6vsrw/4c1Jxq8P
1d2IVAXXSN8ZjO0PIH8GCobPLyUrM1f5cmF+7zrIoTG53HrWvKS25dxvJtb5BV3lut8VJY3HXPFA
khn+Rh54yUbdpw+h/Hd50w21XTjEdLFkFvvv5GbAwpSuWEWzlFP3QzbJVXkn6gclmrjnNUE9AoJU
cBpIDxlF1kCQVczc9/qs8kZPscjLX1KKOi9QyhNzPQcMx/TslHXSFQEJVk4J6SIC/BzMoZkHj0G1
hnqaXqXLM/oXR7z87ZZUKnSe91Vkxqg2qYHsGOgJ45J5rrlliWRcZI7vDz3yXIuRaFrahATe3k0O
8NGamLQn271kk0QA+7+ne2Jy30mZDGnqj0xjwicut7cTB0crMfqF/YKvTg/+eLvEExCAn8cI7s2r
XARjKhaeJU7ot5FbYDzD3N+12IQVnX9yOcrMzOa8teQdgHM0Jur62ivTrisUmEP8jEVENYt8sq7Q
iBMFx8Oih/5lqH84U+T3XH83KytRPP/5nRcZELefFJEvh83e0pwLiUlXJUlyZeCb6nU+x8Mrgcfd
rulnBYaBL5XgqOhmQeAtSYAHXzzAvjQRZprogViSEKRVa76dUuk0x/peF2DybvIE9ZIt+Hbq/1Q8
261UL4a4W5288c7mFgcgvSVuqdBPIMt+iuodm1feiAgDYjCoQkc8iTB5pYMxHqlJDAAUtNfSIxW+
j2pcVvwKiM7NeiRe1cT5x/qbaHlEwKHGNuem+BW+lKg3jC69SASijDh0gN00ewM0Yuipar/nARdE
elhcRR57KljsbzWGlPUBfuO66d/3Lb9WcGMvisdXK1Y9LLR70AfwHd9Gav6TNVqO8ThfLXPJ6XnL
KPZytCqFs3IkQhjOfArr8eh8D3S6I4OsHS8nmpnDAcCquVZP3zvHY8I2rX0XRHFAvIGvmNPKoXAD
UC8moufvUXIzZsTdOPDVaRCE2YPfaxn+MvJfuVIloHXntFiNGa4vt6YHZkJgUje6I/uqY3Idp11/
sp/kkLDo5PnPSFaruP1d/NuCKxE0JR5Q4W+FfwX6N1OevOjEeWJV2o5HnM42NSu2pSctkAJ7KT2g
EeZ5AlUWpYFSYSGDUKc/B9E6ajE0jTNj5v/CpQvFprSOXtrEkJr371d3hu99/P9IUjpbsaNSydDl
hl/oLpVx08YMTMxocQ4d5+R6s4fJoTdekpRzwZmh0Ee7sGgDwR5unnALhrRMDKYgAcRGniEltrAl
+UF+zoTL4fcEoQ/MGDkAQG2qsU8SFgc1mUjKGQfnYflEMOhgogJCKj1SoQTzGUoHysVdFklS3TZ9
IwEb/geGEi0At3K+5dbVSA8IdEgJnc9BB2i4D+FP2ZStQz2Wz+Ku3UerdlJVzaDVtbiWiLSLnDCd
LjoC4LLUFkCTicxyAhuUFqvYSCVZIizPjsKaUBHfJQ9XudoS4b89eoi4jTIPD1kfN1i7c6PKOUNn
SF5Yn0P5N5qKad/ybZUroN34Z0WKNwwK8A4YHVSGPAOh7NVO8BngR4ZVOI5vtYRAvB3BSy4qFEom
ubND1cvAi6vcT+t1MvljjHJaKfynDsGLksZq8d9oVn852fXlynvUdXwQ0aRT8fIJkWA5ZPC7+Bij
2dm9ypDhWBKm8eu4GVF6y3EvTLOMsOB85dcCow6xN/wBPbB9GCi6iki3qKDF3OGNqKmSeunbKx4+
ag9SJKkvme3PeCUxkSCxJcte/niLpAwBTI8YHCA2zd5tGNq7Ccty5cICjdmPTe78joHsDFIlrQUp
7zXK/jiBdDED56WxwSUjbXbvR6JLVtHd6XfKv0s6J/ZR9fi+niuNMHADKxYDGjO9x+mJJ9M5Tdsm
dXMmuXnuaAeI7fwsnnrD3dTnGttzdL2UXooBhgeenrNL3tYGWya+m35yBEf9TVvO+9567iUlZv2W
EWXIFRDe84aeRi7m1MLw4jL8mEkoeNJp9BUvYiO69ktgYalrSsnHDqTg56F2B3ltE5f1VDZjl71C
WlR5G2P3J8pD4Ci3tNQgwqgoD0Y7Jj+Qn3qOAlBD6rfCCEDQcythtwk/mx4ZydUpRFGP+c4PSnmZ
ix7CVyi1iPmJMKBVeKBlEd7Q/T1mQRN0iHO7szDeYKIJdnzl6QXHy0QxtYYC/+xGFYkDl9uxVS2O
HeIMsSktwRg2o8amx6eH5uzRnH7oiMxQ2h4aBmVManza1leMekhv6suaMDBlcQ8r+tSlvKMSasXj
gBjpsgF6MYmn0vnXr1YCloIkhk5dhg54Y3PK/lDa8pMeS8zsoQmFfpgo+UlSlqp/pzbh03NR/Rcn
C1WE/qtjODc4qnhBhvvcxa4MVxoa22A7RNNxNwef1IG7cMBnu4kKQGJjDvn6o9fg2dCa/fuuuhiV
8C1QjwQl2cMzmpxwuky7uN+M4S2b0itXSLRjKvVCUrNYLeL2xQF7V9nwmS6yG7aU9IP5eAwMSp6Y
qvdgq+MDtAXZjZCIEu6TW5ejDUgfhALvytmOg0JtEoJ/lBUtO7tWgnZ0v4E6FZ4hVMGGJ8HeIs/7
9AfUxqfnyFeFZwyhYRbq3kKK/ZnLVjxTFEIL7LmB33LvNr5Ld5arX1t920nkwCKPhQo10hskoWLX
XbJ6YvD7byead/RN3zdw4JV1k1iphRLG8zT/z5+tun4VnhlQhMqDYbghYQIxbLAsj8Fd2CvHKmhs
a9Eix19EOQcBokxhKUV4yNzdZPZ6EC91Do2I/bFKBu5bb6P+8N0bKPTQqHlc2U8Y0zdh8sl5rElI
aMzWfd/6kbMfi9zoDZsim5xhOVR7jpnauS7rBpq+Lof8T20TglGwaQEJ2FbgI4GCpa08LdREZQat
c+bPuyyMFIze1hDyGQK730QLkIA1v8wqJ1qU60QUw0hoGOtc5eLqIkMQlcPHdqaMfFUMOYzPk2aQ
gBRDuITxo3irIqOKq1mMQDQO6q/N/bblFehbYMsnbIEyhZLJqB+AaK2yieH9uGoXP6KIJ2pq/gPt
CSgGKjxy4HkrqKrOf38HmA2mk1yfwELx/i4f2xBkf9RAHIZS2LOHlQsZWs15oQn/4t4RQm7SRnF8
JDy8cOmMGOFo9DjcxQj5e7FDS3fyap5SY/aOwgX+zYIBY3f0hKJ+g8X64ZfVsCFLHXT972z1xP4F
zKh0K1RToBzXAYOpOXXZJU/CKO9fNZhdVJIPayZ0KO/bjJ7mP3M8buIh9TdBRhSeXwZ3unsT1gFw
eEL3dypCznj6INsECyXr1yZ3BcXF0pxwvCm5pBjz20C0v0CdfkSl/RHpkYHVbhrYq8hEbciDP0ux
zDEbXfznEcH1xoBHzHkYU8ZQap/fPbJ1YM7s75FZmL2a3Dq6N3GTpjE2njSYPZc8+iZXMfrYiN0C
B23i6ZQFecOanF5kutZ4UrGUcC7clu3wUbgFNw3cHtmpy3Tz9n9FesHtuyDMk4rZ2bRdrK1xRW08
pfjMHu0VsaCeUnY8LbdZY7c/30Pimd4dEs3YdbfNTBPdz6MrCqJiQrIN64NfC1R4H2JWkCQOpcmY
0IsvpvOaFSIw0koC0+WHPd1eS92th3pIsReXxaGmMazJuGR1lPOQXzH7flSe8w+29bTQ3HXPzbVJ
CoidJFqU4WPAFf7AscXB38WnGodGqx7Id6HKvs+AwMcvEz8LzajvpgsQKZ4OqOkLsrpDApdhx6Ew
y9y+d1nKwInJ7HOuGqOn+WKm33t5e+4DtXZD1JRfZnh6NjVDtFoEx9VyAL4qWgWSYCAFO7RKWIXB
Y+z5pa07EgqD1PrJJx6k4qoXnlZAqHs6FR6nw2bXMYTsYcNibxM4RHfBYk0yHe6O9YHGU4sfQICo
NO7siza844XzBvC21dzkKPcxRXqTQpVjN2HWHOkva4KOiGFj4xhtn8dyqRWcJm2gbaJ50nfIJ6cF
F+5pmE8B7d1s+1RC06OGV7B41ZitYp3+nDIkyk791qeCeK38THMb8uknPJrKuzM3kOGz9/3roVKJ
yIhdJstAY9GrwCvhm1m5A9J5DRnuj4RqnX2tneTXdL1qTevfYa27yx4J+tnum43bFZj1+0M9C9Ad
bEjleHjTGVlV2i6hCT1qh0/c3ylfCuT1kVMaZHZU/rnqDbVg/wH7+xbrXoVxKU2Z3YLHxwdx9nT+
JcnOyhsnxd3tq62Jjv8D6u7qt2ZOWvmpT5YHuZDRA40SSpodMj27m3BDKlSVuJkugKf1s6t+H+AS
DtzNj4/R1s/i1g8FoNabHwfslJjR+abtSjPqA/LzrmB843k8pPyVtegiZRuTaL2BMAluyTUiqCvo
C/usNeCqiMYccGnmOxZ8AHeEePyHSlOoqtuS+VkopdnJ+QqBL8xOZYf7gY0zJO9U/0zNZFiX5LAP
Wq0K0RVa8c+MznuSVp8zN57eD6nq8SCaJk72bUL160aQB8tf8f6vH5VQGa4tbXLJz3gkRJCsYSKz
ttHhjoPEA3dc5HOhAOuenM3UQzwd1RNyzxBaFiaO3s65va0yXc2CGl19Mh2TtSu4fKGoPtqaJmKo
vOxHCHBuKZsC0iboawicXVfjeLrcxvI87wCwGlyAxIFAsCxDg+ikSv+3tKOZtXYa+aW2zYrUSU3V
US7ZK797HLY05u1ZAol86wtxuDyLFl4ajHgnNg2WA17cJTJ7HST+QEMyUnSnnrZQPdABT4zKnl1V
eto++8Tzy9BaiMWClfF6jbFhuyZcjPW7qG9VjUO/VziAI00KinUZq1NCj8Q9ug1kjt9NUcD8b+yr
2Gq9OK1ctcOaK9ZT2sxCrfTdsRYLDzc8ZULUggm+pY1iDId/xBnV7Je8puT4TxOIyboIknUtAjNn
5+GUh1lSvuj/0Mgb5KqXleKZNDzUl+Q52Vzdv0gBN1VzRv3GvErkE0fwkFexHXL7zRM0Se7YCagI
oXjJhhCCqtl/65UJHh68iWCpaXYU0lo7lw+9iwVYZdK9ijNXmq65fQNqzEtkQhO55QqGH5WIUdNb
QasSMetDLNuK/v8p4VRvpSnoyJQZZyQR5xw8qrutOGkMg8Tcg6+6xY7shIb6sQbfbzxez0Rykza7
qxRfCJbLR0mMARd050AAtjGuuIw2p0NW5qaQU1B6ow7teHTVnQXrjo+BXpSn/UlQZ3o0nfiy+Wxn
KYmgKS9/IIBu7z22kEOGV9JBTYQCzQ1YiNCPrA0xN+tORE9piJdJXsIuDU4mYMGDCxPTlwAD8NBX
ANIXS1VGrg6Xwtyt9bMPg0ix/Dwg1gn0ioNNQW87iwO2V+WcUifY5qdQNDbUaupHyHZvvQlOSvQU
doButWZs0VpSkwvPI1R0ncmK6LyZQL/diW1aKw94JIXz7V9h2XzCfgtvWFOP5uXt3ms0/aEvblV9
lxclK8/j+SGfvkGclFaEWIOMbiP7ZRSUfbDCrcVytavBCquruJvBBShCelMVfLHC4+i6KS5WnaQj
9HF+S5mXNmnI7nhbKjym6egu3qErq8LhDRctU9L9panzViwFJx78kLE7kfErdd15gtm4o7OT6lJy
XnjcbFnD8brNg+T8PrZW1RCXDtzSmlhkYWjZ6zBHBsut8IXRwKH6hPQclwxZzou1L8f4c7uPbUAQ
j6BrfWT9nVZ0nn//LzfWyf51z8YDiYTjUF4UHdxlKoVbea/NXleBfgrBR91Dd5KNLLDBJSjxv3BK
+g0avGYhdZ664Eqj0n2KWNr09/dmu8jOrFFa0E+ouqpuwCeT2l1ZHGDI9GqG2dBMgs9XNMlLOOc4
E5KZ8oXF4mZhFBVeeFdj+kUDTdPjSOqiRIlUtj32YpjgNvOijKEWHa51aELSz76ypqcj7kzbn0Nc
imTISkFifbh/8g1tKXuMRZwiCQ33OAhqa19LwTWYgP8wk9wE/ukF99VeOP1APpoaltLQgmH4bjpC
5vc9vBse3fAV+bxcNjNNNrx/teezJ1f0qoFUc0zFv2zMIiHuNpt3Y/+YdogCzanQM4m/57OJoMCC
naV0AHSxRFFebLJoL7KeMwh1/Ga/PkmrrQQJ/91KM2wesPU0eTaUBIKL1NlBV+CYhUeMHkiQNXbB
kf5DwpM7O6+Na5KJqaEC9wSfzXHjnu1zIWrwe80ZMOPzsDMiklV7tbEzWf0M7RbElAES6a+ZflXr
NyCYEqT2m6FB4Bv6rlHQggHOjbEMnglgVrxAcDwS6qX0lf/VwMtlLgfxKaQR39PzdH8zYaaWNFmN
S1CcNDg59Es+QBUQC0BRNxI9VijadgLsWSZEzQKc+mLi4TWzI4/EiggipTAd3oX/vrJrTc469cPB
MthpRpOI5M7/7Aw4jNZ1Nl+eO7Z8EnFC2CIUzNOlSR+8VIriOHOprMLBh8CD9eIkUmCHxCrFFQD3
B0JFMMtuGZVmYMuuaJAl0Lzt9D7LGflPYmvHxKm23Ql9/c+0Kt+6kRGoMzIgsnimruOzHfU+rpYy
e2va2Yx+w3IIS1rGLlsM6vCGu6v4vkKoxZ6tVNLtgVUG6XyoeYbPncVpLpkuLjFlRgXKTABpCIK9
ik+OOyboB0D6GbLofoY+PqovWTyO1eeOqOzf9AStGj0I3ubKjimxhw5JsSyffPUF4+rClc0leOrv
giqqKDEIb0Rx1/xk8njrw07x8EOtC9IrnHHGA46GbrRAuOetOLArtArhzcXZvzYRgj9ZTZ/TLH5F
iSg5qEbPFjjdYxloMa7eQmkqsVloNYIWxJJAX94zvio8gmK8i84/ObueeGtvmVv6FSJyC5QBxqqH
PXHOfPNtl+NfHiM4Xj2e8lGo8mblrWoU/xncL8uYgIckgzuLqQGhEbIf6978FgDaH9GbvGBF2NKF
lNLrSMC2nxBa/e/PNSZQeKS0a9zhQ2C6MdShoHbSVwnhQFyWGl5Zvi2PfAABPv606t4QQwLZO/xZ
ChCzvTmvxe4zi5L7WUsf9aZzXul6Y+zYozvlmg5TPZV6RqSH/ap61m8w7IR2EH3uXh/GqEieNZNS
OB3NgzsC2IYey5xhtUISBb0qW3CtBZEo1ULN9q1ImOW5v1fmq2APdzM+Hx4e4zjPetAja2gM+UGb
UKAsAhw0qBPVgS6iLYfvHAU7nksYBc1uUh80ZKSlX6kuVvZXOVLZrL0rFXvrea9zhtcwy+IHexy3
+gtiBGc9/xwiu4IAFg8oINxobWfk4B58c4+2PQR6UGazPI8AdYpRCTlcift2U5pPcJtm0TQ6HPXs
8/kTDnmdTorFvzhLG7mTrscBYZXRsBaD74BcOdpu5UX2aLESUGP1oKd4jij7hPLrNhZj5oi+yhY1
r4rB3ac8/5bWyAp9Bj98+Qh2vxbmgZhlMT4O3ZqpzR1OVrlAmZMf/t2g1uobR1kDxJjIYDgzo4FB
ZX6Q/gJgtc7G0BfWVaqRtIaqhXLKMkUc6HU2DrZO3ZYpJ1jWa0LC6Uu9hhr88RYzD/e84D1WHVPI
OFwPVLoqKXT3xHRVTrXYj5GiLjPc+9ZJFv+B0ushRDTXRXQwpYVZKz2igo4ByDuoVLm03LsiFyOd
NaMcLaZMm9s+9goOStUrxEG1WN9Elezy3rf1DkkEeDeJpUJDXCsue8jkEoLTaKX06IVqVlf6ju2S
MIWe59FyfDVkMRMgrn3QT5NjbLNp6mpAZFwnK5ZcRm+NOnTTlGlWionmw909k3bSpMBGtHd4jsw2
Fxaq1Hax1bnY5W+bbMiZsqxluZfPfnHAx9i2jOmLMq4HV5dMDWLKq3nTZJTSx4gGJo2WwNKm1nE7
fYOgyC6+1NHHvki9Lq135VuSi0CTwsUYS/0BtSFtSEK3bPUG+L1IrtF96++QRX2l0FrqIse+7Tqi
Z4Cdl8kchRr39K0+UTO94q8nmeSUFYWLkfT2yn4iOHjbN7rw17fDd7l1FxAXDC/Euyo0WJynU4yK
E42EkSkTWN8KvyKM6eWkQO6Ry96RVBX4uo3FwLlmMqflrnrrZF6jkkus9BzmVXmJL9gFJ6uBgOb+
3jwQm2Zv95QzKgvs4vgWl6wzD+d0JTweAf3KAh1kx/Uc/AJUdjk83MwtMHX2TjUZIbFfBhaatCVI
GfYVWBAj8XwP/p0CNdycG4Uyq9D+BLhsAb+m+hjYk3AOsv5sGKvjo3hixC69zYdq0e5SoX/pmOtR
ltlUAiQX30UzHSZ344PZ6nRLo1o8UhbwHRC6uD2CwQB3/x1HeA7N6bx0tAQ2OCPbGvf8cHSB1IkI
HhhFP/QBq7bITyIir7iXeJaaqE3Th+7ncretSnMqZmGfZVnVnjNm708+s93857wf5sV6th0pjQVY
aXN/XEcIvfXZOIoErCWE+dus3UWVmSIoByH+VCo8DMm568bEywnYhDL2VdDZuWyoDoMUykWCnmmI
2FinR+rHg2JFxW5r2b34RWzwgR1HkBWQ0yn5jma1J4lxV4hIHPLGGI5wSQ4iwxKBqKRWzImNoWC6
G0Cmvx84QeLIpgKgmEeBr3+Gr7GSLE47dQiyRo8/2kSybXXQNlZb1VVHJC79/4aRTVVWqxsj76Pd
zVkiXBooXslwftlMHObGpHDMULxvNbIp3cZ4BXjgXyurV6CUWIt763k8HageHHWmVhWn493+cREZ
ALzXI8G2X0L+WI+1DeKo+MAd/3LBIslBMAQjmlvu5V5TZ3wk83KITbuJHq7IChqFfDNR6xiwuzxY
J2LT78RwcZZj/VftOak+JfcWyK62jDe3mWL1GhOCf+m6z5QPwE+ER2Be3ri8g1PfiMGMebH49Hsj
tn1KqXwjmX8/G67V/CBZ6hssngejPb+Q+eMqHMuSTBtD2FwLi/N53I+Pq+od9xIpddxPEQsQvSnb
ZBitbTV7CUXsFy8mS++n10X8ZZ6YsCgMgEgoueG0WhXxQqwULQblqgJ7gUuNnlKzwLu0HtDDFGsJ
0d/P1fw2jSc9dpYfeSdGhDwLeD1RFBFwuZL1lw04zFYlnVn6H1HxImva/gTtkQteYGOFv/6Va+GG
2zbY+BR8D5xDqg7AAFhgqq5aoZsAsnH47F6iLXNJy64Ume81mqIKwjBh9n1s5E5+AgQmGAPbNy/F
iAJR43fx7omKkhYx4U/0G/eSqORHbCUvu/xat/NVv597xX31Tt9FEIqczZtIq6/Oue7ZgzFr6kHn
vhrnfJABpqExXoAGlV7FlbJjrxoW5Ae9bpZDKqJO3r3L5X5QOcyKL8KCJFttU/R8/dTxLhKZ5ou0
6MfXimMch2mO+DAFxxaQydFKJ30qmh4ryYWFk6tqOeEk1igZC38f04nHFuix8CjvFPnr6NyjKirt
rTyTeZ1swRxDFsmRX2R8RsfVQjzqSnBtJ567RrFWygpIojW42B2icj2IpCnbvBsTJsJZ3zWrbdl+
ZKzhpg8+fN03hQyZwyeik0/WFj+e6qpKblfRewX6eLIp0PvWAYcXBQjqj4rkBzobgvCGMQI2VyP8
KNdJw6ff0izKWOvajK/szUBc35BZRS3YlZOYXU75PyudfB+VWcw0kcLRM1KrI2viDzl6PM+8I+E6
3EotikZf98mo0mEkm+YKfpcY+PwZsOLV2+893nVnlT9uPeAZKUNZAK22qSidd2OPfFr0Sm99fpSy
Hlynqx45I2cc1wgknPVsj/EeBTJ9uCQaTDZ9EED82gN2FQHVmA5+ng7v36zm9z2WGyygsx6h3jNP
76RvaZwAY9FwkjW+2LOTH8U8g2lkI7x1SGfbdVy887ARR3hoJuVPsFlSYpiCZ9lvVG/2ktFhbXCQ
4gEp0aCeaOxrBOXJZZSvafR59KEUrMCXX/XuZGlRP7cKrquzb6mtkD3tIVG6W/SH7rKlxj20zQRv
v0tp/W5whLEcsQGeT1TacqX9b0q5vg25RbN4btpgSNSu+eRmpCWBQ0UCGzLJREcMD0IXTAV/OXiP
Rc8xaOMiUU+PZ6PjI/d1OtLvWnQjztqbq3n3mA2xrTbMUtlWAYZMM+15JhsuUZkUemMvblX5Xdcw
twfqU8oVO2jP3jE18n9bKGjUoAY9pFUOa4UKwab74Dxab4yEA5FAFYEmehkDHyFu6Hi8rCY/UPD4
ViFlVnVIHSY289cDq5UAICbxD5HN5wBDCsR8YgChDPxZyP6cWnoyjGbExLE1WgMzt5SSdOA5Rj5q
voRVMSRksFYjGxPzC7aI9DbV7TPBlVQZxyiF16OHZhBkzCpu6rno3W/DYsCsP9SpTkjjpSB9zSyk
JTGfcHxrmMsiSJwp2o5uRlBYX/d+AArzIMy9ur336mCLDGNYDsPyp1/j55sDOWfAJaLkFErW5WaK
knCyr9pkl0pfhABZoNLnV4rE7mHiGDTtublGHtkMEf6+kEyKRyAXzuRYK4e8qqopa/w2W4qJE4kG
o2UVULz255w/S5nfKyq75WeH7iQxuewzn6RrvE+FNOF7jODuya6R4rZQk2E4V+cfkEvG/UP2Kp0U
eQk1Mc8ZY8ca05p0nMZvSEE/iGmpJo8PV8Coo1Qhyt6UqRQHKQJ6HT19vZLVUUwDEE++Ye9u9Pne
NP/Ydp3rEBeMO0Y7GajlAYdxcfCKLKNZ7MDUNY3N7d2jMGfF7RL18GMmmjoJGcAnFRCEajNkZWus
ebKpxuxYEv9gOVkBVcgEzRns9mrwpIl13o/NfXjdvit5/F4zOpU+JWmjquLXzCQf6vly/mwBT+Rg
PdC6bbkZyCCKJnLtUz9s03jpYqhaLYuszSdRB1AeYICPdip3LpOXZQ98JrdY2Wwi7jTzsYivESn6
RTnDm1Yr3IHd1ahfr7rnko6BLEebtbW0mCnbeiaCZy991xrQ6Rkj5CZaNtoJS0hvL2NRwFTQu4wL
kn5sNprjtJULXOdMm2yuwWxTXTQH10Zpr/aRuXvOF5opuPFyOLDzeJfSHMa6r+gGKlXCsI0bbv4y
O69VgwUAj7eaiu5HeZaDKZ5voVGtcR8zWtEiWeCJ0aKGcMSR2Jy+I/XMSef7XjcN6iFbmQysOOL2
FYMzbP51iA9eS6YEY3qVEzzK5ix7C1lvXl7sK6IEZukDG4CqCbwnuJRgKtZ7Ok0jxPVZ9kSAcRMO
7BJH4yKAwDttsWFLqHtb94sQn4FxRbQamUal08uCFwwFbLupxhTw3YpTTW/tc90/cYT1XBAC+qf2
1Fz4wzRaXfSMsReQmvz0/x2CfxCM5IIkPxprypmO8Ym9WpnQmX2F1MchodiwD/wGJeZbWbplT+Lo
4HxsH3rGt4TnLEGncoaLBJDDUPxiw7/K5TC9KLtdEkuZv11hwO0R6DKgpQER31hFNkjQk85MJ3kw
lofVCG7wZjjYEYS3ptflVOtKt8+VGeHwfB39Aa57uGMlDDJH6io1QiBQ5N856vVZ04apTaBT91wL
6incD17/4kp4a/hYPsMJT+FMEmAln00ZsO+e0o7gXyQMzKAKhN5w6AM4YG1JG8xPlBpOFsrbehXN
E/0dPzhA1Di36rJsygkObpguI0dGJa6uRqa+xXfQL3ghjCZ2YjeUjMq1peS5mtUREiZVAFPgP9/j
Ep0CA6yklkKYIdh4+RIV4bmsoEJZHCecMAGUYb5TPB36KV1T1xyLF9mKFTxsCF/zNW8RD3nj7gBQ
/0CnTIqMDZPLV096r5CqXiP15Q/SZy/5dI8xkBPuHlsK/oRvgJXa8mskpr9mRjlOo+wHTabBxCP4
REruSNXiGL8xWnm2Pu9z4gG22kFGzux0ziGvIVEvtGTqevPHyVRfAGoXHSXZYxufnV3jLZqEWup5
zFLKJUJ7jy9lUaYY5k8qOov2SK+HQU5TySvJvjuVnr384QAzw/P6j04DkccSmJQDDaTgbyTC1/yz
VHf3eBMQKgdyLe9I2xkbySOhTVuXHprNXk+oPcSm/oEMYSm5bWdXg5zn9jwEko26lhw7vu9luriA
bbaa9pXG4RH9eEXgMxVjeKFmXH6ZgPaeHtlSzbmmwtiljoa884gjg8j4xb1e1MPMJFl9sGZ5BI8+
Ni7Yfzmo6ujIgAsbzOQNyi51hEMKkGMnOVVI8ngm7IuGWQBcpiqB5v0j+2ihCcjDaT7eQ5soepox
ypra+7O4dhu/6jlU3lZ3ThrQNRjbQOd3Tpt2C0MbV6Wc41UsMirfugLY1dh40aBOC3dhZ9zcLpsY
nP1xXVNtT5fZr6mrUsGuHVE2RHtVBTFHpZxXRsxBCpKNM1m5UZ7EGf8cJLXmRNpAFpjmJiui3+G7
SjbpmPostOKi2no9djlYJvCS4VEyt8JkkzMtmldeUbrB8b5OgFHQVFT1Edy7q1LPTV8EwXlfgZAh
o5Dmi121gYCie9n97jvtnyZC7zQKhFOtDOUPBA9oS8k/ct0k50xwHW2dJDpn+rFOJE7ZM3NViZe7
M4jGR1PnIQA62PfBTCIFlfbiz2bQViybgzLMSveUPP/JWC2Cc24bavnjx5lWNpQyTXQrxdsjgtkA
d+z94NGU/7qgFftux72QtEG0V2ULY2eAjNtiFe8WXV9S8QZvi5AaUByKjc2QJFbf8obn/0keXBdh
cPHAAZEcE/g2IzJZuHQK3LTnq+VvUaTaz50EKyHFjedvi3ykPKRLORn37Sn3o1P3tpDOI0i3srWZ
pB0OyBqGd3EJAtoe38+3X/zA7Gr/iKiKW8LY5wvSWK1BggecptZLIUkgER5uxBB6/8tjH/Ll1Do5
aTwlvsd6ApluKpM3sx621lYrL65mgXF31t2MSUXg3XhSDgy0mmWdkCHNhAr0xXHUauUHVsX0dWRW
NX/JHpshUyatfAQzvky+12dVJ8a5t+YfGvGoZa1XzbvybGETMUFhFP3tHNRxWIXTUIyWt+QuM58B
vKoIpZFrY1IEXDwYVLQTIWa86Um8mcrCGfXQq/TtLqL/K6S6WPZX0kUeJBE4kB6rdcYpjPE9HGVN
/ZxWAdTKbsWRo1VbS1lBpQzUxT1klbPVA19jNbvw40uQU1n5dWj7Y2COTdYL89oTz31Wb1W6tTwc
odyr4lyic0aIfoBuY/4muxw/4MTLYavdd5p2ls1djSYEutXIwCybMCyBCKAbWJo3+JVPCh/xiaGJ
ohR9XFK1QlDz0DVjCaFRDuzw7ww2/70DO+nogLecYqcFLvnmYN3o7f5aSXsnSu3p9hCIda4f2jPS
di/u+1lVVl8nknu1stsMoQz49C/gUq/Hw7o0SXSe7LdOO4/Mw4gL/UUJpDz9VOFPstBbTTvRezzR
ckjtbK0+oD4zsLpNZ6CKamu861VZnxIp9VznvasTlSLJhTVkkWHtJQTRHAPrE/FDc03eH4dLPi+P
B4DNQLoCth+4cublk2Mr7MI3yaQZa2Kr65EghWsgce026cC6ymcxUTKk3ad8wSfmgDvve3aIjrSD
k+wOxxlgGTWV66xpBv231DkwKX3Dn6CbJ+MBgbd8ILKvbqxqGxWnzzUTnPXrjb1h7m+sZOK9fET1
ph+XsW1mZoJKAnCOVmSjK+Sk09ZYXwX39JjNhcZHKqkJTdzDAE4jemu2YTWbAM6It6TO8t6E/AEh
OiG6v+4c/6Sx99nixh0y+dznWFWDiLecAChuA/A7H/noVrSk5LCe+rkApOD4Gl4SU6bmWB9jHWdp
sRtxkvhVhbTVcx287HkbdtKHaQ74PVxQbvRy0QiD7CxHt/ROnZUbgrxevfhtjtyP3rDd3VysMJao
gPIMCl0bVDFlovneHkMy3k6Z2gv4F+V7MJwEE6SEsI+zO63pEQTALdCE5JvJ/405eRip2cnZSpZP
GqHVV2LBD8EXWd81m/aoqyexsTqnzZyj1MZga2ekhpe0PW30WHTIslhojh2d2JkhEOULqzSCBSfe
8wsv0QlWK27Rgx3qwca2zFLWAY66lGn8vtWkFARqTI+0wym1TvEcEjvSvKFtvPN/l3e3mdwj6jzu
zXtbukMWa3CA/OflkQQxvmxwX+IKlzkD2pgRrsWON6qwrOI8cyuwmfoTEpRHlCSH9a3NsbYWmJ/q
YCCAtAw+g/GVjT74rGrKTmSxu3mxCcAgnMWS53OTygWSs/Ym6dPR3XJH3qSxBvth9A/BfgwlT8g4
hDvXfHBpo45625yBfb1rNAp58U2lNtbhedg6WKw0+tG1AourikCUifEVOX3GO2TWnjo5JKOvlmkG
AZgjynPpUKGlowSpp5wkXWoN1KWeBVfJRGSnESQ8ZlC/BRLCcvA1TJVIIe7susPMQCdh8C9zgeF3
qbM+6xgCiT1UKFpCzKu1nDdf5eJS8o9juWYdtKvjwbO1LfEPStJdj+Ca4jnByDmdWcj3EcRVtt+p
vFIf76lr3gv3gF8aWz02bpLvANeI67/Y3ZRZlmRXgDtb95Q3ik2B/OSrxuH3cWW3nn6VqVYkY5Yr
0iWgvlJOZJac9IjARchx6xeMLGiDvJvstIhYjmLjt4OUjWyMT5K30JgM5nY0NMIxCXVpdaTlpOCK
uLF7DxphcQBG7XtSkMc3Kfz26TTf1ApBUjcMhD89FUB4TG1mDvWIYdggkteI3ZYxzLGRzQkLPXGB
BVGEw8Wv42BvFm16yBQYHj2g7qxp6X1AlT+JzqbwyOclczusRPnJBqm1zzFjQ3x5onnf+1iYFzhv
9imdWCHjiSuoRq72s+bnvXFv8136W5+1f3cVzPmIxX+CgwWqvkLB7RJc217U5ijU3GtHuOwj08w9
WFO2sBu5IjH7ipc1n0zDZYeelWYatm2DQfNtP4WIYYygSP+9pQwDOY8H/W6lNQpI15qqiC2qX9nH
VUhT9/E54dEHZZMfigJyzAZZ2gCOlZUMyu0bLNQlIw5sdmO6PDyIe5b1ybpkvXr5PX+dKzJbEmTW
fYyQ1vFcONHztVUek4XrTCCQovUUyg2jcIf72iTo4zklfxjwI5GHrtppDNtV7bhf4/GmRbkNGeOx
NcFU5RAbJ5axeFaDhQ5nn3H0ZuRT3bx4UTaAdeJ/DmM5kdHzQnHwxEQFm3h8Y8c9sVGV2DY8RE2i
zo2W3TBqELjvXiUcEiA5Towvdnu3ZPFup2XxBO21CH2KkrLScf+hW8OOGsKsrD9AaQphJuXR57xu
l+w2avxuyTbYRQ0ayCW9PXLokxNCz0uEjVDCLag8NLPXxs+XlZ+r+XM3Te+9KfZEDjiGrqQfwJwj
hOUyPC80MyzQjpbaa9LVjNkBEs+DoG+pxehtdCvuENgiHGRzxPjePM/ND4nV5RXNZ1yJNZXZBtPB
rvDcUONwC95Z/4SMfzxAQzLzHrAb+/o7wnJV5CEGj4uGa9dwYLcDpYSLalHde0L5Gr+Y/x/QXPjG
1G+Zo5uL69wvEL0weTF499SQgcITanpOFzTncpVkcJa5nyHuT916vr9fqtufS0wIK5mIqN7N4yby
NE/y1As7uPdZksBpQb9ZqDCE9Wp80JEoDQ2v0/L2e3NonXr9vphjmOteWPmp3swUzqnCfEcfDKs2
T/e1AC+NqQKhJaoaN1+uUl0asaJHGASdHWjtqWndReMEBl/1ZQrGk/2ygrHXABUmBQ3tF8Jv/N3p
0hk2+ps6Io0zbFX+dvfLvPQqjg7rnOFeXLplD+NM+KMuI+y1zwcClPkhsFeDFC0k6Fu+vvbzR61r
oUP0QfPmJHkL9sQ6OZVGIebL2A8CCpVR/KsYpMPIM/v11hc5gLSlltx5sX1/oo7+ZarMU9iI09p9
7wbFlfGW09Jpogb+tG14iVrt3iHE7cqHeWSZTegwg6yi2OBkcLQhqo1hbmr9GkoEoLml19s2xB1Y
yeKww0NoOUKVG55rahrwFknZATStxIEZVKrQ009wlBjkjuOWNHIFwLndHY4ALGKIwS/+cs85rH+i
vpz1PdoidjYK8I3Cb8gLBijeh4e+Qi9XYSWco6bqxL1UNyWNDyfAx99Iz7rMdP7KgWDRFTzb9Fdo
P+5wFUjBWuUzqOYo8k6rEgBpYvePkUc6MW/9cCYlMtJ3Ff+ew5Uxa0ZyvKB+RlsdxevLADJMw755
AiH5OIVbOW96Tm1HcgPf+AkqpDkewzTfNjYSOs4jl+mi76pUv4xY1PTqN8gUFoHqI9FCsI0nEyvn
OXXeBdZlSfDpVDfLP4FB1LcdIGSPAU2g7XkvW0kuI0UJCidCXaGt9cJp6IwJ/grzZcA6Of+VQfAb
HqWBMl5CJZ8x9LIq1EqTjhW2Enq2Eb5OhMcCk5Qjmi0eyKp5xZX1RTzEuQEi6wkJOIrItjEGtbK8
iHnWm0+ypBAjMNMtgf65SsqjxW0WVPrH00Gc1knSQLxVM+3WuHNYZUpgV+GXzKmJ1p5bGMqAl6Go
h/PHsoDFHgyOvjaY9+mB7eSmKUq4lzfiqA97x+PIAq9g0wwLr/hwmWJd1N/oaKmiTXsgcRMyt3HL
Kxf4bmpbyheS9NyaQsEniGMyv5BDj84c2frpt1z54+7OUw0IH8+HNWIyqcHS35M/x3YzTon2/Ro4
Ee2TyiTdwHCodzBWiMBBXHuwoygKs4q7HK3Wc44bUeZutRL7xUfBYZrnGJTcc9lfDIpYPrbRmqJD
HM+Hhxr67gP7j3hfe3jZrTQiRrKKCY/CQe+akzxYCmd68p2iBNUTQahN9vRQpwQ6PEUKGSIUXLet
1l0J/sPYODHKXFoHB7mEKcB1DSHYqcRbBFhGnEXKsqYD97n3jhBTa0t1UQqvi4D/wYPtae+EB8Hq
Rum36HGaJY3OYdh1fTjVdARp9m+lEcVl3IZ2qbsJUs5vdmVTtk8/ypIbEWkGpfC4CQ32K5NsAR3v
+BaT2yAQGhkQIkup++u3L1/ULM5Ea6vKpCfOU3yrdo8/O7j2nE5dgIKMpRSqRKMsL46ju4bqzjYK
Bz2Qu5bKFDM/bdeHhlKJN2C/EDdaBdEYHRy7xUOF/tlUC8Jg3fHs9nOoz7AM9SBUpqRsz6qA2QM9
OjjOrZp2XdqAF1ZpVYKOM7B/KXQhfr2Ngw9VD+gv5ZQg9GW7WC3uZZYY5GRqqqgBatgSYPPMnKox
IQaMbvFPw8Hhxil+oRSRCQvy3VqZsPJWvYUo6Zthv3dMStOkhw2NVvU1Ek8cPMiIiLuNAKyevjC4
3+p/r3gZ+ENKU8Z9NAkIxOG9j001jjdZOqxA33CR2wsaqMftcKw4XgCHICwjFc0oHDcvM7Gk/OBC
XaUinJUL/kyV8woUiqxoCNi5KxcAtwxCm4XLsGUw3yJItZJtEGliyNGaqb7XfwsSqA9lvHMGcfzR
+rUxkBs/P1EhgvcBIgovg9BLqWF55BKm22TMfgPKlBRZSkEwLJ8L0kx7nY/3sFUxPhxtiB1Es2nz
vDnaZormdzubILibvo3cH7ut34OvLRdPoSZqPh1qrVFuUlW54YnReV8V1ro84lP6opuG9S7lMFAS
U/S4OBafHYAGE9twrhFsOfXdd3Qg4vR0RgqiVihaXoG7TLwLvAg/4ektgdK2TfP6a3ZG9XaQeAWw
PVN2VEinWNtNu9TBJx7Owh42W0BAZQEQI5sbLvELCejQ3OXy2icAe1MIKVClheKFXvg8pzjUaqcS
Y9K/vGkWOL2HEe2a9POGmoNY0RCTliZyMbWobt8256eRHanVh32B+IXkjfpNCQJySePHAmMfPk9K
vJj9pPu1mNZa33Ew0lJACDxgRU+8zKaxDCewRkwTW2YCOlrZNxJhtAUYY/GyM2RS7gE1eACNUU5H
Kw8mCPpt8oRsng5fEezBuTw32YkWI3D7PrJU1XJNzf9K/Rj5yKL9lX99irDay/kOZZ13t/8f6xfG
fL554W/4tkhBxTdUFRP7qvErW4eHr8G0lREpqX0zaHL/jlGclkkFXrBwK8hXYfG85jAk/8rBYCIU
m2T7E4fqIkGxbckFlg6cJpvgyMt8UvESUBv/a5QRYUP2FHdihTRcN+VUuw0J0pwupR58kyITpfLX
VG+8ypk9MLCEw8Z5OetK7oSJ9pA6os+oX6IAyTcGi1x9237coAY0sD26ZzfgyacerToNYl0uyCQE
tjLyrOfDoNg2i357FuqQ1QCPU2r1yFwpbwxln6Mq/SgAUjqD3D7NXwLk8og5AyHVPdqUL1L8RV7+
GZgrNTUZNtAXBlDpO9iOm2LfhQkVwSdJ0EcgHwtaYEwbY5P/zww5SxOj+84kNuz4kiaxFqu7yStW
WS5yW1OC3vNkurMdxbYEsyEuJKszJ6gsXF43jBzEwC1sOFCbIyyJ/ZH7iNBO9OICgUHH2NsHVkQD
vNq8ISrpREzQkPa36hoqYo1lXn+6CxF9aKz0pybdhWiYfXTfcgcFHxeFI9bzFgSVwCiTSOwcIxEY
SfYZ1mdEEexjhkEY9rlrPnMr6zshweUEokXQakmDMbgHghyS+aT00CBlxIq47iCJNEPJ3uYGgiqP
R0AiwphZYtYCKi76GpU0ksojMpzidq4B7R3ikDaJjNmtHpko7WZZ/LRmO9qEUdT4UCXVO0kKV/1x
k79FRDO8vbpdhfphF4x7TTR5EIKtTAm7ThBGkCq/7XLWempG6LAHxQAyX6L3b5jVEjPMg8VkTs1h
JxWl6aGEVkbQ2JQ9XQyrlbeNHniN7Tkbo+sUEbrstdoAOFw1iGpW3mbHKW+Uqlg74SYLkjHvSyRp
wQXuEMbHJ1/1KMtz1WnLC4FYQk64+oku7WpJd2VS8M0TKL+ST7tH6M6gnCpP6cjAIQWkPU+5YcPP
kDTuZg89SURCAqMYvotwZZNxVZj2qr0e5qwi7CPrCLFRIykYHrRuMqn+WfMAQkMQX4+6vM7VcYjR
FBLwAlogR3Q4cUsdBUZPK8kATINp+AooApR6xcHG0GzMhWnI698NeXGojzO2Ce0ILzNrnXRURbgK
cLMoGG9lBsFL2TUIt7tRYzD9jXL7G2w5QMex0+KjizXWoTSIo4AR1E1XL7a1i0iz42vgxhZLD4kf
dPHiPFGXMrrDNMe2t70088+5Ih7BbW5eOmFEblulEj1yyKXE5xPKOWoRo83VCjQkkeXUN4QRCLXl
SBDNR07rap9U5t6m5dLsHYg0euILsL52d04BRyms1kYNXnbw0CHCGWs/uTiU6tI3B/n/gXro4wHy
aBMYcV2C9/JkkPwJayorAn2Lc35KQ/FN9UwGUIo++bZwSdRU+OhKHDPn2Eu/Fm/TBHW649X9Kv9s
kWfCNjCM0I4h6tsll1eYXjvx2a7Nh57ztViUbrbryJNP/v8gb5iebemjZeuaQQ12kJOeT4TKiLMk
AYQEsgFnGB54HahDw+tyB2rl0IOe99y7rweZ+u5kCZF+oCOom/KAOiDJ50WyhiDYDWU1XnYkre9/
KTvz+fyUfGcBoKMNDHOCJYLVxLZWt6nnEbvGMJ7hjXzQMeneeSvu0tXbA2UKIRRo8SLcBLJyp/a2
46+iIeIQDR4kda8YAvZYyaREr1Vg9OddRax20az0DkPHmkM8uIFlVoPWpuhxaUdp9mtHdcAqLfm5
Ve8iKkp2CmTBaC6XWKKdxnxE74ZkglY1PCQMSFMwHO7b6Ls401UsK1sk8aRct++ynMwZqhIG48px
p3oLqK6xI7wffw+cXuLfjMJnRsEVS9Tlutno6+QhHpvGRa4ac2DFsbTe8q0h3OHHt/qEPu6ecPkF
agsXhKPDI2hE0G6zLkgxsoYeKo7aOLzmGvkKCUlulvwSXVmQess1FuUqc97aKm2tLzsB07IBZRih
/AJ5VpI20mPy2oIq1SLbDeGs0VzoeO2tk+cX/8FdNw/UKokSO2X5dWke9Illd5uy4JitnwTCs1Ax
LH0XIQFKFD+TIDET6SiPtBVGYcQmJ3WLrWRV6e19TJU4JMN6zs1MaU061PhTkOqIZXheCm6Utnh8
ir4ptvjv+iXP6Fv54UlBSCzAeHgUrw7+d+FSUeSH+oBz5GgFkZEyTJjNYjPSxaraKvb9m1WX/PJl
X+/VjnfIwpYl4uoMZJ/syjpy7S3Qws5VC3h5rSOWMQoX0Vxkaw3HT12N0U1VUyImfft0AUAYqaON
b5XoMvIlYBjd5OzLY1F3VAm58nY+ADpH2y4OWKSxYVjSNH3TY2RIZctRaxy1yLVlEdi7WUKXHSdb
3QIIeuAbJ28nkDriIkO/iwqlWqBjd9HNZaRI4iA0B/17xrh2dRkZ7pfFAf4t715gaYqW4/poFeE8
QelkboPu6dS7fZshMEfvvXD8aSbtjYIxgamqlNYBR6NV1dfqTuCk+I5Wv02FPOcHI3K2sA5Yv3fZ
imxk6uupD1Bfd1OL18VkQtLtZwk4cUimPU4ho2l8NM2B1kT2ykP0TiMTBIszEFHUu835mDE250T7
nzmfVe4zWeO7SArqkzNus5hkMsJaCoJEMnMs855EV6Ul9avou+vBRHK08bVklNcjS30nQGFLVS0L
JZFyonJ1KC2VZxkcPdugT08s5dD1gxbyWyScVg/VLzDk5Nfq8od4wfD5yIFcqVsmpT6Nf/i7XJ4+
7Z9pTkD0GxX0RosHmoeLAX2B/rWMSYaJDTR66lQv5toIEJ3TyP0k3aOaQweIyGL0xjQDRoTmCxRc
3kAWUTD+ILksCae7KMJODjJEO/B8+x9E3+aJGEd1FP0eqsKzCNOyDmi0muFRyP5GHRYfmKVjGRy/
Ql8kC6l69rjOfuwhUH87wId5AnPH6SqY1yKAAsCQSZss54QXxWChf01GXES27XGMX6XFD3qLjqeW
N8sRUUqUS+qUfgf2wUGfRMriVlc90s2Avt1x/4R8Zg8/SK9zm1HrySFLx6feU9kKbQ0DPbnFyKSJ
Du4jt63bJ2qLPYfjpO4va5GppkozNYy8vPHGAagAZbe/5VA2t4pDTLmjET8ro8m8H6tTXfISPEaV
QuF9C4QgKNUgDP5gA667vQIeiveYCJ8zZl9ZnUVCCCwMLxymd/bQsf7xT6LYB0YSwKe5oaIJ9Zum
gnu95HQA2Mo0ANfraIiZ3LAWtMwA3TdrlBlgU7NcR9COpg0V4l72wVQ+PKMdvmuJ/8/DuwFcS5R7
1X2AoZxUlx7PjpkQ4RCnwRFat3uKLe+LShR5twpyi9lIB0TWcHPCGmyBc7wPROdBItPKapEZxZil
AyMgs079QG3RsfV3ptuL70iIfOh0iCSTQ1T6Cfhp9Y4Jp8mIv4EkMB8oJ0pZMGEeZvdDBcAOwi0O
AlrPhDFPPIRdYBoANnx4WQ2yjZhzg5QzIxrw+Wj6mL//Vm0anlY3h/Qyrd8E2cudANrMUD5c5Cru
IHbuyojEEvWMCAk7jis3Mgh85heCcEp4950z3JkugipULYF5jNl470eaxTWxo3pJufEUDQNQazyA
LRv0N61gJpr47PkSxlyiBL7gLezCQ5spD/Z5fZkl7fSA+8iR7iCNX07nX0wQvZpWYql57jNKS9er
okaXnYZAqHSCFYRfD5CNtIVl3Fb1O8ju3ICegWKQeTKAAXSBqwhd9+mRGT2anWzTtXLKRv06ClXU
vQeRNtQGpbpIN1Tfcl4zEyhwbb+aMP2INVDwxGIPGgi5ZxKckQl1qqdOzkc5R5XJZXXfprJMr6dA
IVB23eqoPWGcUDl7mfprqyxRgRdpLiQqygfNT8gRKmkImT7dvNXIUJLiddRj25Bpz0M6hZA9EHbM
ho3drzuAJSZvOLX59xQOOOiu7pC6dUhobeWhft886cYYAeEviC/4p40LIXBMt1h48k74S8t7DyOT
QuzVScmop5KnKWgpcRgdVp86jdBB8o2fSqN8gmsRPq3A+/vMOWB+7LgNldw9/CIjo7LE2y7H6F3o
DdR7Muifq71TwIavv8ute3zr/7Avvmr0hXHPnkSZrCXnPk8bXij7MEoRFNR4NpPXPXLRSrVyGrrf
2c0S21xZkXEbeEGYJZwLi3qpe5bpHY4T8nQ+mLvMTUaVS8xRmJPPVCGC8gP60+DmkKo+xlLIQz1f
vNGlRcDoDsItnHULQrvfsrXbuwNMgRAYgcA5HE6EMRfqasI4FMXdFzuDwhrRG/z5a3BqtzFO6mLR
b+WWyX95AaQHLnzjOmRkFMlcV5SBUmJhxnbGWL3VfLKLLn+gb22WH1mVwKFkJDSSSTsGxBLcHCQQ
z2/03dK18F2scQcye6z7WjIvzlXzT9LnT9xGN1vVZJZzQgbXhq7SnPb+pq3eLApFYTzzlzyT7kxU
tSH318aWbbs4VY3aDnfR2SfLuh/qLpQASq1s7qabafIiZvgbrDxa3o4ckM+bjJRuGuY3ofsFcOzq
kl6dEcx1WKHUtovpJsDUSQwl3gDvIq2LS0bP7QZszC0w1aGyaghH8RzcwHfKUa1LsI16AQqrqx5T
x2036aPSwHr4WT1fmt40FChZ+9/PHJeFrPqYNJrco5VZL/izzP53dqTwRgI53USYgAMy01/vK+v1
LKc+dorumjScf59nGYGpSH08Nxv9v2rxehh7fBS+GeV9M7wz7S9gbxKOYKMzldgUwdfoNnMNfWxT
alg1skvqVN4mDyrXCLtF3LlrzPuCYLDv3pMTFUpSi0YzWMmxYoTtxMEWOiYxmsTwpkc910IQMY5V
Pynbwjep3x1yB1dbW0aPoQJNDcNds7THox3j7OIGR6ffQjkUy97FWAo6sIf7TgD8U/5o4POWz9E3
FAXE0vZBOZJueO6oKI6wHkPlzi3094Z3mdGIhPVOsHJYz7g3HcQW1lMmKMlkLI/0gr/1/dXSqAvC
lHZ1RyQzsfd0BBj12mP6+/crY47lyWk6hAtAhboqixcDKZNovW/3McSfwz+iehj+C6MR0dTT7shw
WaP6JBhHlNMv/Ca20sV3jMpwq9xAXd0HSSY6WtXvJKnMtyPUz0HBYlAvO3htoCG//AsZHSUhFmcI
vN2770cU7PDnkaM77ja1+2JqYrFV1mwU6gSuqb7SwOOKkHunAbBg/ch/kGeheZbPkDPM2EIrBHNs
BclbgfpHHy3XWFaWJxkAXs0R4aeIvirKfHpRipwqjj9i0jHrCqU4CRCEWk/hm6Qk49xRqpeRc1w+
8kkAkER57LNSWkjGMAWSHk+2eDSVYJCDyI1j1KuWZFWRDmkdKkkYA6zPfZYq9AGpBAta/BTMPVSu
ycsQDPHcm4ZUnIhmbj2CLJJTi7w6LbYDq3xJaSSrR8/2nfKRw8d9Tp0Ql6uKWyW/5CiV4Tq/KMXr
6vuQSzZnOwnWm4kaJjjRrRgy9taAHZIYcR6lVSNXAt9ZQisNktM+xJBfU4WvRCkDjXmbGUyXVpUs
kNQc2DdApkSdx9SaDEJYJIbrrbx4vkNrf5ifk+RR7RIH7VTuDGkH9Gl5gZnxZhCIM6m1waKBRPss
QUNsp/Wlz0O/QB5nC0ooqhucwt7ADIuhP5bT//HpCNYOEQcXD7gJpItTkk7cf+z5jD9KKtX6k+AQ
h+MyySVTt/GOU/k+iJ+YfwCN+EO52tDlX0SBmd8Ii9Hu/G2hAFjwRLRB+b4bxMO/tHwlWbmDZhtj
+OmpVjza1w1x5dIKOdqME+VpaZNsg8x+VnTUnLYw26VoGeqeLh7t4gB6PZ5GrhvXVBIstxnFOE1e
/itvp1nCI5ZXwfnBAeYKkBXfyyVpTqbXwx15aHQ41JUMR0RRFUFXurkdS2vnz1suf5SaaKwIIdUP
e9qfES6hFx5+u364LM+xPgH7hqd03GJC7uDtgbMPcEdQ3d5HCfsCb+lDcla9dgcbNarHs6qxgh9u
ab1e7euhAiXVirzAyI/dhEoliFK0CBDH687TuASquWVp0YPqL1rAy30Ixd/H6fyt3iohPg+oqbfB
VlOLxQcn+u2YaPe1q2GXnQOMBGAV8vLIXt2WqeDAYLuV8ImlgMJkKoiB769Pju+tC7nMDDQtvE73
je9sbF29Vv1d4xJCXRRHEECeTkdZ4kPCcpAGokxW3w3OCLPs1lORE4r42q/UpGIfFijUjjj6JuhS
Pe9hXAzG2cl3yijuKuW62lcUMv20zbOLnG+C6jZQEwmLFYYiHlKDNaqRp5t9xqr0gxgOYhjmJZe1
SLc2A5o7if4fPjXBWHhuPoaJXMywBNuMnzn4GNBfJoRs4ejbRwUL1Ud3E66atNrFoxQSFx4mgS2P
QeELsaF7KS59H7raqmD3GXhC7zxEP55ImPAHr7hrGYUUcUGUOOyzqss6dl2CEoZtZMyVAnJtlgoT
5XTwoL4HmYT9Z6AuXkOuLFBV57juEu6XK680frW1M30Ku3wHpE182hxtUE000Nc6+BoX0o0ooSse
DSTGq0IpbmZp0w0BBXceh4+YDp/t4omEAHBN6MEuohMEnU3WpxhRQdPI3tN1TFa3mOs2c8WOihWR
G8i9TClBkjKiC49XpyWTYZz1CCUSHGu9AKB5rv3RYXoaXU8B/RRJxJCf8sdrMG/Mjen4wfK4Sw1K
tERN1jCq8jb+E/9nXxVJIj+CvuFtuYzF9c6Xr2dtHdX1vAo/Dtm5vMVwjkDdVP/N0lt12raVrAh5
RMgD6LwYOgGFMOCNuGQJsIy62e/g3p0mO3qObsn68J0eh2n6iPuBJNSRo3qptRV+DLx0udlYMWl7
qDNMtCV7mtJieiQSPw1rN/wmgY2OTsGIUj1bLvMEMFCvA4+39UhsWhnbFJCtHjKrEsplfXTh53RF
Q2kqBnBaoBzftCtJCBPhUiAWsvq1k/l5kSdtdW7ODbrKLXqte4EfT0J+kltDh0OuNrrbmMKW4xRT
eM6wHml+5Z9Taxail+uqOJkakdUvXhS/vBfCmaf2CpXIua9aev10L3/wuaFaWmpVAAV5x5g6QJqy
+FOoqZPS6v0l1D+POnLYnamVOFamjHbzVOAjhkOGCfOP8Eky3HWVjcpPgXosOrifV0woi3bkI0f1
X4JT5MRJFDYC1lSy/DVtmrN0F/Gpx5+9B17Zq5PU+JsKFo60trBAGkzrnp5vfvf00bq0zi0x/lnf
5ik2CMtcrLpku6JzeFtjjP3fSPod9oOnw2jYfa2K6c9FUIsC4ci6ccpOrF9JCxuhYU6fPfmhn4iX
GcqPo9XB8lLcHeILxzjxDpJQ0fqnyJUQmPBWbH5sBG8viTsTbakGZOBOKsBa9gq9nXe3m9hSjAWf
rXq9gsjceApxP4/nUNEpVW4AYJfT22XIqYhIopU/rwGf0OIY89llCSyMeQnADYlN3lyl3L4totwv
OoeOeChMcgWsLG1tGPlCOGNQsCxcUwDb+OaxvT5IvrOP8PtFErrqjciKT7W5BiuNbXV3qvS4Z5U7
g6OUP2IeLL0nu2chqwubXpDazru3DXm3bd2C3aMXzEU5IXXLWkWhiHH71OwDzSUXfBRhmLmId5zR
aMqG5zfy67GLGkMm0bLtGlU9YwxQ2v/q9WyUI2S0/pA2HYk6AoyPGZFeoS2yclDwf/jlePcmHnz0
rrl5jE4NOTcfC0Y/OZTunSWOg6/cu+w6szJk35C1+sy4HaRpOXBlN5rgLcGMiK3p+KerNbabqrK1
lhVfSmOVLmU5CCn29OPB5idCLUh1ORRE/XgYxhuql8UY7XpPMXn7SEQeok7qAECPhnzzFJT9tIaG
LeijmEVin5cx/5R5REK7VwQSHFjoBVi22rQGNSU2cGvtiI1b0bo1S2J2VOTc605FMsriOj8TsAZt
8BjU4SotfKc/Y5g/s1U1qUGgvQqSqv8C6KcUxCRg78KjZwnt/mUyroc7XucJOemGBAQ5BJOSao4z
S8litoU3HY/0L+0jjisFP4uwGfPzblivsYU+reCGKiTN2Q55esZh8G407A5QONwHX/FtfAQRVaT3
yemdZiF7PSbOSt+SWIzqzMK3Y71+LnzfI63gVWB9fKO2d0jKNZKOt36iLKgZ8WhHJQWuWCUBFWQC
VjcISKDcpf5I/ntY9Rx6vPewI2FN3MgJq3y0z//idhCqKBjgu8aefVCjP0kUZ9sCf4o+zHoRz7t9
/+lY+q5nloFPvC3EcTqRht8O9kPmdV4A2xEFmr9JYCzoDCuYr85RD9rf21q16R0moc1QGUP25JXc
TdmaPlZ/3UEh0SQI5J0YqSE8F6wy1K/THJZb1XUbhbOvcCTvNoBKCYr54vY3TJo2muSCGeI1Rp3o
2TvPQ4/MOXA8ihVcduC0iBWcXfGLokUg9gGxLPpWupphid1/imJnLwHx0n27O/JANwMTXFBEAhcU
NPQdwjHiLmVLfd4tiX+D/z2eAj1xrf7t1L/8ONdTGFjC809c7WnWPvlMcMfNFu6S/yf9bxVeR5HD
02xOzQyM7G80I8Aks5BElu2lpDSku3iMMgDlqXeW8Tp1Sz7u6YMRyWILkZJk3h2UDSt/9qZ3tfUU
Hz3Y1ay++5fJu457HHP5xBao5mJsSbfi42gj+4NhMILs2AF/ss1OEy8pVq+9wqgy72RMU7XULFvL
6+B+qDPxHAQ4s0KcDFi/e4Lz43VOjvmwyLKwJZg8LHUV6L7VzmPc3ReAHs2K3O/4O1RWJqd9G6Tj
goASEL7aFsGujxRRl/A0xUOuy9nbdPVHfUQfS0hu/5Me7oZUMLKbmXduS3b8pwj1wdIXVsCZzkba
zVTBAQlNj+TS5N/3NSFTlSFcPrMvwmy7+NwXn5+QB03IQsTBNFUll45OYF9PUqgBoCG4PVHNQRFd
qe0tsbpd5IRz2CWRTSk1nNnNscbQMsCS90XskDJ/SZEFFB80HTck8EJKJu6wjSAYYohnuKBGg0Ph
wBZKgNOS0I1kP30G5HUyE+Xcsu254iE4jH5khv1n0Uppjr2T3J5VSaJwyLLiCguJn5dvE6cin0O1
7bir/wAz1g9DbhHhlCi812u1u+/kTDxCvXYsxIwy5bm7vLwZhNEGB3M6VgC/NgrZhlHgqTUSNqwQ
xwOuZ8AZfquCRYW8NnVegRr7Wq3x7W1yHEu3+Uz1hbv+JfW/ibWBX1477DE2vK3Rc0Wd5t5StBP8
43cov1v0Tg/LZrxC51zg11yrU9VRFdguFGL+Pi12okio6tDKwZg3akh+d0ArDwIprWKXsELRf8AQ
Xfao1dbP9zyo+VLHLqjP3AOhO9jUFgc5jnDKQnUSt2HmA2GnBTjGz+Zx2AHLEg7SxUnNNzS74DQ9
IxuaQJur/nBnCBWVv9hoJi/qL0MvbKl6N5IOdxil/mp5GlpVoeTjtO6fXV0ULTBPJpCmv7fijYVR
567liL6CsIvH8J9obdPmg8xzlVZkp/TFjeVATh2lCWC8+Mv2UMZPnnDMnJ8SaCyuVtfO30NAceTK
FYMR9Vl54tqQs2UAIlmH+zBvmSh/sCf+jqSTcN0Gq/mIYloK6M5Vu9wbvZXdTwanNsECgopA226l
MR3402nZNetip23uIw82Ma/bPElwZBQGNlZ/QnQsW9sZ/wO9S5RvcA+mJPGoQAjpREbM/1tB/EcQ
p8o26mv7h4U2jfYmh2e05e0WiGkDyg2OKcZDpkdQkota3whYutoq5NcURQZ80WcBq4Gl+TjL4dhp
heNDDTbhEBII4jJ1z0ValV8i4xbrE6gX/AK/jbPNkl9NDW7B2hy9veyJzF6+L3Y0IFK8FCq1zxSh
r+g3TpMLb1OldVrs0CYLVepXIZau4d98cHT8XYThJx5DMGaOA4V35VHRyJaQxTNLzCBJr8yts3LZ
I1I/2x8M71K5Q8UJoZpPcQVmBqhH7zHn7uccQMmVO8rB4G1xT+TfLnI64GO2dXsOlhmlLwq3Tiin
SAp7ZyUq6s7eHwrEHmhkcO2xidiFRKTotWAsFg5mfgdsJw/zrrxhw/qvx6kXLPNSgne/FIkish8h
Sf7yRaXmGemBsBU9KwX7+5+WpfcRK30cLVjffLn24UM2l7SzVMHK0lLY1hp/vBRCTPrFEWECxtBe
PlBECybvF2YZFZYZdpMgCAOAi/0Ca6v36qjKvXmgZoBU0lIbJQI+PeA7EV5ZYhYC0JY3eK4q/+WJ
9kGLIbTse9XNNqdFxdOIIxlJfn3N9iwwM95wvpVTplUBqTT0vv9FsCJIohvJvauCFnQdI3XWD7HS
qLBlSbW1miYJm/RrJQ8yoAokFUlbMMXhy5vP53M2Df1AxvnyuEkj/O8tSOGU0YS67h75j2kZSKkK
cDO+WKtVHB2vKl6UYfw97xeIIMk0J3u/7wxUgalzFFxQb6jL/I4c6v0lJrvlw1lldUUvsYlo/u8I
aRfwfEUN8G+YHsCQN4RUxV3lVcJoaT7CGSHQ58iRpuZ1Lvo/EygFgHID3rnLUHcow42HAnfovqUt
LfDyhsQWFwv65wmvFg5BL3RYxxZr5rI6qg7UrLMBh2AL8Ac6wmA8yibIM+/kKyhRjmlXS921rHgq
tblDTnUwBhsc+gUbYS4R80+fR+vwd8p6hkrh3isYvsOP0s7JGn6GhR2Dda/ftOdiUz73AxH7pYCc
h6eHEWDF5HRWUqHCn2JElK5RhwcW0H6ngdVGnMUuHR39uLFJk1ZgD23q1a0cDAcgP4Qxci0XBfAp
ItmB1msDYbv5nZzba95nVY5YBesJ8uP2zqoBcz4ijGRUlKBIlCr0q9rc60p/Fp7Plh4VEsw0B5/l
BAfec2Q9DxVwa6T8FVs0+dhiE14UKiEYdRrPtpvFTOeSODfK4ShcLB6sSORac8topVJhK6xNh7fu
QOHhIjiit+SmW3Tm8+Rn54gXYcZoVFwgoTF/HHcv7cGsgSmJbNwOKLm8N0YP49+17bPVKmTpIcPr
RgMLHlbwG2k02dmaUhACEnBpAWEJ+DqsnU8COanNuMjrG/MkaiKU9CpcwY+oBTlWBGSux5RmSLHr
t6bs1DyuMUeaKWiLMUgPSmIwZ+Isu/b5I/+OR1TwdeFRELv12+J3C+lUMDNjkk6a5uJDPhQmw3ek
55UlT1XHOPCIa6GzA364Y6pBJNjO/mU8qW7k17qZCtbhAZbrwDb47xLIziq/dCgcn0lw88vaIDVF
8niAYuziv7STDJg+OqdSAaoRYsqduIj6zz7Lg+CKb8dR5IqGkUXw0u4YgF61PpmPcXoUa87WinnN
0IPgIH4aUo5Ce4RCA/5i1f/Eqsl8yPOG4KCt1/OsAOHS2B9t+nut62VgUC32oDmT4560NZAPTQK+
/Mh7k+F8j2MYlqEOz4sAYIQ0juuoNJNbJNCinOExXVCyFxF+izKpWKzJcsq6H2Og8Zo/iVk6zI94
Th9iJ/34Bv3rf4dQs9IChc+OtQW04Q95QgPIPBH3qGoY18nLQgRcDgO5r/vISFUK09XEpk1n5kOK
RkKnTR4MQ0E3yjdgjpTQJlpoNgcKw7tLw1wX6eY/bPXECbvz7wYS/jXISDZmPsmWmHgXcNYNH1na
EarshsBBui4sAdTgPN5q60+TLUP45V5YzwpCd7jSM59F2oKyPgsi+4W0DMdBzpYflbYMP7RIFm7C
ezqsTXG/rCwHSjm2OVr39w0eOjxrgqWJXf/ceh/dO1dr7MYO6Hg90KU7Ork9NA4qLNWzipyKe3H/
ZKJPUp+XQeiOzy8bQOfgxngWjaQb7Kh2cfpiGJ6Jf0y401kGc1atYQSp1bMh51pVLysC2VTMr23p
UjL6nrbZANGl698New+8lhDt+QDO3p0CiDCNQQUhV3u6feQpecaqO4/WAo1CwGduapkfgPv/zTyP
hwVR+xe3yNhyczFCVxevd80W1U3LAspcZaPiRUJB3eS8tp0piBModWQzWKnVOt0UqAt0DIPm4XoK
Z1WQ/Je2F/6rZtVXEy7NpKmnIUV84nznKkbZ78UpqEOnf1RbPV9ojlcaXac9cDq7epHp6CiNuuqY
2JyEJI2kUTJFGm9wLtc06hPM5oJRW5/TwtWbArV4n4ExlDWpmx2wcdX/TtaWPYVu4BtXTLt+sSiG
yjoOjssjJRBweBM/dkbADWXoUduuEdZUcqf6Sz6QMxoQlX/F6W+Lnh3jM4Nu3Vd1jDQuVtCSTM3V
XV/jn46KWmJ1jgwpcy1xAY1o/PPsI3D2VewETnOPzY5h4SyJKt3RrmCaTVmCoeitIcsaembaFFak
4vcFoj5xrlZGOCiceuimEWvdKtQkMntaZ58uyyIJSnOSYCQjNGCYk8xgjshSB4qW3pjPvphUqIdG
9hJxJWguWMIDY19nftDzX2p3SHJ83TjQ17UNy7TOsrx8MeBCXf+UAl3J8uzEHZkV4S1qHRorF75+
CX2Ej5BBHhgiOugoyZviSlKWwpWlPqqfqimgPBrDXTTlsL2npeapdR9FEjQi0gm5DuhgUE4mrqRW
13FkXvl9gRxt7b6LofpTi/1HWZ0+t37zrGrHRjaiCSSNoKPfHHHaOMt8nO5J+mLMYO5LFA2XAam3
8Uutt87iTEvh7hWCamyWJ95fof2OnPZQQfKp0QAvfWTS8kiSNs7rwqLl1TnRS/Y3/Ngs5horzH4/
v/eO+5AcHKYBr8qLSMFhAoalHtC+tPLU7/3Dvodgc8zsNXlmZ9XWB/+MeIRBbAiM7WNovSfXbonB
sVJhqt7UwwiBJFgX42qXS3/LIqc/Jq1poL2yroGbSHjlUpnA3fCYc2NPu3wiqlpUbwiNQ2KweGAC
xN1u24jm4MFXWAXhy8teP/vAR5gquOEq9prm1r3940fekcdM8HMgKS37di1tOyAdqjy4aOQa2I2u
LhxKYs49kwQROWAr93QjpysXSX2Qz65FnVAdLsK//SToZix6cEWyckni7F2UchXT6iUYXf2evm9k
Zj7XGq7WQKINzyBKTvgfCUrLiRn8oM8vgzJ6QbEU2r3tr0gmo9x/s2dqWSQAU7u+/4LukMH3Wew0
LriZmBLwZhuh1M0kCsMun0xsvSjGH5z/pMAHLFhATEnLBNEzyuy6CCJy1GnlgT19QoE3D9S0gX08
BiYB3MHJSAG/kvQH7ls5jjTSdhRWnYW09//VEECIMP4s/MhrqGkCj15tqT2RtFQQCMAdkK1GldCc
dgocUpJ5+Tw0MKL0dJWqRKTedry8kWc04JjwWn53qOtzXv3i5QWDGa2USNonxqOhkhoR/RwnRfLb
OPrOaXqEEshhnlvH8X1V+MTgI6K7bA7KpNHXbxpuyl2oB5sEl18Toua8ERaQVGUTVpbQyZ6AC3O4
ske1maQpJW1X1AVPzvjINCLfrYn08PpVhnbb20yoVCy2n66J/u1WA4ZddjVSCXM8nHWy22s6hcxG
d+Qd+uCVziyyNh6l6NA3V5CLYX9GEoyURrlIl/4nnaCWVGgl/T3Tezx3uApEgws4LoxSF34XNmJB
nFsL/q6iUkjM+cBBS5FgPuuwKAVBiokQiHs2t3rgTFtKJygRdBjYHq7SCofYZqQ1ndF3iP1wt8v6
p9EayvYgi2JhAZ/glsUswD/N/ICa0WnMIehmLjCPlOaQp85UB9t1M/0I9qUKlwL04/wL1Bpzlhs1
bwifnZKyunEzUWMAy7Y4R41g3drb2kXF8/eJL3UhvjXMRuMOzaWuUOsPWIh47TafkTRnkhWctPNP
BPErgwub2YSbMXTxPvjX+h5CBhaWkCg27GTYNxZkmoOqhycY8EoUD95GQj9TJ7ENa23IBaFF63w0
FBHyqIu0k/tPJHzU6Rwy/QM2QmRihRA/PZZc6LtxBe6GVu+EdkFTy1HhhoYLvZ0cDc2FbscZZhVW
VV2rLO+EIu6lUWNnf+V8VAaIsBJh50eS7UpYhZcgusPfQRjkWonfxvmWsl2AfFAMCwwfyqgUlMhD
wu/PjWv4/M2QSnUSCH+dDjtumSTUgJrH07Jp6AnIbG4r86AVozjJI5HpViJoqhQIFEW7yZfFRiI1
GKjVHX7b/vP7yez45mp0Yo5XlHqR9HgMsxA0LQcNaRIWeC/Fe/fUbFp87U8yyYUeywjE6u5IDnwa
jqHkKdpQx+LebeKDEtiXHJkffLLQ+A88I5lohG9WHyED16SQWgIWc+AJdU6ZXTbhWxGMmbdwhDdd
K0AFxfTb8XFJgivY5cEV0d79z1QZx0iMikyz64KsWYd74MJFZY/uZH6oCWhQH1eRckSrIVLl6tNR
0V61Qh5y42djcUg6UqxYQRo4Ibbp0CKjz+AVm51BX6geCSQ8GkRZXhaI1Sxbx/lxo+5aGU3jaUVW
ff+r3CAiq7gaQrLVETrQdJRnYNeLidbP239HF9L3HHTFc2BEYm9k/blgFPXOfG71nuXv2PPTzkSQ
Oq3g+6qMxFcL2sQFPE5c7o0cNL033xvHDpJJjqUOG9oGbfcaTTPasQg5K80tdC4dbXCQPotNYRbg
lRn1O2HO8jjFldHm11lp0ixlQZymbJueDJedTgDsHsZbXCAxMKjR1YUoZv0hM5a379mLgmBwb3/n
1IILfNu++//in0VpQemXub7RtfU/eB9v2YfodSE1A0Mcd5PsBq6IGUh6uUtM2Tje6H5Sgpfy3+Xc
XoP8zkLHgc3WcYiBIzLpiwXLTub7+1MoWKLkm0BAZSA7mZLKd3oNj2sFznksxywsLUx3/E+kbk3j
vDkx/5Eogx62AfWOF+LNM9UE6zdTazjLN1pT7uBhS6z/PMCKjXxs/bIaM7xLCHO7viXT/Z8sW/v3
DxSBLJMEIPWh6iK9CIwDZV3GX2K9L41zD4gK1BAW+A2DNrYuTP2lEX+e7Lw6j+g64OKblzZcrPIE
BBq3tGROUSVy/A+uEaMjnYtV/99+a/YVtoJ7XfrFx9RQhiEjhtU81g4cFf1n/3G3tqNXMiJDxFWf
oH+MihuPMwbZP7TP4yRNnCi11KK3A2HPBsqeCDUe4b6Ks6p90tvMPALhtlB/3AKxzfJ7S9xD985R
VYgyy4+CPmR+Ys8SRoDLJ0egLgdkjswrv1CS0pP73f6H1StjDVCQUXGbRVbJU1f8FOmhESWDD2mG
j3uXc1UZMxg5QPhoy7ahjTP2GDm2iGJz0uXStz86Gd/Dni8qA7kTSTqgiB2lk/23fP/tkkN1U5KN
PFadaPG/4iYbsOaej9Xe9pLePMr4P4DPvKh2vdGi6k33aFjuShZi4qXozM4S5ciR//rYFN6v/uoD
AbanKnveUlG0gPToTvJwsDRGjN/To9taozTHT9BbTNiSl515o52IBYfFTm6m0BfXVkIUYXcBX7FU
xiVRsCA2fSulLsHK0HfQmZMcu/V9hqvOjT0KZ4pa1GuhU/2jqc1YeyMoBuMn8F7LB/xNtl8fhCKa
bCFp//mO7z9h/sdP/8Awiaf5nR84AIY1OZiIFcvReRHw3oepxKIlTO+nXHEDYKuSszMWxEXlNREB
82PL21flwg0fS+hOPrbiCkVunZZaPvmnsoppgdvhpsghue1FC+JHAHfd+moMdCQm9LC+uDGtW9c+
bjoSQ2MP/T2sgg8KRsHGshJFgEWH040lXsZ+VnYf421V4S7UuPBCnZZDeexKOL6QwY0/53ZN1NMk
fhvOGXrBYChUpubALc9Kf2yThWOeRJgjfmv+S9rOqJ93iK31yN1Rd4Z+a/SEr3zwdZCNcY4GmI4J
lrGPG7Fp2zFvHcN7nQ8WiFdvTtPi4hyDZdGLxXGdKrEeGlXVIVHGv5+wKHknmHhV8Y12DoTMN4C+
JWgljsLY9BTgZqa9kjWD0+eMHfvuq+fbGlTsHZCOV30xoQyinwW2wFi72KMQQQfaiCym70HyeUqz
bQorNpOqPqqhE6zXv+g6nPws1WiP2LOrxdTRiT70CRJMwMg5W2q7sU8KC6ABaH3KewMDrSJNFmkM
oOZ5brjrTMQQptklo6j7JTMTQ4KC7QRPxp/7ZTAGPIyIgTwkLfqfVdVYa2cxdeflnz24uAwJ0oxO
S0aC50XuONZ15YQSV81S0nMi68WNmBx6YOlP7S/7Kl6cTaOGJ5dHBId+x0o3Bvkz1v8ROuDzWmFt
K2faDAqwLj7ssR+VMW+InwveLTNaiNcUitPVrkd6AmNvh7BahLv85uwAsAVZK/l0SoiwYvdaRIEb
2ph5kQChmOHdrZ3chJDV1LW4SF7vXpgDs/CZmHA0ezu8sk1T0KQe5o6cPxNLSkWVplDbzRnS4TsP
WpPmUD+yooY5+TOwKM7xfu4rgrGnWLMGmfiXAPbsixPZ6QSRwi7eqIOO2ibI98rCxp5aYfJZsxQ7
CdW9Ezr9/nTLMTWGAE/hBhkQvN/ZcO7eZKE1g9zsyRIoUEqddvQmECGtwJDbL7UWWYysSwtMd5wp
4QBJCg5MNme8wMtAx+kjZhm3DynvPN8b0IDSy2/G3tGsI7S+fxTfYDRMXgx1BwTyXCOsI1Zle/pm
5Rs4egdfdWdszFS9q/lgQXO/OPYd5QBIe9PIbSwOlJBsX0OjIZteAeARcXFGvTDCT+2rRNuiGtl8
bVUy6XwjRmyQ1gv+ROJM2Uw2Fd3qNjaVlrlWcq5ukDhPQGuUZE+3umVnRxnKqPIEdCpxanMDw2Y9
9ud6SKsJxMYZUKwmFq+SYtmThHJp9SzxV9sf/GSSGvyVZHO0j3njvxMHTnqJYsMyxEfgvkf8N1tN
mdKXAq6aAScaDinpvemz2ylTrn+qxjE7sff+jgNlGskxR8GmE2uTMaXbR+cagWbIQc3N7NYJNLHU
xWeP3+Qk5+9y2epiUL2mcP9io9y1n/7zQ2YphX//ZKDTz8Kpc5bYsYzYM1EylmU1Op6M+mr88syF
K+1ZLEOqNC3HTO6SZ1MOuMQikJOhF9X/oqW9lAsT2KFE8STfMPOcZEkj+5z5buvYG2n0sRJGm+G4
ngFWNyiXDqgVpW49+n44E5IkR8GvXpyheWRDNkUhkZbOUHwSHZLpHgUe6RmfhN+il4zZut5Ky0Wc
H3trTlUAxC0GEAsHWR0yezMnUkVZ9r1cY1AnBQ1Ks5ZCib5TQQtJuPZdh1FLw+z38I9qYJ4O622J
K0QXMfe4bEBuVLLRHu5QX5pm0XqXeYF/m9D/a3IQoIJY2CaXGAsAhzBtkhs30RFsmegZQEpN9ZH4
vhA3A4eQa/F/wiNYVyjhauAfACNEWPnnrqos4eA7kpYgaoRfQzbKnuSiJ9SMLx/S6US6eO+yZHD3
z8arIvfoRPypv5q20It05XlNNVjf21ajz9HZViINjx3cIorOH6/Vvpzi+QVyAhlIg+7yOcp5UdaD
2KDq2qoQ6rhmiL7lpZjHNFF1PsFPBw2h4WqkakwiRE4KQuV5jgwtSVINGNb2x+vj5Nn+mgqOtjDD
041sqheoZoQ+7tzGUPvX3HVFSPBLj64jlgD8w0XitKMdJxmyX0ChvsKXz5Z6mpsb/D6ZfDX3EzaI
KA/cTTR6F/YgOjBCGZ8gtyCsvXRH4OiHtSgtzdf3Dx4R61SvjNmuQZvQ7SWgOa/Q/ofX3C+/JVIS
JJEYXrJSrQboiot5R9xvgLOLk5oxyN+qMrSzrrNFrBmHygMsAAmUWDiuGN4un6rh9iO+J0m7twnp
KJrwD+nzqJDdyjXfAzks1eLUfa4tngWyTWIRayIJmxE8M4Jf3hwzSTWwN9C1nnvHJ2ZXD9LEMzg8
hPEx0Ktn3r+JllzyXK321K3uCIjvyTxREf29MRYdfa/NZfzon3FZvGkBUYaIfGHD0wnjdSOoreQv
84Ee5GVoi6yeetATCSNi6iKfoHpg6M7y3EohlldqWSFLoG74L7bZ+FC3aWKeLNO91FHq1EYTuunI
+07NNoRP21Vhw2Tg00INnlKhmpUumQy1CPTEPdUdevHnE2AuoXWDS4hniQjX6szatpfVerDXe16J
DCpnw6lExaZgPQExMpj3yORXAf3ANMDgdkmsL900cybI8W0RYwmysvXx/w/B5LBYyoXSiszacG0S
6IfvPVeDYrd/1oqYjreJrzLnwq/MvMqd58p8TcsyVGeOXix7HWT25xFNlmZd6g4iAlG2X6OlpGAs
ybAuD+Zdz3YCaLINd1x/W2ZibCOOEweGqE+/4bOfSKQ7xWJTtc2UG/Kb/QToaqAoBkQXQv9f3d8f
Ac5U0MBtjUATmER8qbdIBknoflF6U5824x+P6Ljb9iM70ZCI1S8SwCprOKQJVz2MoA4YBn9/mJDh
Ssg69aWjK/257ho0JjFHnhHQALvKRheDuCI6UM3GRdR7jw14bj8GZW3JGbiZlr60jIcD+UVzvMwd
oDyoqP0JVETgfblNCQX9+BqP5+5q1NK+UcqtiH9yHQ7eHpvvqm5rZnqFSomNUzmERXZS5SqDkqVF
3Oo5ssI5uFWTWzmYoAepqSCF8/dIVqgPaT7gJTbDNTFwlykjEm3TJgKCRlj5y/ld7ATYdUbtTWV8
t4fhodJK7j88qn3utJb+b9myiqsQq9bImPDoKLYiJth0AaUzTGtccWa1gySuxB+lnrSTrOJiZYuo
hCg5kbyYn5aJ6WhlPETcZAVp04WbN51ib+5ev+XXGOI93Yc0oqGKpcvXrEFrzglXNgqLPuJUjQL8
dUKK0eXKXPD2rJxj059dI2hppExa79XWxYb2bMx8B2dFEVyn/B5iQg+5OGpeaUTK+46XQMjlVaID
o3pq5fAGk6MfqxmJsGmRjaBqDrEGe84C2UPSc118YcH1y2Wia4MLLxfY2GNcl39ftgjQ/axyMwYz
QLIhwR563NuoVJoXCzkebkQwNh19elFQViq+dzBKCfPxNC9bV0H4Qa2VWlPQHyPh+pdHirWZ6470
mxe+8pqfgSRVOqHADFb8ynwEwYwp8bAXj8nK+AEiaEtFEVdM7Y+/3mL7qTk3g7EmhxkMUihKkcN6
yb/gAvfBaThad3clcdWd84vPkkw6RcILKs75JGUlk/ZNmz6brCc0hWW8Afujsn5MS5omJKyGguoa
CA9JvAFKJnniEJ9NeE/PK6WmZRA0ngHEjJX+NcRkfSzCRndIro9/mIMb9+rXSdFJzMZR6OdmzghG
ZFY1lSFBkyz4r7wKeBtgk+Xilcgj8dTITcfLx2/+Kb3FW5T+gEv20+Q0zIoB2sH2UVaQbZikzUa5
Lm92lIah4Lq6asRUFuvVzZmHH3SaPOluIzX476adOn3hloiulSmUn6OSSqhtQChSjUNt93IeXSyH
kvLCnKLawe6Kq97+HBxzO3gdkTzKVgXeN3CDGNObFBX2M2xXuu5l1lI4piikzrT0SwYAHO3RXsmi
3TSqaBM2uevUjpOLTEzseWeKqO2R+lO6SgydVw4XhumLQh6CPXWtCQsqYS2pMDAMRjVUTM4NTUB/
jyRALqogDGty0AwM9YTBcTfNN1jRKDFWmiTyFpGk+GDws9gaPg33II0jX9WBn7Xr5HhqN5Juo3Rb
sTsiM278CAMiFI6oiCJ1sLGV7tDVwhog0ascBkOWGYgT97v2dfTkrkCm3JuFm8BsrRlynh4Sg5HA
WwB0LAWxnyhqMuOcbGg/FQa3xz9tLcexhkkiIS8k97qN5EEt5UPdg6ScjU2gTWfVJTk2GhhGyM/V
z2NB/nmdzrq/Tr2MGcMBaLTYB2YUr0iLyLFs9CEUisUg+dK6xo/NXGAocCfh/GTisHyhFuiVXH6N
ginKQL6hEBzuMpq+lu+cMHV9Tcsy32PsHVBi8h9Y8JqcSKjYRl8vbIczyQxWJ2jdyZbwMU+vyY1B
k20c+tHRH6GE2GUfWe7zg6cMCNv0j3rCyRTIWL+palco4oOCahQ9fhzOsXKS7ONcC/ECPddJYcss
cJt9pic9LRAAIraS3kuYXJyrSqmP52lndvSiazc7QPB2vk25SfXVBwN5Q8hwS16b+GGFB7paE3Gv
efHOGNykpW6JMYfvtaiNCxntSxJ4blKGXM+dpJdHhUl5Cz5eFS3fuU7KBtPG2eq6PW/EEmiuSPuQ
BncIftYeHjo6F9F6IfWk9pu2AIFC6TWzuulh9Ij2mY56UlAxH3zOpQvWRJY4fJNK2TGslX6rvUBG
++3tqZrYjTXLHy00Vo801JY+IMQLRYgBSXN742nscg7vvRqjQmkdV8NCGCyPUXiFjVILYwqzENiQ
hG0BG/9xxWiADVqD1NpwbhAjGJY4h/YWkG2yu9e2m/nZg4z4jURiAEfWQv0Rlh0EfeQ1pQQijWBG
He4QZI7T51boKi0Mbvm1vrg1/9kHuplFNVoar1BUbnT1wKDrLJjvAdzvACDE3VYkfhZnjekKFekb
LDkELs7cw0PbCwFIrTmipFYfQIH9HMrnTE5Ua/pGKCornEfSZ+oiMjkdhWTluLt7qQa6nNVIpRvI
8xto+boeb1tLlIzebtpjoaYyR9hH9KqVcPPe765P+s9tnKU92c4PsxawXrfZJ8JnHB/yqJ6e2JsO
53MqmMcabY8OYRIw2MRuy6Kifonp/LYPfdEpJx+NIEsNnqyU3+fVnpxAqECqIn8B62gj8uEc+c6l
5h2mbSmOn4OEyxFpEBjiX6GRXyQ1qN327f/A3lNYkFc6mrq2TLb7J6kGb3+XF/V1N3u5GQVlVykM
9pulcuzxNsRqHjfVHKbizWq4xxJSBKg1Sozwm5z3Xh50w+KfDGcMGKipSXG2TpSZL+wJWmK0CHBu
AxlJHzY2zMzQT2t0XhLDcQh43nKBQRhqZJ8vnw3+feBVZzLrGAr8c5ssVVDOCzltufqZW0kq604T
2dyEGbYpXv7ZkqhzXTOrBimeUAi/8xsBlZBySV3mvPejbs51DA0BI7MjUDU1uNDNFbgKPbtyjcQ5
jS5Xk7HTK23pduYsSutla95yG9mmCXoy+LhCO2fNW5FHmk+fg8uF27NIRyoyJGaFjpSeXOC4BYh6
35HmzMFhujT5nnPJiJfTGr4USok5tiNHFcpV8Qby5bPBU9cvoasl8WlVS8k1vl/ZcT0TUwxhT1wf
ytGNrMWAI7qHTTzu4FGgUAIi+/jN9mCvqMRpN0VQEXxGdog1XUBz4DDzNFmlNdGDEHD3UcZQsVU/
xHu68kLdMyBciukVfDeYP/CacGz4OxHL7UQUbRBXOByNvuMr1GrxzIyark++2AGRhHMdPJKJCtMG
clHLdwVfB5dmebZ/Yz+G6ryilEvrBYDe3Xs/KU591g+j1m293h8n9lX/Jb2X+f7KwLhyapLHFQMf
rABws3BvV2L3E3K5S2Kq4hvTzPDIaKHbkWoQK30ODqh62L+l1yvxix6uTgls7MCv0h29MJl923us
oQaJXYvF7yDPjSJb9jFGAy2yBEGRPHg8wsjkrcYSyCLBEXVAQSqmlRXVCralcju7/Nb/8AD9nKQq
uEMxeSfcApbCv3i3Xmo2CQuwpc5ACQquQiWSk+b21D4ugHru27RHN+DbwMDM9OQYM2BF8woFcaYm
elmM/SLXIx8lFRQW62/7ymTP1q52lJfHuUtC910ITp4KOTe/EozTfe450nhU5kPMTH1Y5G6XVxtc
5wSCwqD4aEtIJPjhgOXk94FwDyVWwdfPbFcpsll6aoxlspf4RPEnc9jY9ZdkjGqAJtfywB6AD1vN
+ORmAEkmT4RA3HcvfwiVgUQsqGce/hGSdCL7S6aBHi8jB0lAKmLS4SlfNFHo19q6KhwMglxqtT16
BO+FKojqWJcn/r6+bNTveF+LpnLM5BVhL3z9PiH7ppg5hqTKtO6UMepDgtUr2LdrWajuKM4NmEoL
SiL4G5BV9IQ+mB5YdUloEpZTQRaxCQiuf2X15Dgc/6glq7xem5eLgsu7UPw804/54ZZroNDrL4Ka
S3SVYup9gF4EGRFgbkRhiqxkAS5e9qJUdkdkNmhyK0NXGN6DdZpuPLUpawjhbEHUWP769weSu6pv
pPBbts05xU52peh0jjU5eA5cYMMAcxkUdTUqhq78Y08fwxGTnBsPIxSSMkGQODWQECofolpshu5t
msxX7AABdwpntMTnsHmdm7V/ZQTy+XkguxBQgFFr6/zRZ+7MUA7RoDdKMq34zH+17fXTfc9gchbl
3LkN3yG2kIyf7cesT3B2FB5N0Pz/WX77AlibvAH0iFYrTk20WqmiqPjpW6WctiswClqNzgdwul6f
LPjIM9MFZgZLQimrxGIL1aQ2LpIyEJqhaw4ICyQvZ04QwV94b/QWZ9jHUpzR1f5b7NtrMqz+SEUI
3caicgl15VE4NWYvP2XF6oSY+a/xhsyfbkP8Tqo8kR20lIlvoXQpSPv5jIbUGFDy1TlxyR/T2DJz
8GEeYhkjz01fczaqukgNT+2r196fNNAQcqpJnp+Ip6sZuUgfw+xICLi3q1A533cu9AW4YCBUrT4o
R5VJv0cevx+8Cx7Z9zvci8gPbILqffDrRTo/uymZ6MH3dzmBv2ftdzvM/DzVUXcZ2URCuOyOSdq5
iBdB4ZywV188y6de5ZQxGOtYzLa0H9RMkt967Q5pOC2SHXUWxC18JDsWTMGtB0JtmobUcFL0BfY0
eQvaSaLzcBsoWHBjjywpzKQAVdcUI6DC4QAaTWsWlN5MEogPn30wK0/vUrmjWDKp8PuPQOM2fX03
hgsRVWrvAZEpVerwN5MdVBLVaALvMK22kd0EGUxeH7FmFYt/myLDRm7Qw5L1IY2zEx4jokG2/mvB
jtL7VpfVfsTOcKXON6y6adR8h4pwX50ZxDcrOmOQsNP81/g5Yas7ycx9c2oiZqoQc6XgJAjOy/3A
DzT9A2rvJrWBIGddwZ3QF/JkCM0bfOiT/bjeM7oLuUx4/LFQegN8iASPUzpiT2tHfxqqRd152v7+
Lpm19U8f0zOShIxxnYrWddX3MOPyEXJS09lXKoeDA5wKdb+4eZkhxSD6aqeJHluU6mgGbryBhDMl
0EFW7LyT68LULfbKVz8JQknKyZb7OTwY127R9KUHnHHL8HuN8a5PxpxrCf/5rfb5xW+z617rYv6z
j/toHByVxNdFZPmUNmeoZdit4dhOtUf7zsmuVF/KCPGvv7JhdYvlIxYXc+5G3LIrMLYaqC3QeRSD
GXVi8PsdD2TS02WWBFhJKQxmhozjvEDwToMv/4Yo7HelNrJ1rTX5/+wGM17f8vblCysoY+jqha3v
sFreTiykHYxewirQZEwj5ctivvFNtafwww8cBwqbVeGXRmn/yyTX9cfaOPBHUr0dDAMIOFpRos5/
rV5eGU/cv1GxJkj8fy1g8WOu6rEqKnCzd+2HwRU/IvxRAE7DFdc0kXFEfnH7VicxV0dy7iVZKC6h
vQQnV9DHHQxtvRy9BvIsc0SSRClX0IdfMSY+8qgZOule82F6F7ZFLC2jX8vqXK/NF+ZXffzxEGIk
FYqqiNpc/RO6xmq2gmje6YdMGEd3KWxo5J49VoBGcAMr9RlPUmIt/CZtkLdecKw6B5O1HfAK/uBN
7WpsS3PZPqTguU+iTriLQbL46FJEUc6vHZVVAALBEHRKF2v7H5U0BcI7dNWoEIQM6a6IIB7pCsdo
ZjcWnWcdlUt/NVwBj156z2rfoU1huhe2oHsn0xE6aJ5a9/M0AeUlj6aoWz6xFtiRy1lHLVyxfKck
GP9s/zYxjCjoYgm2QrH2FRDcvwBHA+qoeFvs45qokbLc0iiOH6iSY6pdXNw69A1C/7MFQioG6SOf
tNBVkAsBXA7Pk0AOT5hQj4iVqMUcgJaMDpEu+eJj1qW6bVaXCbbFSFDpgcscBuwvs4OlbGmSrCeS
eDHub73BLPIG/VFLhyCjXp8gQ7077SIKDdV9pNpOjAsw0YB0zMs9OYbxKsV5k3MGMXYQr01dzLfA
uShwnAE0MnQghJX2W9wQoHBbBVQDyRbdMZsJY8vHmePUxeM7yez1HAnMcMfLYEUukNaR49Do8/Z/
5UuWpbp19AMCNj0dlbCu6dNID2k+MKIWrBG2MVgUZdfam3NbD+2LLnzGdZr2sCxqC2Rq2OA6sscJ
wdefwyWH55RNqXi+hp7zEhJpDdrfIH0E1yTLoYS+KMg676vcLKzQ+6Js/PbGQxlPD7FAURHpwKt+
XoU7GdFXkepZ0FUh6/2yG8NolqvkvtO9ynfpbZDBtF0h08EYm4Uz4blKAHzeV8q28rQEiHikftT5
QS2fD5WfnpoTWK+0jdAZk3FuAr90sdhSzVyut1TrUUlMvEiSNH5PLJlp69vFfTUL6pil6oFnxObf
YHlGsnKaCMDXYRSVcKlMq9DxreETEFHdGxd629XK7HNbUUvV0Wx6ZJEj3cBnzMdWuGXU+fhM1hIz
J0piMOZpkWMEeN1+WmbzjNcWedGXa53hH4a4Rin+crZVM2V/8O/h+iX77HJ3PROhKbBdBB+0eSHw
7VzIS3749GW2nMDKAaHXAtyr1TRpTEtR0+MS30boaMoQ8O7aG2SvWc8piM0HHUO9LrlXUSi3b41F
sUntEQ94qYOKuUFgN4diADiD+NhYOGcXjh3dzmbgiCtZPicgoaqV4DLngDeHaKQ2ij9panEyIJhs
oeLqjp1O4M7Dk0lJxYPluSo7Yuvn2FU4e43gnI8Nh/1wmh4bIJ2RGldocpmerNMXyQmMlCGONEXO
Q/1R4AiVcJfBjbKJMEmV2/3IQCKpReHq++vq4zjJCG0/EvnTsyrkjWZlmMq+F+5cT0uY2CiARskc
iaR/E1UPfTZOyE/tNv9626cjumsSVsK9/jKp4DQjiZsWxqS8sdkRWTN1ct/+rAsc0jBChC4CB/Q5
9CzTaZ9hUrkdA5oy0fQmTRBEwoz60kg0bXhKKv6KQ3oj7SMI5RubWM0tWbMu6J1ZMHHiGiVUBC/7
weB3nbvwgczUaF4sAwJTwH8WE7/a2xs3wgQ5PV2s1370lxZKfnihBGKYWeP/TfCBSNSVd8foIqVK
KgEIqXBrkGVc+36zW1u7t6FXaB0gxTBt+2ycRmly6ukoWMTFSV9XdhAN7obxHpDyQoL5oXZyyzf6
mQHpskRF7C9Io5HxGfCeURinOBOA6sPWBCiRTvBTzPzRDib02J7GWxIMYmMogIXdyxMSAvn07RWK
9Bws1ez3AfiZ2gaFLAj43ZBi9HRj7s7bQ25H4lflZHg9ssmIrDpYjaKFynkt+RJ23+h5ytU6464H
X4LLyjPEEaozrDWRs1rplLvqzi3mXOKkg6oRw/R24PPlhWfWftjukMVJlSIZzwaVfzQHSKWY4Xhy
U+gkfX24/eD7lD5Vmt2KR1JCq7Uj1eN3iAou0K22NTfUI9LV9RXWyyCrgf9AVWM5QepYoS/tsu1O
0LayVYkIOKyq5lF1h/5Qgew5ceWbnNTGQtR3g8F8wS3hIYsfvOL7/JT71uOtqqiPDILhGTd2D5QF
x3mvlJRcErXxpN12YSV4AhaYuU3hEqG1FlURYkpWqPgmn8Jhs7S0RK3mKtO6dPu1XWBvvCLDN3Dj
ScPRM0w1N1156amfmiul8afeOQt/2OKJ9mmxVIi6r/2jLhu3Df3T9oW66B1Nhav9fizNeHJuo+8c
c4EvJMnWRVo15trfhR3QY8HF2ah4hpMP5PRnPTKc2FDKZ6Xl7ApmF6ukqIg3sq3NDCzMOOWWhPsY
nMiK4BngujiNrcpVMx6jOtXR79Ns+FJnRJBnZURtZ8ZR+lLoidqG+qYr0uWRw7tJhN+46gvdP57b
Empci92frE9CoLiBGyuJLOHmALFnmOdtnIqS2Rx72B51qQydX+7ziAsWEuCvQYgjNEpmkK2txuPK
V1Ctmy4tF0aJc3C2BTgAx7A+UeWIa/wcb1j/PnXqRCUfjnJErL5fnuUY7+Eg4tNwctXweyJUyVe1
yZlhNNkY3fVWuBXuqh3viXo5NSkzrM0q+7RtN0/4fbOX2GkKkmjV1psQ6+x8Y7i3Hq30gW9j4YvS
5LPhNpLQTlAM6uot3rw0IjVuM72QNtR8Vt/tH2JoE7xSRRq2LJEyqflJERMxNGvlrYg9TMpc7TSO
TqwaSaGbpgH+Zthc/j5tyYwuPTB3OWpQOxYblL1jM/DNU0uIxgRKdzv1nlLUzjXAwN2iWxT29Mtb
yWmOmCk08XUf2QomXmxUNbMtID7C3bb/42aGNOswUHIdq4Uwiiydhhjb/Sm4FvZqhMLoM5PtQ/WD
y5V6T45wdNMmkYXQmIYqXu7TMWwuRDBcUpYfERA3J4pQWmcjjSvXYN6JoWEH3ne8bU4jEeDbTl0C
QXvqiyxacz1WYPhl8nNxYl/nTg/itubOQ/pQ8aX76Exjd8vgJr4fzA/0mThDH+WJ/qreksgrLkSE
3Nn07p36ikBfhSFCRTshaFAuVhuSYa3kiLK6uPngSYTOH2GRyOQuzrltmDI6ERefAJ8MtdyelA/i
uj+K4A+HsKhETgkwHVHtlwxAzv+PymjWKkZYI+F/XPaDEWtO6eWMVz3fv6ZE+qco85tyvOnjNsEY
P+5eq+l9AcSu7uDiBaKhKVnBevmfBdBiRF6QZFLCE8rx9W9E+nRhu4lz3shG/P3AAy+DAEdHbRP/
fwinIFi7frVQANGqq/3R1A7Eu5RITutus5sTuRYlpZB2bEf19/2kmWS6f0VfMZgcb+cYOo+XvKhP
/PuzNuCLqzitVdpz0S0anF8A+H3vXYdRV+/DYRIwyA/lqW+cBaGvSPgh5jNnNst78wswy0v/0rEl
xs1cPErt2EVDHnUOqp2MOjZD4IIYo3yI+ZJ3Jq9ZSjqUKr/hm9i3mBQs8x2iSQxhWXT3amP65m41
yRkKLnNBgKKILHD+R/+nWduHRYYD6XEtXuh1dIlTXZfeR31E9O1ZW7wy1GGW6/m8Qo2DDrZ+6EiI
ttU+KPwMUiJmgCo2kHrwdV6JD2HjSurJ91Gas7kxavvIkxOEQ9kuApMe+XI14HYHghTWbcMG5Iau
shl6n8H9RFHQJO/xZlBI3WLPgO5cwaZVmtwimR3r7w0Bq6mg/la+111aBaKb8QZsRmGAQLr9qRzH
mwnBBtoRAUfOwo79awXeZKAkX3KagM1LbLljslqnJkmjVbp5fMW6z41VVarBdgx29JqbmKSvl2M9
/1ULPO0YqETFu0tD4K2Aqe7b+1G2waVkURcs4UcXZS86wZ/ZfCbE4pBx18dUU0U3SU2p2UYn4qvE
ZdDiyloSlIPW+rIeMjQeXugXkjtKWZA+7qr7JgRUERvQrIz8f8Q/DCIAARvYOFog5nYwJ8tt1LhA
DNVl617r2nG8eH1M0u0z5Q9I3fn7CBf+SFTj7gRYhoOy8/sb/CrzLygw3fWl/l5EtrBskaXfyEZF
LajjgPTPymwu8fLTj3zDpUd//vSOedJUC/NXQDNe8aHmSJ2Iy/M1OPHG+pToxt27vHOwi23WbpfE
ye/Al4F8ZArYDeHOVTWEi3hmc9dgzXi04SI6skuaNl50xuhoR77iLmchv+seAusoUsonrtX177Wx
pW30osWG2E9PwZSZX4+2kKxyihCxLjq2VnN0uHFRGo2IeZlhODPODxm5hn95pJPeZPucqDj9TNrS
j6aDbHmd2oGaYFekFUQklpc3PMsLydZS6QT1TRk2cI08CcFwaLojyFKlFq5eA4dwqfGliZ8DmPsF
EXxZYLaUfXDPtgLmgbq/lwb0K7SaBlVeTimCiuD0KLeBJO40vEnNRTeAw/DYMgYtslb+r9traQHP
CDjREgl/1xAdxTmAdRS2mMS8tXiD8ouLTRRK3n5nmxDPbUETunF4u8XlRMY280UC/GCUxBDxpNrn
wuqe0pVUL0vfJTZaLPQFUQRr6w0ZZ0/t6F0PvtRg/nkSUnCLdUwawEiFGxW3TWH5IAUxdUPjMQIH
aBFV0tKGM/mKhAVQz+l6PTrbV1KnfKDa9Rm0pAxSkGbwpHPMicUMPNzlZaJlUarHkN2ad8UHsxRN
iQLs1XXEmPhERORdmW+1QUuMulaK/Vx841WrVXmuVM9lRUj/dIxSbQt/j9b/pYu3WmfUhwn6STXy
7oGl7KX0VAjx17HWItLeHOyC15iUDur896djDumzUoXQZ3xhVBzMKfshNhHA2Bjx9hGNaBvO/IhE
M9rCSXNgmHXePivocCYqUJemBtZndzKCnUWHx2IEL4z81DLS7rqNF7uxHcGKFx09Hgv81Y8UNZ7K
rqQMgeDIkthA755wHWVgVcxxZaFm+BYhm0koNWCE+PxMlLXpJuJuOnyI3VYsWpqugDt+0dZ9+x4o
9eqMpUX3RM9Mgn9F87GUFp9fCSjpNP8TK2SkbNvSTIufxbXiQQ7ZW8ZNYJaKdEmylCFT2K4Xer6S
HxR1iLSbauy0iPZaPv7ZJzWmEnXzocWHMikOoWQNwSp+ei+Z3syQyFs9QywuiBpqXZeknNoiu0V5
MMBT2RW3zmEHJnlQFI1a+rPekLiZrTMg3eaa83QasADpvhy0JSYvasHRsY9kwhF6jkWFwaoMbiHd
xjs95G6lFyjgzG75DTmV0kr6gOZ8JqxMUbuYV39bw3OBD3hdTfT8tOH6imJJv104/GokrG+MxAQH
KYdMdMeRMIXStY2U5zaGkXnWdmurXGeCLd9D1UyWf6IoI0kReMpWNBRIaa2hujqcurLdHoYQGbFJ
TKJMy+6mDPn9hKEiENSsi/uD9ZZPsjAz4igoQ+OJ7g/FBdOPBDV7CiYk2eS3V2N0PqdP+kxZwDDb
kOzFrKlmOyaBFeBCcPUapamJ7fiE5HHRuPJ9Wvy4il7QexGr5Hp60hbuKD0tu+fd3YG5KFXwcBti
u6392Ns0EHRFe49jOqfmoyK1Ux0yiyAGrGKSWwrVpUdt0S1fG7Sinoq24p/tGP+AloDR9sXJjnn7
wopJN3GlCzqO5jIlOeh3idV/6OA9DRP4yb9JbDN6ACUEcIXqhpoc/plr+bUZp9ULwJSBror8LkAE
eOJrIBdx98P2u+VZcPJaQMj2Vvjfvz6qVh7A0qnDwyZRYV7YNQNbKEm06kuR8Zrh+FArMLYNZ6wd
GBmvW01S9hm4VT7OeyHCVOt9xFSfapS4Vz/OVWgJk+DBwThrPQ3oiXkdMEHQnENmksGVTpKVTUPm
yu8paSLCg/s3cRafnJ8UF7L2rnIcPM+MFRc4y1S6pHIXhqwgBL1yFBBxFgOeWoS0OjCpEpi/x82a
UMKNLrMZneGZ7M6WyWBbJywQJX6Qbol6sg6B7Dtwdl84O629Rp7ZU1fb2J/0njke8rppVWrHb9j6
jw9Z9cdyDAoU7RKt7LgufXLpAsvjG8m/1dtREmm0xn/qy2GQXWp4Vsur+tS9jjHtAHqpm1gKekYL
RZSG2wL2vltQM0Lqqfq3QgyCn0II9kjvNsL9/V+qc6V8HBLk4kEQy8JZchrGrC82OtCArFXJSQuu
SDBNq2ZI7M1nX5Fa+DRCYj6gMIuNCR4edYULwhTpld+qT6zzsE328UzdY5EIN+2xcYE5vOQg75xs
7CmvHzfYapGwV1NuIrG2X9LhUNiLTn+6y6NF7dC3DLzk/Vj44CY+8DsXWPlBC349ktqBFqRT5wTN
SX/kXOQFCDJAy3keEbyfezb6bfdyygqSZiqkoWAwNvKCYZWre0dqM9z8Zj5c+mW1Ed6D9CPsX4u8
P/8xFwdztYrDbelMQrZJJuNS9bWaBt3KwkquHo+ifjn0ljvO0GVVWC1UBgw8fM7AblZhQ6OO6rSF
9pVjtNMROGlGFocax81kHJ0Mlkp70c6sFTt8HZRKK/WIwmVoClHJpgTHqyQaL5Zh3UFeX2+A2DxY
buUc8bJ7nB0aHfnxY8aH5yJiSTVMTjecL9LAnznSX81PeN/vl9+HP6BIzoGMIjaNT2z9VZ+pFGRd
mInd9zymtLX4WzUWx0c9aNaXZjWB6PuRS55R+FiGIcHmVsMQpL7eLsVNBvHiuQGZtOs7RK4p7kYI
bcOIspj+k/GxS75Y2Wyu2bK456bCK68drCt9NnOPCit3wiWgH6zFBa0J2W25vkROHbjuKT/RcrTG
a17iIMRaXU1xbuzf/V+p3LFy732Q1+SvWj0td5gF4j8097rPY65MGkvtI+khXNdlgLuVkPwFxgx9
5Opc8jhM8pPd0rlfMrWUhNnS6DFz08mTLehCI/75ztK20tQ82ZyQSC+vfA4e5jkx8GtwD27sgAfm
RQS9BkZx8RA7eQokIiaV6NWYNa3WcxafHCHDJ3a1T8E2nijtDKzGeUMIRHGJnso1UqKYbsu4aE/e
d8uUzCbnv7ZBpv5hPQ6LdTMOmGDtqxCtHsO0Cx61zgafj3DB4OvTcX+xFH6KPOa0yC42rQSXWZXb
WZnMlTwjolWQvUceW8PCnyhyIYs8dr0r22lkPUBABOK49h1oRnCOTHc4EoP/XMBYHAM91zGtIdjw
HdFOWwOTyQNPlAuuc4KE779sG0JI+3XQy0FrtJfPzIJJoY/m6ZqSCIiaOpgrZMlzljwQgNZPk782
0SxCfzMKhA8iHszGPfJEd5hSOTY8l5qe2lZxML/J/gi9MeuA3oOQyuxqGXn3VOuX6Q+1ajc3OJL0
BbG3RbMl2f1k5a8nAi9skWJsAREUkXaG0DALH72SScxk+aCdfKSs8IVNEtvm9juwYwVBzZEYocO6
aPlBtvNX1gacWBKyFWQ0otzw3gDZYt5D0IP9ukIxelKN9kRW8wju+Hu9gUETZHOzyviz0ws35U/i
Iea1bHaQ5etgt+TZgEqd0r9/HhQmkFxgbWYp3bjqJVVdBwnBa5c/wA2nCUEfTo8GCzbTy6YSLMgo
o18TXK69AU1rWR/OROAc3AYj4PzBalQOEYHVuhJ3dV6qQhbZfcb86ETeKC2h7ULb2PdIsc7yj/lm
Imxky029GhA63EhzZrE6kKYsSlfTWRfE0iWSgFPev3CF0qF7wJHD4Nf34I4XypVSnc+ljBx/VqYn
grDiUTrYk14MUdTO61z1CMiNTuf3UWANhMY3Hjk7uVCyXOoJP+H0E0t76T2K/8D/47y90TsNQR4O
M9Yli5SEqRQTIy4BkDsLlQTSzT8JhbAy7AuwgVvhkpxwYh16aHii7RonwA3i+vNNi6WX31q5XP0j
u2xldRd/T0DznJ7lvcb7KqHIrWsSZ0Wz+0rLvWTB2ox97+327pJgvVxDYmJMshs06hGHezUVs6yX
sLW8MhLN5gORdhkXUYLzPbMoUUQy49/frWl0R4u01IT+UtbrR+lKIEg+lE8SdwhFugHDu2kr2y7q
KD5zuO7MoCLyZTyCOcx7jDgc2sYeI5PFaoOJchfe8ry3pS/XIVmyQHClneO7rjb6JIywf4Oqw/wh
SYmu21azbYpfcXBLWLJtZOMdzQ5BDiOmbD1GfVF00Btzs8Hozf4nk9ljCYZFJTWKYETk4rnvNVvG
VTzslOTgIK2r6pMFNPqMJ9nuXzUdVBY9ZkXP6veAt7W/uEOeag+3QsQgkaR2kYQYF6Sxjd4ts2jD
Rdj0KIoz8FZITmYrQVChP3Nxvh+FVUIIc47ij6vENphbcNrEIej1eVyVxRZ0GXYsOW0XnWiU4hsR
/sLvntmUuP650Yg5R6kGsiIfkhjwR3x6Po//53eR+0yIiFWtbefMY8EB2b40nmN0I6crh4tBgoD1
ywfRrllV2iknGXgGK4LPEcLJ5maDsNF1N+vSFM+v7+C5v0AaeaLjwXRI20TOkYTBW1q/ytVXkybu
xp5eiTCES8l+Fh5F4jlP8PPz3BRK40euLXzRKMwt4wacaqV4Eh3aM/bEamH/cSSoGtJOfgT4GAQL
dKH4La2HF1BiKB+26K5Pj/fZ3tGdIbOA1tCnF6xMkBXdOdG2WeLhNswjV/WFAxI0gwhi8EvL4MZv
uyeY6zsUWbZDUBHChZ9WCdZ6ZAp6Jz1ZhbHQ2XBEtY+5Nqar8cJ7VNBq7rrvgR5S6QIXjSAogXvv
Q4S2Zaab0aMlZudLZTcAQTiuIn0u7Zx1xZoS4q2KRqOiu0V3rAFq1P3Jho4sB9MHNYJIYs7ZtVcB
4O/f+pdziPuJ9DkFcM8/Hqsgem7Y2Q3g+1YdVLakiUxVES6NqtpCy7gICYbiOo4XlsfQPLXYRGaS
oksLV/D80s3/LtXgWsvzhUG11RIWzcQSEGCEkIXeCw1VyD0jPkQ2sRZ10Lk0Tz74OMfEmR1t4u9h
a+E62eDjqG9E1bk99UiLC4vyHKOQWYjsIG1QokDRwighTZeJUu/MjQMtKkDwCMbTgn/TDJ6mWEbS
waDGRnbQ3dPQGP0uEdjc/FOWp1oF2oYA4JM9iOm5wmsEnoGoJdhp/U2W7xL59+fO0ESxb1Kf+PTD
lmI35s/k+cxt5aTzmuudToH5+0SRuNC7NbRL9WIdJxICOfWN0OekXoiGnl53A+VhfkJmW49BTdmY
S5jstOWMlGjEhQCag3G9n+lH0yWnDXamjorrPPcIi40hBq61QbE1N+g3mujZsW3Rq2HAZH03jKdj
PzcCHpYT1pzhy9IXJH3v3jowehQyLXBKyJ+Klh1HB+QPWNRPpUuCZ+kaN5hkN+sjXLn1eI0OW73X
u1Nvf66Sfa3AmCfZHdmj4fr82e9PnKo+E2i8fTZFh+kj+s+9fNQIodriA6gnIT+vxkyFnVq/CQdl
Fg53vs95KdutGIx/nZNGQIYjGY5x///1aqqcggbTs7miX1AlDMBW3aRM4+zDEWKVEafzVys+2C5h
ui5f1A7wJ6M4lWQDh0kUmo7cK5vhXI6ONH+KmF5urT1Wotx5bwU/zlzDq3H5j5avyHVdd0Um72Zl
Y+SP6MuGxSwbqvTySs4FEBklcAnlkuznopeTlm7nZ1jujQB6RbsvRQhxkCVVxdftoXoZblt2eGbF
QA+7at1WjebzUcaQIXFKh77q7u7JRVK2HGbr/+mv0A2WnpKUWpfZPZ838NYU2MNymjGYhVxjuOnx
n2Yyyd7U3HkVF5bGz1QRqf4IyBpmIwZqnnTkXVFAehYSv1G0BPGLrQ4aXYSCSck5CxBFHprEZy//
gn+g7BOzYJYzjfQZGIoPR0xMKcY8jt+Bog36R1f/P9FPfVwgY1WzXvEyJ5vtjZctJ0n8zQR3wsVS
fQ4iv6xiicR2Mz9quhWeSKf1jdI1EFsaYyqzNZN04VTnSGPqbbnQjLEU7309zLu7ufNEr9+3CW1D
aK6L0Zlgflp+OU0Z1X/df+rnuCt62VVWKjsaHj3+bilO2cjdcP+I+8d+PSrFeeN+yNCyHaRZE3DY
NAHFVJ8c9w3DeBEZ6TcH+U/f1kyt9yBjQb6xfjf2LQa88KoLkvjUntY264ZUOT0kZorllVp49U5Z
8pXeUjMOxyK84MlmcdXY8RcimHAIOvq1NAG8U6RtG5REOq1jN9/b52+OiM8pVbOmFjJB3GqKDNMZ
FJqkC2yh0pUYjHOVzmxOW9pzCp5oaneVfeLRfHx6Kcgm8HYybJ6AYnF9eFUpF5vCJrGgtbXJZ0QU
5/Ct64Px38yQlOnn++FbeL0ZhFylQDGfIE5H3Ne/zxQnpJGL3uyH4P4sYAiqONn1QBXl0laVf0i1
8nnbPRrXqlpBkiSFTkLPdYgYc7bj7yy9dLWG/2g33Xcl9moMKkocC2Kh5HlT8sopb/ffU+IpsSil
VWgpdmNuJLdR5/fXOFZ2YwjwI1XV9Kw7X4SpJprnGvV2vRyTqyJJjMpeh+XT0MgDXPA+wzEr9snA
zqXfJ8arfJRzoiXyV0Dkw6B2tir1kE2Ni8CmLNhbOxY4NIEXIB4lj4MBIn5R6hJzP0wNR6PFDw2P
A9O7LFHK5GSGziBgLE7WXMjLH673ZeaXd/s9lUpBx6ifgRWM8re6nnocPgRQadERN0S/XAJsB3ya
1JCGMq3+dkGO6VXPIxN91pfgaruKjh88AavZNI4QPB8/0vjn2Z7X35VGVBgEo0s68ZhpBoFX2bOQ
EUQ8jeK88dsPWaGj8+TJXzGF2Oi35z1tD/5Y7S4Rv4TK3R4zq+DQ1eFMFE6aUsZ5hhp2XHaNkaQw
dHGFxg2iUVU4nTLol3eGbyHVtXQqHgeG23a53Iy1EOgYWWfnnQlYsc4IIM2qJiklLoIGKYKrSqoe
X8DhLztWHp4aKpwXZ+9cnfLLs9lvNozlfCFJNP2KapcJcCstOpn6WmHf9yQLRSX92jJCjALWOrQJ
LLziqTYErHzUd95FTBoOWZ/4Ex75Oka8OH0OcEiC9pRcYWIIPlT9I1X+WOQ+14QCYGbkb2tNlw70
d/TxQIrEr7KNpTCzeBjZqwDS55mt1BcXfTWsKg1KPDohJO1HrSfrb+mVkjCFqeXyM1t7Ng9JJRNg
3CuofvWqioGuZenmkgrVUvwxYVr9GPXNGuJ/bg4vQ4PW4elJkTuAvjBD6cU+DXXGr5HNnAuxDQsM
hfaRnhXLdwVrrSjPoOQ/L4H8C8szyd7oCrwWEK/62cxHssuhxwXAWe442LEwBC1z55Ghib/Hj0Te
2dgE2qwByO3ZHZO04SmVuNWU6744ve4A/2HDmOt/vERkPdq40Vn2FmeQTFd04Ib3nKr5bCRUF6Xi
qsXa9kIR2SUwFEIucB3dskd2d9jptLnFQ9qKT5mtFjciPRCEnojUjlwO80OpdySSUGwE7ESogxCq
DWqFsJ7UxGEjUxDUggtzBnhNJaXyJgeosIphh1XzRisYSKtfR/7hbII04vG7bnH/rG2Eqsj10F1p
RQmw2L1P0e2KZmnbp6H5Jx1HdL+zGsJP53Zp25DA3hLp1gMOZPmbO8fL39XautjemUErQqAtpL5T
z8//lmCI3za3uSmk88KCEmwbFh2zkQ6DXN9/rm5P8zhNwpWw7jpPY4RfuouCAo2//PEdIZtxxA1m
JRI1C1h1sufm2bI8/nh5BpaQRKGTFhLmKHKRAAwFKsAsiDGhWNkkb74v3zEjoJcoXTsTZhWBcd0I
KLZEilnWd3e5smjzZlKJ4LrH9PnBEHBSttMGjVB7W76nYIIsLHFTN1pTlDZpO/uuCTUo+fIKhmb9
SJzVldJLZ2va9XeNRii938FQV7t5vFDpKlYgYIcuqP4pDV+2SzXy9JMsITIhVRTgpHjywYWDYtYX
z/OZv4MTNbFEHppy86C4FpoNdfo3xeIL9NNJxUSQdt++QGgnacUJOFoAECmxwfHeURs+5ln2cD+z
OViYXtyKAY6xWIhRI1T4CDYHDYYvcAJUWO3QJehftdkA006pOzShrP8aIbS3svbe+gAcM5PffAV1
qNWC3KraDKJnGvL73ONmU5+c9bnVneLCkBiMWI0hx15rkrAiYxvAWozbkJnME2SbX7/GCtrc+38o
H9PwVah36+ANjBoGeTXOZJiWOgoGfD2weMdBMfKqmIBC+iK/ZXGWSuA1SjUdDrflrLdtxr7vGfqY
QcdSRjOm6y80QwMEus6EnOCeGUroUTGtVl2ERyuYJnSBvEloDQ0VnjblnJxggE/nBOZqwKUQfA8p
eRRQ6pzN4QLXMDe5rX4tNHKG4D0LI25Q2w+LIthqScIrnRfuZMhDl4ZfaSlCUNnYKyVQJUxg8ZR7
GH2kS/GCw+lzJ2MpfcIn0N75A6xB40zjZGla0zWHO1Imm8s6E6V2vB19jnFSWsIVoUgIq9UkNWbd
a5wVjaI5HxPRgqURrJfUdubrIHCadwTg4hDGk/uSLZ3V62M5OWzu6fxXvGmxpWdghw6nbhS0ahwm
rozs5y0Ha38SPwJ7FrwptI2ovxYmTpNi8aEMaoq+4nrQ0pSxbWlqOD0FBYpFuBaPlighoPO5L9pB
t2ei0Wx4VsWKmweonwDClZwF2RG9GpTIT1VP1NW+jo/CsEqmeMXUEmI/aPJwH8dR21YSzfcFje75
LspgcWYFKtW4qTcKdDu3vMW1L9tYGUK+/gWtfhznOJNjcxywT39lW7aRswPfp9gtkeLEEPNx9kOy
c2+abqSr/4Yy1G/+FTq/1VXWHAL+5BDO86afj2ohr0b/7RSN1a8vK616EDXVAZ6nfi4vXjt96udB
HTPW8mvxA915tsv1FdsPCCcyZKGMEW2RU1z9zUukfnfwRtX/VBFKQtWquigd+yQHkQXsuOjqjHNK
L9BOfu/E/lUYEebNJlUzLR+dC7YABSjc7DKU5ssr02Qe0YksJnJzBWreNlHlXLVqYnDykl7B3+dM
feeIRmf/zMzG7DDxYFPbeIH7+/RY5waiy3gNmEjCIJekIDp9ptPK1Rd/Gg2wvGiwsKhIpRiyx5fM
gx+pY2su//kyUwnPhFW/tlzEoc3jxmVOZ2SEoiPZwY3qnLF/aM0jhhPtRpH13dIdcxgeAVDaxGp/
YR910LpH9iT1QkOvoU0PC8g68fdtO3ewCn2Bmm6zXX7V1Icc17Cei4QMUr3IPRE8Fb4R0k9SCpse
XAgm4rMsgyp/nzdWTc7vuFGQJfJ0ZyUj4WukcNpKYz8J9bRcQp/o3v7GeFN6NbogjpTGtLujsKbi
hNgt4I1TX8e2rAKWlRaCY3K6UxdNIEMd21QSFZqO9sEZK/p8oEkqVxhSwC4JiYhnyupCU5vli59p
ueOTCEcdF0AKT2pzzgmnak/xH1p/aQfKvX+5w2WxTao3RX79J/ZLOB8HNzSGtJ3IzFxwnfReXpBc
6kQvAVEBUFsDJZ+HhWrkeLq6rVMhti8xNZeek7RifDp6p+oSnXE5Bjx32hO2AqOPdslqxpUZ7db+
a1hYPGlz9Q5YqqdvrkHoiQGrj8X4wZ0tXA92WyflBZxow1v6bWfvbIZGkCx1iod501eOncKNuEWi
iTpMpSm5u977bm6h41Dg2u8EWfbeAxWmHFUk8vGyVqRJV1dPlKhFa+2ipw6jzSxn8mxE5fdTQFOu
r3l/smMaUU1uujQcDclIyBOQX/JyMyJlYYlSzSSPaKi+h6jtgPPHWKRsrRtGggImUL25rbnCSJD6
qjUiYuO8KDNplfwRHIiuEJeZSKJ/e4hJTDbUO16La+lwCdH8voeEQSuDBdqb8juCNFlnFLUK/gOK
Vu2q/P3jvLsYr/BvT3yVwXRzBOirXCcgJExX+QaU9xAEta5+xknFT8yT0V74HVbLtt+XOnp/tX6J
rXR1Ba/Zukalov9+qQvCP27aDF4of0KHq0a/It1ggd7kABjIuF8Lpqo2+mKds4+Toa1KSYLzn+MP
ck0cTBSSfAxzwzewj82rgab2uFucvPsWUEWQa9xvuZx09FVO72eo2ea3G4HdwyhNFXDfoo6Qc7Nk
vLGdB1ihg02LWh1iDrANKiycsEnJXPsM0dJLl1Cmo1Y6eO007PLk7hnsYB5RvuynrLS1ii0GphGg
ZOqwBtRgTe+qi6MbASwnERA7cvZ8QcALpbcUmrelwr8b2FxJWjxdz1HJ4F2kFtqTFZzM83hBaQD3
su8KK2+OfC5bF6CvZwTICq9cCH6GnobF4SVaGXX8GCO0HUZug3uFjlX9UM4Hx3myiASDJ9chYpVf
rh0mPEtmOOyDKe9IkdzA95frrAJvt6wSwHP0cqgEIzKmeXcFiILsqY4ZVoF1235eOr0+m72ElmQD
UcpkWUxNCz4QhF0xgqeUWoF9c4ErCOgPd75DxHO1cqZPW9km2gFSJNBWgeQ7olJBuz6rSmMl3DzO
zYrnuGedVv9e6Byk1QmjDX1njMm8h/4/+jQ1ZM30DvcLII3wd/f+Oe3OekhwoVb1eZY4SLiHn3Rc
JU5xgLmbH6+MJY7pdcHe7VpaJZeSeWqHW4l7X5RDoFjWuKrOna3meh3FgZ3xHjaElaNQ/vmvl2N3
ya55xTwFoGwyP78egq8UJLtfIspvLyl/6X8yJuWYdc3VckGE7YZl8mySdIOaxwy0rrUIwYBCwGRL
hy7Qc85G2hF2bXgM026SWoHgx4FRdwvuY0T/pmfAcAbsRxC5wX1Na8urTBQcjcXo18EiEAO5LCGM
SbQqSx9dDQVNdHB7asTLP9/+L0wU8MDCRlAsQkzv88ctp9v12pMfNM1pMemUjeyNNDKrtlKYrBy6
UvfH96Tgcx/CTgi2na3N2P5S9VilW89SkR1d/tPUrsTmwGDchycRue+laQXZIpcIukKIR5at/8oZ
nWOW+eLBOk1LOTCd3Dvz51IzddXH0KMaKUXog/CvCEKMQY2GeLhtL2EPiLCSBlnTmkxARZWllPsB
Kf3j0A1Ouw51xTMirsA+LDptHPp6kLu6Kp8UIxUKkqbXb0Mf5OJm6cCZUPXCUFqEjuejuTw+DUIz
9+QxcLvhlELc/6fOgRKqiMMm+c5lHc2kln3v+MnKeTV4ecii5KVgf+/76HYboz5awPRYcYhxeYix
9yMCkZp4AMf2AZzWcuH/kQmpG490RiSVq4zNIl9CWb4UrDDVSE7MkGwm49G/7ecugEjJN9wS1VFg
ZLZrOadP9vrwQ4YKlc0EqFP0WPt5Y4RCB2uVhHvX0o/RHlVEMaR1JmIbLBcdjUq/9AXH2TAnpykB
MjxSevewF2iBcEIUy37aEEQ+BGtnzkDeukMhRzDM6zV1Znkfix9DhqHzd/bzdme6ubrJ3v7BwNXH
Vuj8S9x841Fl5HF6erQg4MfbKvmFkXtVhcQuF3PJ4tG5zZXjBSB+3ZaSqMsAanQ3bQppPGjQGUbU
+bdNIz7SluZWvC9tx8ehUKkOKcBac3ysHL2wk64CsCXspd8swVne13przaNfo9b/dZERxLzZ8Hlj
7DEoLl2SbtAPkW29UJH9Dg4bAOkJPIslQ8DtE0QnHFb24dkxb1EmGbbwKqr0WgxtVTJhZuBiHf8S
1fCws8+/YhqoC8yTGN9elasMK1tOYxNdYzLG/HArVdWeJEvR50brjag1wr5o5dT/WqdhdJ8P/a6N
WeVIt/11KB5i5d/iyTC961MzoiD4OtXthZyGj0bqR8VLNklbi/yrhGMutvrkEu48G5ScyEkwRDhF
zA0eP0gAWk4ZukTSetMvOh9JQ1RhOfQf0Hr2c03texg55oi4LYQh6yA/boWXhlji+7Wo1AVvZcf8
bWFL0mR8SbSmgoDHSDeFz8cKyoXJfv5SlxAyExVp1vwEwxstsPIIOa3TJAb3jOhhLoMOos8MnCMT
uHNCrRPxxFi1CZAs8B9AHUKLCZ19kHGQCXwa7a9BeW+Khbj4wWcTLdluSqXrCSyR8sK9pzBncOyI
4XXDyt0bX1n2sgIuftfizciFFZGUnlukRcRP7bfXKktPL4NemBrNRKgB1vmE+pCKNu58K+YmbfwQ
KcjF7eoxEgOhiMCaB3+L4sZjVaLy47NkmkiWcLS8cVGrK9qBVqBX8T6FRjIQMNIwmiZbBR9CAWcy
gZ2/j8RqyYVgVECrbarz3LI++/MBy40jlmfYRuBDyC+TFzsc0mkdeGLnMdWhwv9qOXzq/ayfNH87
QOonFZd/U2moAc8pSc/uoz54o+d5zxfqZ6mT/qn2oR3TD30wYw3p0I3gNqsn108DdPfvJJa5OUhh
7FE6moYaqUx+PZheDUco7G8kChlb5gJ8eYGCU18rq65NjyDtAxSMoib/jaLnPS4hQZplKm66I/S+
3WZ4qa+mfp0QXmjaQng7yGKG/Pup6Im/oYO/yHRpfJd2kHsLzeyVI43OYXePTw52fZXrn8qtguRx
tfGwg9MSdRWP74tPDt2yVtza8h6uL0RaWmXhmHG85VSK6/JLPZtot/b/iEYJTp4OaBJTE2D2jxS5
zVtKP16g1ZMmFD0YtwkEHQGudcgIZ3QHJhfHsvTyrDCjaDZUVetn8Xzhgsw4IU7uP7rTy89643av
g9fs7ifmzkCEpCZ3CNI1IAMkzrAdzonVrKcIh9S3fpKG6zziaqggvyyKcHHRzafPdWlUI/Zvgno1
Z38JHCFBSf4oiD7cTc6bBf01ITXpKlJCmJOIeQMfDQk5ARriEC8RKPjD9tM8fuP5dBCep44ogycQ
OTdq5PFMiTRk9syDNSIP3FOrKAp9r26ILUe3nX0O0Lb5Y44j+yC3jcKGov2Ji4Uf+nRgNns/tSGx
sAg8mdl9LYA5wYhtcW+hOzxBpqho3jjNwprukxkDVj9Toi2SftzmAFGoWOYZl+YuaFlY+lqtXqZr
ubibmCaHRb5tgeEnS9A7hQKjYY513FgBgbopTJSJ438h9Acih7fhf0MD0/BJhEtOxl/6XSosNgAz
UQ11dQaqAUnaiJ/Hz9KPMnbmiJx83rb7H42KDSgSBPaBZqFsNrfsADg5Nm3Li97tI3qc4eJI2woU
3Ble+cnUrtrkJJi7zbJoW7TvhB7tlugDcD/3QZLXGLobOhTZP1OaOeHjtaiixlMz7DcZmZihGX3z
Xa5F7RfPCfQwEMX269maX/eSmML3GMuTXiz5igAAjI25G2Ht7noH0s8DTHWFhMWn1JJ0LifaFFO/
8JT7vXYBB1TS8bqoS3RnkcS8G6Is3mvNQs1okoJrBrXGAHxbdvL27y16boILZfyp/Lv0PaicV+NT
TiMeWB5WOQfByUs9CsfYIEgEYVWq419ZtC9JNO8o+osvyn/g7JHe2ZalwDXXcD4B7GOeaHXd7iz/
56lNTJJRJgNd9aSOqNC3zNwSjQ29nijSWwl+9Id2vpa/Uw0AqEyUuMZcaTOAlj7pJ6aQlT1hTY4/
9j7JATI+aYrqvUBfmr9knnY2t3Mr2Lx0Ts3+iQSPWuvWMxBq7+DnQH01A02LfJQOF0zSSDfB1oIX
pPbJQSxmlV/eG0upt3+8HuTkUdXSqgPF46sF3nTE3RKXSt9kVUPia4h8Wbgbzg0avHLZY1+fHsfO
/HaTCNS4TNkJmwBbZKLYlB5Hdp8D8v7J1J+5DonQWlrYvKyQZcEEZrwJccWTIJWKWkNegd85u/bl
ExmZzgpg2+xvIs5ihCvPu5S4m2OzAuEpasnehhGp7zpRB+E1TQZ+Aoj6a4rX6RkWCxKEG8lTQqpm
whI/bwnR77EJiM9rIenMgVbDAMVaRPMywfe30h3+si2LuRbBK3dyuVU+oCY66RjKLV3LRMy1wGFs
zuiTcjVacIAYaOTS31EKGhOmdDZCpwdvZHFN2W55Ueu674MCB4a6+ntdj4dbBZakO98hQ6xk1pB2
25SYcpecTKHPXEOlK7iYjVFFA2kBH8YqvkacHEA3NiD8LmIfQIlToeYBez2YYHtKpBceSNA0Jif2
A5SeIWLRkIr/FbVpYdxdMDGJAHPQlQ1ju16OytmHS1q6RTDX3QGIShrzP9E20Oz9KELO4LJJuu6G
OuOLktPrGQm/er792PkcMr4ZD6mrz8jeWyCn2jZEWiNvDZ89CdpFXXxTmVPpEjfl7giRAGh4fncn
ls1UF/7hOip9KnCEHTPND4M1bko85BqosogZQ9Z4HVofbFR8RSyX97SvR5XghS4AQN2m6Tid9oYu
tHLUEdw5km1/su+Z0eeNDrk7GxmWViMGOON0sJ5BMhusoAzBUfY+0GNHvAd7p30aj7oNCEMYfOQE
wxV+Gbuqv8qpNfMi8ADxko8aVnFs1E/dbUX4PrF/+zZuKrCGnr1Y1z23AtYXCLibZGlpIg4TtYVU
1xWmj3qSnGNZLYzNOXE5W5FiKD4HwPDNPU4XTyTTD5UUp4Ja6TWecgqCA2LpPmLtaO0TFeOL6Tss
ASgyNr7i94Wk6XlZtW/0INllVHgAMgDenS/nJDQN/9CdfgGDpzAaCwkT6mId+TybPY7SZq0zRLwQ
GtD9SDtdjmrkqrwQS9gKZh+DTKuXWo+BGOieHkEr/y+rP8aQiKHAZZcQJDWJi6Bcdwk/nN/kpOE4
LkTOfQV8vATtLrosiRG/8f4V8McQn895ch9o2pOJ1zhH7CqksKbfUoi2IjsLnNKZA2Kpb7e2ifmm
+LX68SGD/EG4/kS8+nf7kGUs7S07KTtNvCQCdD1kmtyC+QYwGP7k6fxMYP5OGkxQXsJlvFhJwrwP
jBBs9xposdRP7H0zXdrUhmB42tTy84PY4groeRb7BwvS7UMJrrsYJQATpaOZjeh/TT4znf5Tjc8n
RwmOyVL3xgwTH1J3Ap0oRz6lyLJ92m8f3yzgqzo+E4twNoOhaFF8TpLhFlZqG5y1RSqc2DZ8mIb7
FjWUhbSZYxKWZu9qHOMOsBj5btm/mYwnM1aVFdQ/I9cieLg7ERXtfeaRsWCNwdsacCfIronX5Acw
pkuhJsJ8P9p4nqdQJ0oNHCG4cpfHjw2/Z0l3qjJOc+NB47UHbGXSIL/EOQtoX03wtJFSSG5GwlaR
jJ7gPdMEjTyCIfbr3AI8nJRgtv/ZIAgZaC3AHhzYKJsJwwWFqSyMm8kWDtibynMjcW+JiHq+5MLl
gqodcQ76gmyEwWj+tIB7j38t2OmZIaqzc5KxXO1Gs4J808qxElSkSq32pOuIoRdjHSCs0xHjPu7m
o2gsyS0hqw2i6sCL+gqWEoHwwOJihCp0Ch8+ifp1tDbRmq4FRGudhhskSFatxKCW1FgqPPvDWc9d
zwwLVVsONvel5L89Nn2lDm+Hc1dSbShRUFiFvAeW3YcqhwGDObgrrpKr2x0bwEsc+yDMbvlbDGHG
e3QBd+YNeTPUxFMoxpwKg66OBbQ5SX53VCwAgd7kqdJcW7sc1wVDdjPKfIaCk0gq1vPYH/gqLTDj
tTtZethl592bWIYCQryC/XKhpHpu29VtCQCDNjwMsP5dwEvlncvu3jwYuz3GShZfSus+osfQafk7
tSvZvdQmMy9ey0o5cFjzmtWRVG9ph+OXukJHDpEu7sZlwfVUEptp86816DrdDVBsN7H6/5SxF/6y
C6jArbs5B1Jt9EI19elvt/KLhCW3YYm8hU7BgVnKznzbTDxcAx8P4l1u4SvBHEwHrtGdY0IrMnK4
X6GgiakBJr9cu4P3s4FMnzRbf6mOn9vQYS/1D+HBv9jS9zj9q/W0LvTQkELr2mOt8godTm962iU+
QLGu4JvkM8BvxPsL5gPrJnWjKUY5QgMTDVhUoITpYt9BNw38uzMnNaB0ShBfB+NCwMB87s5Mbqq4
U3cb0fK8brI84J8Lf9qo+WFAUINdhH9crpiWXypoAxwNaL7vjN7X0jCLlfGSE5fiB9ms6eXAsf2r
Lr2bP6WuWz5yVoYzWtQRa2Bn5XRhBbL0QojA4J1apwEd9uB5ZoG0XSZxKK7M+YBp55wnXTg581E1
pLmT/gtd0CEtT/j3T2jCaHcUYizQPDZFzt3+Z9P2IWXcxqo0gw139Bfr3SoO9ZTSsUENS5Ojv2x1
7mtZa9INFXlnV6DAFThMVcr2xaYUq5kSK89NnPwsm68uuYxXsfK0p46zB3DRxYabRC3RrI48vfIj
JotIHY0/1OrUVcqXFQHox1//Cshbnpjex5oeM1ebt5JnEr7qBmB7mD5M4Z2sQr6TbEd8w01uvwX2
xznPqtUwpKiHt0a4U9C4GYn+NWozh8KrD/SU+sbZo08k2IIcbpqx/O/ej4/XQb63SJvGHX2jDBHO
SfohyvdIE/iogEIREgB0zc53jMWEf9vMXdMDL6A8wgbTI2YltDcR7WLoRsb4vKn3bCr6vT6yAkJQ
3Ia+A1iZamxUNM/A+7woFLVlAO2u4+k8KaHo3/eTbIJXRDxQe2aNxOEZDRGzO62GLFUZ9DnIRIuH
Z1ym39JKI+MGCXWpkADILqNZ4xFNGBCdCoUDmk1LHHVIJFIMEuTjhyPOs+xZ32COfugZJ3Qxst37
SL3lNjWSFFA+mS/yrWcAsTvgIUaYcwqUcsWeBpmC7QrIIu/guLWIR7ppI17ZNMAzM/En1y/9oCwK
TF0hbwIpTzjhooKPWEvt2SqtpS1DmN++RsOpJIaLnKDXynhn4j8atpNvEJnuEiozqRBnAOP29FWR
HsftJK1svG8BjZjf/dak0hpiY3VaKFeRf2bY9txyBpuAG8s1ltGTt7mVY+JQt/zLQbZBb2T8nnuQ
WA+P0IMjq+7QDFgb37Ut73LaPLyg6mce6apqy+6G7LkDD0/nS4bwxnUVWmKgVRlTYQgaI5xjRCgG
rYfYe6NgrOHkugx7WCvx4/VSrW6B9BKolfgRpA4IQXEqncbJsJpIOJ54rhQ5rK8wkrhrMq7ezcnn
LG7pkv6CnbMq/9mTS2JYZMpFoJhU6YyqCIfKlYAZyNUqjylv3b3snv8c4QRNkGVgKvfLRsmah5j/
wmR/Kaf5+gUHuDOtf7LeQSl0FiNNHohy78Be2fc3xzh6O/cl/mdSyX97/hGSNP9t2nZriBPQArqI
0miKQY6/vcAmJ6HOJ2PQboGNQiCgMAsa9jReFIzUfSx+n0EAYT/RN51icneVrYW87ZuvGaDCwwgP
qcCtMSSMSa/FTeelBe3EkHVElLeKHxDzybwJBo+QRw6Wb9Np85vSC3KOIUKP00RdbXURtzYKhckL
IzNHcuipV8pxjrKqOQlYIEuVSblbOlpl75Mjp0apZ/ARFlIZsVVygLcDYdoX4KPUmVE51QoTojUy
hrk4rGkNYbueaplHLEYU+Wdo0KqmIEk/XrDf8+bB4F7xxW/a+uoCfE4MSoBPB78MD8P9XSB4b+3m
KWskDw5makQkmB4p9z8yDxzgpa00WSRt4xJ4DsU7dZc/B4LVesRhNeZQ+jxn3xZWMOei/1960kUr
1BP5ewgUM3myqyPmm/cLUrEO8fJBTmdprY76v4MCaLxjS5fR+gIitPrWV6TxFHgMTlXUAj9EoQD0
3DgYqUzFNuO5+ovfITBhc0gCMrtRQOHrJd6HYkbqq/qR4KkfOfFWjbGBhda4/b7LIQpBGrbdef0f
jndntVF5ISfsR8N2srdGlMgT3RPBLBgeESk9rM7EgEdPp3YS8gEJMnmeaG6MDcUaOk4eodaULmM0
OkaoRawJlaAmj5F7YrsV3AfWzp+VX0CNF+JFIiNFGzTaQtReJ+IDAiAzrSO7rL2u6ecw6rfu6c47
JX7f+3aEoV4M/JAvEPqRdu6mt19EPKvz9d0SXb7Szzg5sJu8ULIGUwCrjzn1jfNlLe0byXapcZzi
LoEgTy/BkHNAmgOHRwMymzyNMFXiZyMq7WnNHZAnOsP0FquYMdvrvv9ok0A4WEmZVJ3rFVw4RNAA
xlW0TOnBMzyfzyC6pUDPPoyrSjcMwE+YAG7+Y/d06TH33LgAsil0X4IbBsVb9LjapmsL+gd6tfHM
i+gfefJ1NA8Ktl7XNuPsk+tjcEUBLU+WV1uLiF68vlW4uMNqrKOM0CQ6bLz7Xb0ejLvsNBzboJZC
LqwhBDtvGLFcmtjdbVj2Q6C9PvDegvJM/7IHM0Jxb+5NyS16lQ2l62Dz1U6PpcbOJnWHzNb5sNdz
JnG/tFOZNiexfqJRnllAilp1v7Ob/cFR0h7ekkZZJbyxS6CmFqfjVzMZQwaglwpf3SJltmyxB/yh
5zWKn8h0LuBCzbNpMD9Ah3matDcBjtdfNKfzrsRNWBnE2BxXpPRCAs0nmKolQR1cowt3P69WJJlU
RStXdsA8hmlUgaoOhAYDjKjTRA2kmx8X+9kYp+xf/6AfT1Cb9ltsrKa3v6rvwljQjBZO6oFXsSzb
PNYe9nCsCJzOETDtNccxrnLAXI3yo5yMQUqEfKvZltrLKyasq3MPJtqPZQQXy/ydvW+ObHlfhXRl
PdpYIWguVjKmUHrhzMUCv30vMlOkVo0LLU98T5JGBISnqJT0/L8mfLQNFs620+beOxPi7VnUjm2z
3YzOVjz/m9lGZkikOrwJC36PyHxYl3Z8aWitjdZsCSzGMH6UzOGNGxy9PnF9R7PH4XP1S/h593D1
7bgF2Kua78SWN3fAcK6nTV3qXXZnAhwpj8GjXlHnFTgb6ZQ0JdZdcmYLmt1TyU6fEbkGfqIvM075
RhBSwO2TnjeqgRIy80QX+RkIxBTIPBusJdVMBlUhzvIfKOGca8VNX7G/RnCgIYaaOfPA42AcL4Ed
/kPxZlE1OtMPF2stBaFFtaOJAfe35XR6uTgACg11eWOKP3vKSS/e2oKzRRhlWUGxELLIgUDArhci
0WQGAIfDdZkRKnb84GCz9V9Pk0KU6jcAy+9DdO9NcA6Iuq+vbE4b5gwnra6VPZm8FPNEp36M5fqB
OMGPCNSTrYDmkziWDeK/E+ccK06/Ka8KWR09KQuKk0W2gBDNMMO5Ke4wFT4lLHB3J7D1wMWO6MfV
m9M9N1D4eCRd25vuGyRLZq2Xye0Ng4anzfgmKMpZxAcvJE5oTsyHWq+x6SyWr9vhbuxdnCDaEaCR
UNMTgTjtwIk7Nq9JOArC/mqHFM1r34lyblbMHGtETowoIEdCnxbIwGhu8hErc4Saq1DaP2VtxhCP
ROMUKtMuXg+xGuoYWlhw+aTARVLt+wXdeJ+yPPtpeCrA/OUXs/GEzqlrZOYVqfv/MFaThq3bamnJ
EXmddaMCGz91edCrwL+SZip8qXg2qGb1AL2DkjCQEr/qQtace2ZGvtepJzrb+bKm3d81ZitSomlE
SgC8KENS6w43bxHs2FE6SQQeBkoYKIUmiWFzGffXvKFzHT+qSNkMicL4xkZuCYBuw0zXAXBXs/NW
EZ6+bOUIveCneJQXgeVujfU3wU9AQDbMOwOv85hVqSQTicE/I/jBbaq+R5LmGmFo9M849YVUt6zL
8sRbYxi2joJv+UEu8J+LmW45rL7qTe+T4ZnKbHTghAvB46272G1pubuSifwC/sTDspnWo9/cOi4w
ehQA8JeFY1iYjSxkoRYgvPNJpl3YsCSzJymmcF11FPZozP4LRLXGgsCfxxHjTdlP+M9vyZIZT1uJ
/+kySEDTJwp5NHMBVvE5CxSFqx3MjnM8ylvN66OlK4rRgrydzg6GlPCTND2hjzfAHcs5sX5EfshZ
TA9USfu00w7dxqFOo32Q0SDK8OzhVGlthKkAVkldEDbOXkBEpLMG43hhig1Y7r55aOuKdDU9FPVf
hXJfwSmtxhSaUyvJ1w2mxUVCgd0Ne9b0jDK2IMzx20fIhwZJn/fDq3haBfrGbyafyzNtZSPKdIFW
BMlgpd9u1KrLPcpSBIU8PzDj/+p/wGCu6r7bD/+WgiEWYd7cxpnV2ycLuCSmua2Fp5IY69ztxDW+
lU38XU3x8QtAcImZ0lKX2NX1kxTUPnfmBlU1IPhsXojgh1YFw1Ll5QkkB98PawNVJKffhPKhKGOF
4SPxuju4kioQ4+WvCY+NxgVzUF/1l+Bp+ORW/XdICqT+4p2I+mcpbuXAvs+vuwmQtjcvfZrV6vAg
DBPyN5x/Sf73errIg/mJcTTKd4K7qgxLgeKqzjoF+jzFTm/nDAEV/L0mzaDgygAi8tdtV3Ye7Gk0
a2bS+pR59w8CpDyLhFEwCSMKdBrvh8nweAdxCxw1HOrEx+AEINwf1jkpO9MLIvsTJ71EXuCyCyWD
pcmMbH0jaw+NEWazzQsBx1yR1wWTh/2mMTJxo7E6Iu0HGGg6yxuyxapIEWzYqpSl9Ng93FLp2lGL
XP2tYKN/Yz0NtDdXXDdBtTJwF315GLxkAy74YgLY2kD+rCJ5f5WDXIdc0u9+Y0Y8jDwCIv04cKFB
ATYNC+c2H0AL2oWH2Ia6RaIaMp6xSEgilJcaFF/Tebth7QGD97r47CTO8WLisgCZRGLAxEHXd9U7
sHktoXFLj34ClVV6L7E0OnI80GX3Vp0w2kWLR0899/FRwIOxuSyB4J5aYZIduVg6xoBxqH/BGdvr
1L2Jxd2xPUOfw/FCkiE6jyHUtvPWpP3SD1c1T6xtcDBhovOrsZnSaeAB0UFtiMbtGQhSiYHU1bKL
c4t+vf9aZoN3sMxUcdj78ATb9gKfpJh/rxgokAyI5mf2X9cpXM1LwjEYF2hZM4YGKzGmViEdMudM
aidABT3nTFqLVsPDCVA6As82hTTvZKjMjWoGdNmN/diNGCvx/M7gUeGje588bQtAXS5lPoMW+4ut
J8tumu+r+sVWJ4ZIcR24cBo0R0n1v24C42ycaUrp+Ta8WHV5khguS04YyJXJWJ4q2Alu599gQpV5
ot+g6+gEj9ggwcrSZhWMlxdN8DfaVb8TMed0KKr+ys/14vngmU9hneZympuKe2pRSk1khN0PZuWl
iDpN4D55uy4hWrEJ7fEybVks5+w3/BdScyqSTIpg1tun/qC1ExbpJn1MZy+Wspwea9NpydKe0VvC
BVf5ehtHzNQsQ5aQq3I8C2pklFFwR7TLM2tu83J8hiEpc0gG8ysgxZ8vosCtY7SL7IhyFBQdmMbW
phJV3BngycBir2BU5KNa1F7nVrqfICGmmPY9Djry3yWV1yqnm4T65zf/rvUS7Uf4wacwD5X+61+u
jTaHhIex6LpTysButm3MlwWC0bvKzQKht7xZCTLyXjVVaA0uZV5aNDNmZ5wFBAOVcoGTjitfW9zL
jDBFxTaH06S9FW45wb2yI2mzfnKY9Da+arX02vm3MACcUF1zB3LLRyiiDkuYn5aHnXECq2hlFdYq
aTR0xBQnUY3PeA0E/kpsW9PsfRTb0Saew7EJr2ps3gs3tidHKXNXBJ0fwUfok8csD6r6Wao1VDY8
lOsmDlLNGUbPSDcl4+z/QqZ3oswADwvFwThXuSVaGs2S7g9OG0p3NvdAjgPOVgmicwD/T2qnYrao
IRu0fAE/i4xY8G3wPAZIvvS59Xd/qU9/3f8R89G1rG4VMIhHGXT5rD8QzluIH0MCKDSIyLPj2LV5
xuvbVPeKp0/DkrQK4h3LwjvBB2VArfcrM+37qpzgKqa+AGFOPgmmvPu2nbbQT5MSn4edV+LEAv/Y
qaRcJLg4am52kG17FL9U9rIBsGgC9mL9tuYbtyY0dNQzf/dGhfVEZWO7giG23mojJh+JsY67zu8S
CktYD0I2NUth6saRLBY8U/ZfHOfJ1PV7zO48q7vg5u+VI1E6051Ku4yffEO2Py+pA61a34pG+gIU
oNBacO0cEo7nBC814WHqiuoiO+JjNh7Wbiul4AH98vgt47UTDZI/wawpjUXMNSOXLDzPdtCQv//4
66dT0y9fVPEPSYXlpJAHUflu6c0KYh2cUmi/eiqMm7Ovyhj55gxpD7u6vlgMT3OqZ1gnJWxqL4GC
TLjJy7cyfTr4kvNcYGMMVPmYUR6j3Wu8eMOZSe28wbPZobKkxwm3HaVj3Kqu1dW/lMiUEbTTNkiT
CqmvhRQYKj6++/zwa8jflw2zzSmk7fZRYF7parpT9IXICk3ezpjKDZzePZJlVgiz/VqzhJ083lvc
xYB9ugOPMe9M6jsTfgwwddTihl8EHaAE1wR2ynNILVO57OSmFcsuFlzu2m6j3mNYwsJb85kSmmlm
lRibVU5nnpFQATptw/KJ26Zz/yZcivRVds4MGDo6krV2Pm0i8DHCHpbaN1F9vw3ufHCQM3NEUZo5
cUoxth4leuaNru7EL7GFc2QeJZmst6laMbWM5w+9sYSM2iTZoyuMm/BjhiyXe8bO5pSV0dmWw0+X
XKkiu7KejemwQRsgeaKu18Kzmdwix01rzLZ5kuxCJ2IKnUJugmNi365rwNayb4HLkcITyfpF3Ym2
7Qg0e2ZSFvPV6KvQGOktSy3jpf8BSxXMy+I5QiINi4fhrQtJkgzt3tw9gRuMIbn4kys0C1oCt0jN
zEvvgeY8UKrDbnw3rbPgLefQ1puYe5vxhbM7cdXPA8ak6QaXJwTzUKe5t2EchbppiQcmRUWd39tL
u/ucLPmPKtdgNSnXIksmpG0YQAVSGy1VSGN0FY2NOGENVunqHLJQsF16E/JDVOJw8CknyaaxYYow
IFcLOf+LiPRcPV7h0zYNcvbFXwWah4sz4zX4wUzSrZLwOUliYnTtEGVp7/YEwwlwjgKe09yLOdaC
e5X9NRGlBpe9jwW+MFeYMF78fc71SzVkWhSfOupzE8G0rU1FrZi3Lhioko7TpAEIgaL2OpE/YsZY
qtU/Ea79cz0ZYAaccLtNwWAaDksZ7wnGzeh2GNb+HVELNALfV6LYfsbjXdCi9/gwZa4bOcsTwigr
krcJfQIAFzyOPSZuI5QxIfTmBFfRQNK5wAMJDdvCeiSpAkOzv7zKQ1SFKsXbSkTgzel+xciByI7/
QYuJtJFswffyzPHGHYbcaw2CQN3G4IWvRKkKaU2dXSAP7jDkLOaF9i69DgJDRr5fAhOLPD5F+Bi9
IMyf8DpGF5KEXsVkeQ6MqPBatz3qzPbx00VoyFXAW62GFyadGY7MSH7TzORs0yayC+edyuTDcfvc
f+p+l+jv0T20pGw+lSPZ4xVXLZZvLwnSeNzIVG9GbdN+UojZJTT4Zm+YC/ZpDy3LMk5ZoM9u4GGY
Ofq9Vwc/slQWlQPgcLZnwWW7UFEkBg9GUifygR4glBmW6odO/Ptl85aVYHyZ978TFcUyVr9oDhdY
T8WgRDKPl4HTaZQCn+J62G655fuvdNAyAsN2+s6UDuQi2RYADbWz4YphikZg7JIG8us3AW/gxKyq
ITXOYRpWjmfMdBolofNWProwcT7Wt5BVy0ImjUdS6ND0vyv//4amOiJPCMs/7fXQoPNqV6hIksmb
4psDwBfmlehaTcPqNb+j8EQutl6/BjYFTumB5NsNDcNs7ECCpYLtlQdZDCXyqUUHI/NpDAdq1C8d
EI4JUj2ZmffCPPepi388enmBPAB+5+ku/jRnCwYGv/++EM8U7KRegPnVF4eVsS4y2eM5K1rqIcam
CD4wsgD2NVma++mjEKUM2SWwCG1Mcg18tZgVrThtTllUbMyeVuCS5ZEc+Jhg5IIBYjeRIOpedHXl
RmK75URr1LFG+WwHXDqolBeBJ7vFb9G4EtCyHVT1rxrn6F0q27mX851N+vIiyGw9VXeGh8d+P6gG
9nYizFnWCcHP+0s8sKTl64Rb98uuVL1j0cja5oLX3yQzrCYT4IyO498zbtkzz772jocZy6L8NIqS
L7A6GxfbgnUWRY4MGrRS3iMyxiOWAGzEQ7p2sAyh0OWwWIL7D6u5NPkm1Zq1fRAthJM+MbPQnZuT
DdMSS6frHBH4iE5PRxQRKCMHAcAuwga+KYeTCNL0EVRCO4/u31SpnTjLscvenxYA9G9OPbOLfzlo
iv3FymCJ5p5g8icCTcieAfHIEAkLIMfLy2rPuLX2vLFEQEygF5MjyU2PAf/K0sFv94scxgzGf++L
Pj/loxj9eieB0Xc02O2UjNZuBZBiQkbgAEnEwxuk6PY3Y+gbeSMVTC8o7FzT7bTRupte8j6hPP8g
gQ8ivppYWpdtks8ty7T+TP/NIjqlFRJjw1FfEgCI23vUA7gAEDNZBEM/Y1l0770kLgmeR6tzez5o
F1ITSR9QZrunvmgpYdxMiYG98Wh6+L/hJQ9Ws1cTIqUEs/IPz7EYHcEDu07q3lkzPApQMvlco8Y0
f4IcGCt97XkrLbC0Q59iahyiOLvQois+65Gwejq8zWtwPqSEd+VIgBQuv3ADKqltw+41j4id4AOU
MO/v7N0zgu2Fi7rDLdHBQ45FTYbq4tYECnD1BxUTVFlVR1gwj9p7QrX7H9Ae7ql2Xu62FB9l6MX9
zCj823I14C1+XYKMfSfUUl1UYZXtJpByWwRAHD2E7rKhAOt2CC/D1gspP3Q1iayhVpSrzf+dJQ14
E7oEBjyklcHWKFWRhHeGgrC/H5h38vPeT4GCtV5eV5hbucLda8c8+lzbHFWN/HDJSUrw6gHOVf1P
jbKuhP0rCdRC7w+tq9k/4NlK7JcLYTpRvL+wOMmOTM4llecKbtyYGO4t5eu843hIBeik3WQ+pJ/A
DG7CWz7u/wLhQUh2MsVzrcEujaUHYcv8Dhrzn7xqyHydTirejjeuhXDBpsWpZH1WXi2DvRMlnkiR
ILeTuphj8oYnUVSefSmt4U6R7+Zf5lLXlPm+zy6vIjps3+EgYp3MOu3PQ/kI2uI9aF6yc+PYoQ7H
JwCiw+oJ+nv7rLQ7puG1m+KtpMQEFEt3/Bl0G/J40RktNNQpl8xoNdjU1o9BVGjVXW3oxm5DC7Qp
11gY2PmVoPUV5+JIS0F1M8huo86loWkbc6v83hqD0OFKEiH/JMOL0EldAi2Q7oVgNGSl3jt4U9Jt
MR72kwVzKK1/QJxGb4OaiHPuz8lu6ErPCz3Ll9jb+8v8fGQ8ZbxafKVmFw3S7nZW567tHumwgpgh
DxxtooWshjwUypK0sPqyXbvuZ0qD8vugndqhRbwq1fAUdGLF10z8QHTjaLiEziGiwxACAXDpgHbX
Ra3r4kKvdqatcFgfrxp48nsCyJeShTdT/AqaKHPEf4xGBAsBkRXaCwVv9v4NbS1dPFiLMWACEKZb
OPx2ouOtVbS/AiopBaSBZ0WaypzBprz0yelQQuQAbpQUqkhysWqAH97236LbHT1fDn4GVg6nwFmN
4Wvcz8cg+TyLP0KFnkAV55wtKy1P3xaSHvna6xdHdCP8ieo6XPd3ryb1cjjhGJ8DdUiZ3sGKY3cQ
XnFWItgTHAZlR6YoJsDt9a+JJU8Bqhe2ZzZudBONAA+N5ojpJCHc+uQLkTyzwYoFOF++bFZ7e3SM
3Apqe7zgKerQtQgm6sR6BdmB97dFafInfvExlIqUii8/+AJMsiZFTDXctcwjjzxGBosvE+rYt5+k
Qvc8ZizKf5ji6F87jqV2rhCqsAnhVnwz5DkKRpUYVd4s2RrXeiplc9/IDpuOv/KDhGl7zeVXpNqF
xTUpkrncPJx2JMwD5WkMQ54vfDsHIZDPsqIBNKF7hyDtToyoa5N0CV5uUwa8qNx5N4NRk7W7+k6W
WwRQf8dZWXhN3wPniGg75gUPMspX0yRTxFTqnrTJZXRbrauLHElypkDN4VF5dT6CFpd0vofBQz0C
QAKK+E//u01jvX5Ujy5utlnfsm+I4uxRzk4xDeVs0eduZMi6wblysx15BfC198wHphQCHeWCEXBy
kotNsw66OHOLwjuJVO33V7zDhp9EaJGPr0Aupg0XPOptG+4B524l5F+eHTr7dmtD4mX/8cGXZUX1
HVxvS2mp5gxM5sX7dhraFa51lpevMCgOmuqofG7rEWyeCXfwownjkuUslUm46bRyhHJmRDbOdU/T
5yqTveeX4mjae1wewxw9v1LRl2UmETrycTkEA9ONEchlbfBGG4CPaR/TLAOZBD2iLV6bbx+1z/xT
ZG3+Naia8dFKeLLvXnilDD0Hzi5k2Ce8T8g26uJ4/PSoM2OjQnQzqBUy+LQsZtJ9/YJMiEmXZGoe
Mwwsnbu7HWi1IlTICYhH0Lh5y6vkA0jrY4yhNxZfQUW0vaz4wHyOZsiv5GXXU3hdCUEqHq94WpPh
aV1uERyrnrBgf3/SZrgkCiHef5XARKWm7P+nt3mf67HMutHySIbwmCO8s03bQTy4EMepwfgr6kaU
MgEj/RMe/V4wWKluqdJohfRwP21eWYiqyYmg8boKqcx+TcRR2i6K59WippKczkHu7xbhGln4RbTY
7AZk0HFpt2fumdzYLoGrOIJZN6G0lYs5LG2P8QwHINbXqJOAtEw67uU8dTCA5X5svjdMdLgX+p4K
RdD+4cxdff2M9Cu9iRqui1jA0mhh1o6bdjkKfbkEAUjijBI6zMj/sCrq0wxjgBOfVHbJEzKo/VUN
dmatd3LFE6eoMbRky/Ha5OthjfbrwNKqvVD/0+RC3q/4r9S1n4wm3vvZLF5mLUeBUnnoQ8YYHpx/
ZMVmXy0fniaLiH66O2CaL8MYC6mZ3xquQCTWW/3DHM7cdAmliDHGvW0DoqhMCrqq7T6YVbmMylIy
5s1S6FVS+/Nx2Zams5gzQltosGqEtqTdS01GmVBak2erB0scXmy6acHS2J/FzuuKPxwVj/d0vmLc
jO8spgeuNPQ0SxJOM4IAkU97paPTT8kjfSBEvtW18O6K5p8dAI8f2cw3gDJCc8YfhM7+xSkC3yH2
r7eSzg99Tc7hXN9T8GscfPDRrr0j48fza71numteEviAZuZYKgdvvyVeMu95KHcoALLEpiCbAED+
FBbHEaqB5bAqyuOgoO35oTyOMI49GovV9jFlLpYqvdNuhsjM4TdTV/rC0kj6IxFq6yJs46p3PrH1
xSIZ62L7eEDnev8hjl3Nw4sKNQ31LggQXIw8Jvmoce4gtUUf0ZZVMRwnXr6DEfvA+HTHvSGCLsl/
qdbaqinCwy6/j61G7v2pPF1VQwq3gRLvnK7g1FeEP8tfQNHvZfTDgwzjEUTyuH4iklZxL6jMvhoX
oNVMVRvlbJEeu2MDKaA77+1QvVB4DfshaQ8OT9OMv63JRTNsZRq7CxwwZ1eFnw3717H/I2TugZ2h
5reZZcWivQvOj19IWiVunmbEzaTmaqcFMU+6AF0KSowKyDGUAgpqM8BIwHIx164D4nRP3rSKgGqc
Vt5VBuusxoRLkUtyWqYPtOnTqGEuFmcVI3xgLzabQKRroRbh/dWJURl1al1NTbpzqTqBCD3uuPqx
SKTavnsXltG4wHMkbioJ5AaD2qKK0fMd54QYShMt9i3AbeOU6rHAUgvceZnyFa7M9RoXHJ4nLdCc
9SwlRrG6ITRU5RwUIEov4jc6AUQSyKV1wbzXUdCirVGCneuiXM8tZezE5ZlHiOTJmLUfZuCvktM1
ld4SiC4Rg106Cg2+bFzjZ+saFjZnSEdUfexzEq6G9k77obiM/JaFtJ44VQkRw722iEa046ZY1ek4
yrlRLHgHGhpuu0VZ6y3Ft2olAt4SqA6uZK1i6b3SclNsaJg/S4npdJkMoU689uwqnAj5QpMyIgxK
AdtTsP12Cn7aisa2vcBYqmyuo3fYzBnfP63Aed/EGenHVP/+2u8zDFbVWAjzV59j2fJhrZkd3NuH
D+oT4EtRSq43U12vuf3INluBAGSnhU3CuUG56lQrmDVsy2Ah0xpMf+Xs0KbHwgkrV81xdiqf73Yr
dfP/CAYKAcn0CZjCq2lwHmFZaeQhUYQCIaJj3nps5KIImr89bD99EerfvJ8mnLLeVuKyff93knXU
Ep68NDoLq+u3di9FfHAc9zLrFd0WLbBc9SZ0eJmACO2z285k8PvRJNB/GTLe790ZZPunRK6hXIuG
KWD6LdM9onmuHtaFG1I6mWDxdgaDuPsM8BRM2/argX4HX+WOTVIPEjqxjlKta1lF1aJj9UUVXIT9
SaboOexsNWsCsMZVknabOIrmtUyIVCbHxId/hae/zBvm2phuaNoU7eFu5NXg8fxjee6wlEy7OYgO
/FFekTGavvnSLNH03JW/b2rkE0f09Q3RtISdWTFVdixmpvPvVuvVAtlI+MkpYARN0pCVYhd+Ip8u
0rE7HyTSEZWNg3LDmyPEd6OFZWe2s7FJGWjN3jgjA+egsQLowbnY4iJwBqBtv915pYgDsudoXHW3
ncPajgeXjMkr3FjedFKLVk5tEDs4BTpu+GmCyrqu5uSpv8N2R6MyY+VBFjoH1IXsbDf1WfntYUOQ
3PdtBBQxL21PwFSzAUce8GBcUqsVi5XxHueOUoL4mE17bO8ggbemijGNM8CF3UbeTPSwrLkJ9Pxn
8Hu5VtQAZKDvZwcmN9alq2M37jyr6gJagMHQKtshkqtYPwNWxUqgP7ldYz3IGbXWj4fujsE0Khz0
yteosfbiVQixhFyUO+bE9iVADGsgQzuFz49A13gSqiVR58zTHNi4bKHdmLMMEYlSJgQ/B86ETEYD
oeEqZMuJzRZvhWYUv1fzXioA7cgLH65EvqsfVYBZsO947mCbYDONLPBAeVi1nF22CoadFbnIFGcp
8YCgV2VHYLLld7AKUKx+LVQieIao9eIqFab45KWw+ivqK8pdJtisJc1VUJclRErguuWrs2sbGY28
TgPgQE5Fo/F1e3Uh5RqtnOjH+1dBNDfEWfl/YCjKnx8WBvlSUQQhjkK9Rv5NQMSANLxUI5e4BgB2
PX+v25Zk58mmaOZc26AH28enKgXT3haHK3Bc1tRXYZkq4rCDEi4plizdHyoE3Pm5JVSfkwBfkQaR
yhlYQFUQj0EUd+4/k+EzknQXj6RMdPNoqPTSuNgk05owxOPXBZPBV7rEP3DalFv3xkjcqzs+rBKl
UvQly0xQX3LeY3gkwXRYRHeTK521yIBXx5B0DYrAINkag8oEzI5Kk+dlYr2x7iINNqNISeyQwl/V
RRfBvVgtWsKCtiQkiyXowqYFsUp1QwnZZJjx6/6DrYEwaD7eg34UKEF+0aRe/ud7p9kYcbcgae2W
vd1eRgagT+5zBZrccBITFfDQpOor+ncmil44GygRiIz07IuT3IyePWlu/nntFjn5CI7axu0Cet5N
56PbAZ/z8YxRU8zI+cELrBE3dkbgVVvtlO1GBp0AAyn50RiqxmN+4vrH/LWLSEJaag+W+jH8ut+f
6Ro0v9HHv0wKBEK9KkB/HmSk8apP/aoLOP1C1XqixeJUdPVdVnFETH+Zzyxc7Q16XWOvs4CSPln9
2S71ztf9DV9ah8v8mqgV5iaQnPX53lyVFHWJ3VAEuxIsm8t/0FT744e3tFWvmdhO3YSmWgmlG2dU
itYdmkiCLfTEkm4JkkBdMwP3nRA8QFeJniv57ITzZxPzhJaubcvufXdd8P2FYptrKIOTK5/eQJOz
Yc6RWGFTtBI/gTFIBqoG2K5on/NjQnD49vrm+m/HPmA5OgPeu+Zi7EngfvIAOkueKm+Io32kZQ2U
2eRcfcbNhmeiwN+OgYjLk6qL85Hxi3zREho1NCSdbTYE5e3HEFElpJEcUASBM0GxDw0+MLccYIED
ui+1T46JyG3bd8BsoZlHfGhzVcP3VFJW0K8CBNNlCDsBRAkLW8vjkVyphmP+7I2VmIA5t6OGYOT0
aQsZcHWcxdq3JhCXsCnSaRhneHou0Dj5CbFmLRULWDYC7hvLZK4EaAtFgo3G8fHMPUHOAZ0538TS
eqH5bpXwE7iR05lKMgES4R0REStBeQfRK9zxiECEB0qKirMjnsIMSSG+HJnHOCafYWO/oELMYfAy
WdZkCKMGdB8cAVRp/Pr4SJ+YFdsjAufstUpY6fLv++j4BTfqLO7KjTP8wEz1JT1XMkEThAMH4PLv
uKP7MhFIcMqp4UyLxjDHyCsvhJjX77NLLdmFJukaj1ancCdZ6fE3UN4J5bffVuvdnuhLoJFIiJAD
bSrUqrLqzZBkqAG19hTnyGAizfJRNOOe3L+MmfTnc0o8KxQkgtR+LTjt3hmqugmU9IAXAtTHtoi+
D/iAIy7kVtv9GaJkZIIWtJUsdzkFq/nCriKvAFDdBIXUISRnpmup8dMQEFl5YxmqaFKY/LIFratT
1Eu7KQnSjdGWNT33EqIpMq7IGnTMUVnEfV1OmxWAreqEqh0cbS97s/AEulCwXT03I78iqwN8tm9G
w8qE1FJja6d76YGrQBOjNEXWoeDk3y+5Jj4Ita1R/F6s0JjCnsp6ku1h4x+lie6ca95WSYGqztXt
n+sPfz0113e+NbapR88TOCMNmCPlkkvL4DWQWh6pIiUDqVh35d5OLNp9Ge004T9d4iyGQ9JOLa7m
Iyy8NsD8b7hAjWHi6itP+P9xiHvyWrQjCmQzG4Rd9lRrETcBZM14NNPnxnOUQyiD0GuMygCgMDWi
2BAMb08VUmTp2/d3rs2+sx4ZoXDP5kNcPSc9DHYN8TBAqpS2ZS0rzlZoYlllkEnj7C+BXujccvUo
TSlKELGbWOFxg7Ty1Cr6j/F3MhHjU/R8Jq2zCWv2dXpfINNcPNdm5C/WivLLtiw3KEEWPdDaY/KO
ZE8UxbhSYVNm80r/A6ymiSVUQ8gk71bc0TOB242LE0zwlpu2lXjIo0pPPbWmW87jks8jb7pKa1m2
2jWuVx/LGijNMA1G+4K5in3gkpNLI1I62eN2gZgWWMI+fmHUbpAyq1g5J53DFrvUYjAbY99QR05t
a4HLSt9LT1ebkp9CLK2VaPG0PPJUFBF0N9NqIsWXdntY11tVrpAmiTKD9pb39FOgvgpsNtZsePNw
SDbUwE9RqddrXMPX6JNFPLBuZxyGe3CmeiddfNCocRqZNr59/q+HaLYq70th0RMMlq7xaaVt85XE
mbhJIHbbKVrqwTIRmh3mt8zkrS0QHqrYpkYjybPBS9SnEAJXGaTzOzV73tFqodKTgymI5UjIa7Q1
T54T8fZuLLs3+lVf5UvfLvEpjx6g+UCdTSyIVO2vENTLxgJVTg2F6EaShEHfRMsA/NhP8HJSajo8
UJIGrFSnKFWHGd1wp9m/BRoFxqjP1A1JPkposwuIMpvMBq5eCDBT3I/gd7ImeCzas73KHPt7Wp0Z
LUpX9Cbve/FLMayb1sorgMbj+LR4xFlE07iqR9videqBaS2DxBE70AN4+YCZXTQmzcr6ldgT6h1n
rUYm8czMHIztZvlnK0nQ4mC7Rp7BzAeREybMixPtbGreYsqDtDV2L+ubILjIqkoOUga0rzNowzBp
oxM458dYRGBFIPpwpiuVLatHI/itSPC4sM9GOEBj3XBsX7jEjGDRX3OoehBZcEvV56ycQjugkEX6
e4gbo+UjwZam3EyAjqtExLc8Os/XQKAwslz5jyh7aE7DoB+Q4q6V82Tutls6gf6YGyliMIePxfVh
H3FVbR9fVnKau+ni9jQkxuTDryv4ZiBwvUIfEdlCGaiGytkj1Smf2FNbXw25l5ACL8lqtiBLQp74
AwIkt1Ze+ajvixsL8B1meih8fCqtC9wdEOwUGt3X0qCXSqWQZu8AXwA6Rai/MthpxYHvb5ZnQHYl
yKWK4suz9or+IBO5JKZcbqdKb3YYz4r4h5zTI4J0XxpzlYqxjmX4tUZrcQg8W44hmN7wGfFW+E77
SxvPj32+81nkDvEdNxq+5KlokxTWTNmSFZT63t6tksWsfPT/bmLcK7ZBKa1uprYxj1jO9dXs4Pal
+F4mv+kmYpd+aVkYZY7B0BvRRTO867qoD2FJxAZN76MMag2Mt63+tjX6v4d0jBodr8Trd6SBTmmw
O0MZE3Kuob4KMiJkJd+VijkZMuOsLEc4M2E/Iv3gGO7yT4IceoURmvobNmS1mdWZSkPwG739Meal
gH8VYLOjpQY+NMJ4IRDJHgAK4Oquh2yhsx0PPetbWCuoVxxkhTvizSEJN4LhVQMtlfCgxEbdjqTM
D6RwI2x5N21YGpPqDzWNGqPVslqg/oflnL5q087jjtzEMk3+ZfaeKVsx68nUJWXqfGYYPsUgX78z
ILBv03kZsT8fDDcfecJQL+UhtsrTMKOROqTAS1ITHkzoWQGvfZaaPletQnWMRVT5yfLO5/ktGNLA
0MS3Bav4g8Nq1o2O2IaMXlYcb9QnRfbcJRm1dGYVQvXm0z1XsBO7UgXdN5SusWiuBVZOkrnCB+ea
fEuBX0epKW+kuUy448pO0BtW9vTC1QW3paNomSwgIG8MuT6mHSd3S+z28ZrMBPxwvSlzivaIJS23
J9KM7QfGsa/0kDDrwtqqILZbcwEPSPyGVjeEBwLgnT4/npIHIJrTOAgiSZYWaat74JkuhXjgC4bz
Ut3r/axH69lPZHQ0XD+bcUiaogRiyQcUOtxwbrLWSVjLLKiAoT8eELXXIe5j7gRUXCv+buDzzSLQ
svxSB7JL7aETfthB37hpwTOVAgeBLUQXhPsjub+As0BAnk8uLth/GhrQWaw65FhiGLUiPLAyFV8E
Eq7JRL9rGrSAyHnwraDdwFCvTDXyUQpopFHOiJ8H9U6PxJRyWgYOhDD9QgTvBCGjIcuwFxNa/ORz
aGJq++uUPzceGPDIZ9zj65uJXq0Yutj6IOogSo7XV6WzRNT5fPTO3jQbSptADAXS0dBgFSDy9zjD
QSTsHeHWVR7hNu8uKgga1/N+VRwzEiu7s4HMlvZVJ9C0S3fDA1kUnvDEy2Ct1B9i5HKmenY/hHwA
8LrxzH8r2MjzGqk3A06jtW5zc0Hz3jK5rNiZhQt/QFpbB5BrUgaWOVrHdV7AnVMBOwdE10Ia0JZJ
oYzOmdUWd752Aukx2h1T46LmVNwBRO2CP43rdwUZwPb/C71A7c4izpKNIKQkwvqgnjgUPpPv+IRU
eRDOyCo6BvCZxnNDpMSHqPzycqg+/aivFOXx35HOfsg3HuMQhd5Hl/9gznfHTcXAa4brxL6dunYc
4SDd6FLeLoOaIfdn4CIIhsbubO9XyOfnNffw6S2Qe/7r0jseilW/qAhcWKWJeSfqv9KuxPM9ky4h
SY1tDPcAA0pCuOuwWWf+HZdKE1XrGP01CLdlirN0No8UtxbFpPTuhNGFqkTFoql+f9gMpFuJagH+
xrkNHE28wSlglwgtwHFnslumziN3A5RaquChfJeJOufSUj6NHivBidXB1JVdNxVCvnWQUB9F3pj+
Ic/QHOrDNvpcjOKPH8XsNKE6pTXp/oem6UPe4q/ruCLYeIcLtu+sFP4u3aNzbd9tug/3TwDAScqC
tdPpoIJXHNFX+SA8mAWidKSVq+afC8XAC5VlBdz3CbPQlaHN9dLL4w79qoe5b/esiG9sP4TPCg90
kOjDh6lF9n+CgOzPU8TFxgqF7g6Tdaol/W6vaOEYf9qfXnzRTQXRdPRv/ymS3wFyAEKGf+pRPf9t
gi21SgtPWCTA3/O3hy1CJErYGYqyijzjA+Ux+s1RhaKbOUSFDvH95TQTBvDKUNzAkGQkVSgafUtc
fABfE36REic0WHbPLEAswYwSEBjqBv0mpLywZ/9kLsPa1GPnLDopZUfUyJg19swMBmGG/fegD0+0
xSG3HU3QL1TfOyTioSXzkn9djqfWifl8HdZqf0Wx9ycWw7cb6fYlJ71/R7LB1xVssw+rnbX8KNxM
YuWBJHLt7+vETYm6R/fHrA13jSvD8/wUpOzJEdBP0o15ykFH6+OgiPJIxNRleEy6aKST0xuLfFuV
7y360nOUn6uFOQvCY1iXaiVKuf+aHKkwpTvJINuvG8c34MzsTeP9gGTcQgrUxluhwnKVTeoTBmZF
arc3wGEDFYdmQtNgmLGUHYOGwp/SH461GzEqlG1G1th7iYUcT/PrdjJPNgW5Kj6nXQkH27E/Tqxx
ofBZmWEzs1mZvtapXmEymuAqBHZemxDsv+oW9iAYxlBCMPvexvkXTavkehtQzUZHdCupbQIfe9Vh
QHQbWBm3NC6Da2TfziQhmCqALIummJ90zuFs6M3yd360fEwd/rf87fdL1tOK6LsnrkDebfU9NlLK
BwJIBL5pMLPCrpbnN9GA9flSMXPxgwJA9WLh0xvFWmFtKDYRFI22IIJoc20vU2WaB9roSnXf4pNo
Ktqsdw1LkMO8mwp4jwGf5egPQKXsfXHio/IltmWz7fQqwbGssA1lEW2jni4ERjCWIdbN/B4cRUoP
K9LJBk5U3og0/1RJIxidsW45TChLdpk7P32dwnTlkUYpP1LUwwKARiQXhJd9AlwqcF4ONapE2uyb
cswhF1A8Ie8JjU1tm9mcKNNwA0J/UzvfjiwykwG2wj5RVfrEjgGM9dyUOWClkf3jTj7NmhLJ2OYT
Kjpg+SipSYWLB/35uL+x/np86rTMpshduw6Q4ZrcZfln98p82q4pPjWw+PKDrwtL7qy2suH9xX/q
Bips4crSVjmzYKhQZQCZcPoU3y9szqX+2r/d+sHVWDV1JTR8CMGvxX5883SVmEHAAWnKbgHDlN9q
Na7wMQ/xklFbgwQ584WECyFAmUsk4/BT+2SbBtTPG1zRvMsHhTF1cpOK3zsQGSjaobqm2w1K0d4o
kEk/PMqnCgSY5gc2yRaSFJJJwp60szb4/03GAIpcdUcCxdNXr+PFUV36MSdX8qdEVW9fwGs4h+Bc
dGwJ1WeHrF1r/YKHmVf9SOYUr5UY+KRjL2QN60p2JOkH96Kip7tEIGaP94mGIQL6+AF+9dWWRNp+
IrcYNVxigRSNAOTatBaUbxpEsgdOn01AEue2npTwwkHSIOo5qvdl3v1dBRg+kjPp8dcJmai51d1g
NWtrIAXVZIYes8HAhiyeznsJ9eVrcXgo74kVoQ2G+sWfbhML6kKwKOcb9PrTHOZpQZCw7vgh4HSf
OZ3+T6GZgU0sHHLPbvRfJj5cO/a2TmPl4EGJ1CRwB1oCn2quqmDCN2RfxqQR4VQ533vd+8lX6SWy
GeyTZkP5BWPlCnQprfCcRmPyLuNETOP+rLSU3XJx/Gbagu3WuLB3MTY7cHwyghlvbLjJtQvW/2ff
g8INURV1QXPm7M15IKaj4w4J1z5OKnmFtYzu0hNiJF0BXamyHIb/HoECJb+86tBVCgjh67X+z0II
Q4Zjuyzrnpc1dcaK78xSYzIO/xaDraoemzqNBsprfaP0hWGmPg+h8RJzLLjWcDUxv3bV09pu2hfu
70Y40oGco3vLFl0sEubiBmwLfpcBiHagNrxRG8T+kXQrpEYkAJAT8fnhwIs1EJt8SL0EA8JwawXr
oGZMGQ3low5DnO7lj2SBzhm1h8SLvje+4wpYrAqSONMk26lqsaBz8Gg7k85J0yrWC20Anc0aPYQK
xeuQayy8Cnaze9pJA2AKnC6WSIYlDCxjvjN+nQasLfT8P2cG37Xgm0xO1T4Of07e5NmEAEwp12YK
sUXfRg9wJn2ICJqdmFCHVjzff67BDFutk8obuwwQuoXT7w0tjmuBWrukpuCtTlweigOL6ruq2Exq
iDMtcpAjyRU1akQD0apKkhsgf3tyd8TAOVw3hOXTfGj9iwWgLh/680XHVUArulqxQXeDr+AAfWN5
bXbAC7x10nGp/2ZM+82YENPL2PoRnGNDB8UaSZtUheLcMm47/Ux9vgBgdkByRuncZxe/XFtik3c+
NYIDfSpzKHNzSQTdkkX0Dz4zKeB0l4MaRLC/FQuL0ixdpRr1alv1bYu1kVKpCRoitaZfMZ7tXt+L
+t3GwuEfseumZicqZUCvyWNv3piIK1aAku2zobbWlUnHch9fDuhu8CGSoH/v5jIIxtyoJkWzrBdN
djmMk6Z4Pe2zOUe4MeIbrTZrQv8hhnSU32POIHEf3m6uAhYfhyG1j5jsRnA5xOHwbs3g3FSy1s4e
qGnPfKN7RcLAIAk121k89xUbKo8O+w2vvmZUa3FircBK+GX171IpQy/71dh/Dr3WNLWRzyseSfL7
RLHtr+yfnHdx3wcZB6VFz5jS1R6eGizHgbocFlRRk5yhJhY1fwohTk2JgYzBc9OnqwTk3wsEph38
oeGnUUJdUvRya0CWccKXYgiaWNlCak03hQtnU57Tfw+WQzcO05M3AZ8ZH6aswygkg5H/285t/pR9
CfA+4qHMzLwwx8rTEPKXxQH+qxRmgXeC665uOProTVgMuGl2mUCdLVPDHw8FKqF94G3nkmo6iwb5
GYSVK7+zWVn9nsIvp8al8j4FttxImuE+S9ct4bysIfEysOpAr0uJnW2NnwqvVlQC7TR5f3mI7gCs
oxgQecTR1cpkmuYVjHo4wepg/tKsGDxK7pFuFgysO1E4++XIL1deLKvhv1H/YR3VocfIC50cZsst
rrcWgKdd+Ff7HdUCO1weiD2Dz1hKstZZELuYuCiP6RIeN1me4M98Ff8lEzIHw4EiNDf3vLesr8kZ
hdjcehitBpGheeCoMwanwY8y9yi3K87xyrcjdCyiU9zYYxiG7ESTTg/hL8Xtp2bMBSd4zRnU6fzF
jPlkFdXtOa3GXwoMav+O5PrCWjm1PA88UbR1AC9UjzyA/Ei4vNcp3rzesDRS5E+HSSEuMY295Vzf
n3YLhGdfQ4TcmxRkQQNUn/PVShVHhmkn4WVH1XWSwuoPjo3cSz+wgC53bqEXA3HOFV2owOGZ/NJm
bUNjeLQLsleRKOOnB+FkygcK8MzlkdvgwyflrEsnsUP4Jns8xp6rB1BqsKTnHNY17BTbcLpf1UjH
pirUfEL0HuupT3I7q9V3W/K62AXEVhz1vXBuMWkEfl/4tAZoTPzm+zZLKThLKXz0PzGNOpsYKhvY
xfYci5zwX5n5Q01WQrzhiGlzC+DFWJivF3FUHG/EyIvctPI6goTDoApfmCMxGoQYbQJxrTYj1a1n
YYRcEIcQJfdW6vlQgV/cRCYAmpHMJs1KICTP9VPVg1zFnTp/YS0ZhFZpmLwt0Q/gZASw6dCP73Q/
GZwn+NQCWiiteyeY4yVBNlM7LLfcuI0OkizaVtT54R8E9LsIeZYIKvb9CxIZDRZGqrLO9B7p55pj
92lXpvwKfptZks9OHlu69WtrIGvRMRfT48LK8KiEbxrrMTSw4cbFtV99TXLuvEi5Di4CeV6h5cRh
QeJ2FeQ9JcDPl0wVKdD526lXDaCvK8Aw0IVrQLYIqAJm+GOj3SLtZATg2Kzm1bLrylKyVKq07CsQ
ejVuHwVEYebmqnL45JbKMRuOX7zhJjWMPxsE3rI04Jn8/nIcRF9FY1qdtLILkVBLMXnIIao7ueoN
g2HiRxpvNqw6S1ECgME2VlW7ktkl77h49BfR3lkqRQqkNxz39b6f/S6ECRncXL6+iVuWqtoYAw1Q
eRPL5pSFYdEQsMJ54qCC3S1AXGi3f7e3otoQv0mGFd3IGpQTrDESCFvNwOLX4z5f6U1cNQYHTNEv
0bNraabm9i247I4FsUBI/+0phQwoFuUAgUFz7Pz746wIb6L/bmu2OpOr0ooDRgGYxkBkgwMgwhti
lZfA9H/tnsPPWieOyDXRWgvRXgFkFwUG3jNJHGF327M3K0YnibmdFztvyiBC95TJS697bwQp1L2R
sAAWigsMGnpGlZfnOMCDMeGERLdI3Xlf9wwzs8h7h4BWxUaRy5G59C4+4aVuudiGLn6YEvB5gGNE
7EC3wfUa8x8gtDIBsWRIgMdrGFZqP7FoqnkSjvlRtYt1XxC52Rn0r/SZpcjCAJzhP3UYl/WSuwkx
JcXKZMqwacEf1fZOVeuSj3MT1reZ1fp85F/d2y9KzUpbZslDH7rO+DQdBsgI9pcoiElnlWQKbLis
uI1Ql6rdW/4qMYOEMFumgYMarn4/OJZTIbDM1P8lfJVXAMVGEpaIslnkSPdUPhLpcvfhrKYwnwH0
w/R3e/aELFJeaKEUDWDPcg+GWSVuVnW/kE+CSrF4Oo9b3v8pks9SK6wygNTjY3bvHacPj+IYxRxb
1aWKPu3hPpe2sNGQ/h2ZIcljoW9q5T3Asgel8lf9kPBHyWDyK23I4uyjC7cSyxd/OIEkWJZvx88H
KkXAwICw3/KRt4cFBiXPPshPtay/tBz1cpjc+szcCEAbAcEKU+JKywdmmwEZFXvogMvUwcdQd0jN
hJByaCpbUp1863wyXKeQDsRIC+AUradZSu2vWfQYniLn19MgbTqdR09xGlXI5wtZF67OP54MNmVr
RVpy3ru2j0hL3g/FUngLIUgh36pir8svs5qbe/HlEQhuUec2vJH9ItV83F62/6otuhs0fuuNXsF/
31CVl1vyQ8xTpwzcDASGgMhjYHnB686TF3w6fMFiE0trXGOa8Fopjux297Z5po5AWyIepyMYbvKy
lRnK6qXGdQhSfkeMTIspSaRIACf1Bmm08G+X3KinHCs4OIzSv6xNB3xhmc40fr5DlZWatwGTqrCr
tjekjhMEOwQ3qBhDSEIGLIS9CI0YRMU1TmMl95z0GMBp7sUHGC6Su9sHh1vDXMSOyfkT2Uee4wJ+
+OA67nrnCl95Vw+c9wjsgyygo8IllBSSt7uYY7Bl69XO9Guz74h2IqSNxVk3HlcX3BJf1Tm4LG8c
9R+tq+2PU0vhNMAFK1TfjAthGEUjZWGqadW5VBlyqzdgWS40alzqcCnznkMY4XOm4Vrieorneh2u
vW13blTfKV1RCAshF9/bO150JLpFlPqPUrxh881llu5vvdjQK3rnmwt/7uU5uw6/q4hZL8+sCboc
STIJlEPy7YOh0AGfotNr/Pqw6/hAfkI5XdWL917ZwXPxr6ydBM6SgMoYrjEAUTX+9jt+uEuxsnrS
Z5uxwaMYHPpGJV5kEHe/jCSqcyJwleEnJKi/X2OnX3K0tdHhNTvDUNLEgUbaaZCm5RJGj2bEHNcc
OTEvnnTv44s3m3ZLIv0nyAnZUvH7zgGPP1vd1XQCSEsHIO64jO/1GjubLwscR4qkGXx+Yg8VLCx6
LoDhOJojHpQhkHBWp7CPG+yAMjC5cSQ5p31A2sHs6ezRQs/E/25suKotUKLYsY2N/gUKWluwfE0M
WgBEOq9obf6xDo4PLVjZOaNNz6+RwIQ7k9tMM/R0LMivJlhWZ5zPlS1FHYcigWPsSVMGrdFV8mKO
qgKsN68UmwlapUtyG4v769VwTvcmGarAQAkHhKLnHfVIIQhmARN4qN2q86y8cKS/5a0+gqTgZZwt
D+EYdew1nXdHX3ZItTz1G6hDkXEVGITSz52qpjdhop1H55u7C0frdy3N0VuYoUVnzaPzydxNiUvu
S/Lgk+DUbVI5SxrAgOupP2WWTAqoGCQAuGWvzrNr/Wz+LxErFxJP1mEi0zlDPkHjBcORv6dUidwP
JrYCxlXWOwLw8c6L3R3CgzF/D5ELzeR4glDaWKJh7jiSU/bS0Ylh5xOHLG/4X964Q2Tr3QdzdOlZ
nkTHdFRe+DNSHIo7hWCT8cz9hBzg3xRz9+OYaxK4QydX0WzCX493REfsjVl9/g7/Gs6RkpE8JLli
AgI977ollNSBYf/XOG6S1M4iIvd/gnxTQdZRbGiHfHTA2crP4LNGQNqdZAByXPWTfL7LKg8gwuqM
Rn3HineBPEpFY5S+8PDeGRxdTxE68A1jnRSgFN+PRMfC2H+tXu0SxPf8MI+BGjUua8HN9UPKy9ga
Rl93tUe1nhjLZUAIOWUuQji2NINF9r+HUaB2rMb1DIQzskZL0vgv85yaPsy++QKca/2slr2XuA9D
Qp1e3uEpgsEqTsvS3c7uEVX78YaxLWq+CqluCo3sS6S5fXO5hOB2aQh/3sH+Y9LyXn9R3bfIaMvZ
TKaZg5e2OH3P8eKJ4DBLfcCPVEBF3BOViN3unvcRM7IsccFtWtHX2qLa5VTp8drNW7yaisfRo7EF
daQd9yPuFmkcJazAbZPvQVxZZgnR7B0QNT87oRW6g8lxXSFNr4gKVGBwMMPDVxcruH/UPNLZYYx5
IffCu16Zbq3KrVxzUhQwJctJHCRu1/V/r8oBq0cJtp5GQ7iIbd8GlDx5GVGgVwKx+eZAT4tLwbxK
a49NKADXDonBTJxu89cjYLP4rmrohp3UwsGIg0ypty9ts39et0W7itMHVqUZo7DAXVIQRPX2Pgvv
Kr3PpOGf2I5WDatoq99p0z7zO72lXVC9wzU1ZJFOnVQ2gspL7NmNCrPipT9ag+BAhhhEUDHbZdCf
+1eBhlheFtJiX5E7h6XqOFHBFg56fIc/9321as/0QTDT7ZmGgo0C93zpVEAqN1zklgcF1I0dDeed
KMvRNWMAXnYaiWXBpacMjUdLMv68y/s3d7IJgzo+gATXeG6Az3m3q21rMC4mIrno0biKbbQtKh4F
c3XqZ+VuIltg013uC0USBITO1tjO1eQiCX2dixL9zOuwBx9WTM1zkkUTjTCPbbIv3Q57UEZWamMs
MgGN4+MSm/Uw9ilhbBrPoTItC3UFlydDSHuYJOYxIdaG9+4IJbhSEPe9vEzwFPssY+D/WzdyyVfu
WaXt4SWVQGl/Hn6JTCZG78vYsaMQfczRm6kVzLmIXVr4dQXCVRIg/W3Vl6PVm40eBkqykMBfm1Ku
2ksuWiXoSQr/fcgNwYmegKwLpm4ni3kVh/rc+gOChu82ggmH2DesOK+SnNgDJ1hIEJMe3ajhfztF
kwzJgKpjHS/Ro+tEFYmk+GTfxn4I/gB4jZQ7ibdsm/vsqiJRXckAjOKAdpQ2fh1VWzA5tdoEYy8g
IPcz3/b2q+WXZyaW+5s8ONUK+LppySxsZp7icunv4+otrzzdL14O1fnO0tdI0HOk6wR/DV6FQ6Gf
6W/FRe7JHR8iXYxxiiR5QJPitoAt2NuARqA50qzeYK7c5Z29VZAj2vVfqAVnUPV7pmCJ9+zT8UHx
SqHu3Qo4Bc6isjXqzagUH8yjK30YGbZes/mzRFPt7Z7fwDBi6vSxIe7oMEe+yyT7zyS2n6qeTrD2
4lhoCtOxHhSQDNVX/vf11GXz1/O/hxzIXnyOtoETjwmQuTMvQd+iBUzY40YrMXSvZQCyXtJbEHQU
lxf+z0ccTWH5XF3y6ojHeG66Tyb7iGgBooV6xWoRkRvOVrzQ5MHC8MAJoXnsnII1XCiKYFMF3ocQ
IuUaMlfIcUoFKVuiSauaOA72n5/DTs92BeEgN7LjJvcgzlG67/6IwgHRF6oiKJFiZdgpl5IIUMPG
r0Tf2BvvDmmAC2ht2HgquUPmGNTwwNcW8dfLe+LguCdnWoj2Whhd5yy1LyPeBzAobrA/ghasTXz+
O+P0m2S5epW7SppkeGpMnwIDiSiRDFoTEqGXmlrCuecxxhKzBKWyi8WiwnmT0Vql+8p6Xa+rgjH9
dP66jQx3qpzBlBI1947sReTouOQt+8EhKXse0WtWD6st11RWTkIxdlzW56doLvaPkKzvzqe1+nm1
zf09PYHcQt/uMUHbbI0y374JkV3eT4QuKX6IAKNxBe7KDP9Rj076WcxWjicTWKQzEvm1MvKC+3iQ
1YOotWziPKouwHIrQaQXwSP3PmHyUKGcd0+zGg2FuPaNwUkzb6guSwZTU+riO+gFwltJRwJWY61G
bYusbBPRjF+2b8MmGAowmwS9gX8Vnz+Phq7BnbxhL1+4bEeIseOhbjf5XYVfF6E1qgX4i6SGYcFo
pLbwvt1U4GQBKRBaKj/Rb0DsEGm3SzPH3zGEqkBsWemIAUXoXN69QWyX14RmtTDQOXZuRQO/xfTd
uC5TdQ8cTGKPGRlHLsLI7IWgOK7Rg7ytr3fZlSpWjdmiSZ9w6XpsnHkPJi4GTS70+emedG2xRcDJ
/y0112pNq/v4ooWCKvoWJoJ7E5cM73IMhFWklVaZ2brKu9G9u/9ZcALtNwGhwkwlW9eWRAHyDFfI
DEyb81dESbPO928FpnyvBZluT8/gHa87jl7oOH9v8LRefSBzCkwLVnMRgsuHloTiEFqurzalCZ8k
OV5x2HuavdxLjrBdNlDENR8BAah1W7a+UpxfMX2/m3t6OydKYd1rf5O7zVSWjVCbwbaqnX1neGzk
6ewncw/k6f1UPQostgHEvETtUuEVMsV7O6xXukJQJDDkknAiirtmcC4mwR6Fpps9FHX/EoaHuV9L
Fr7q49BTudlpkGJU4syAtymOlqvH7Jy1FxH2PmUAG23bx52RtAD1xHMODnLXSrzg/nZB6czgRDxN
6cQXExJ2r2zDg3qeAcIpZvhjMRQASYCnzQk3HXQ9PBl7w8V2eOUmBtMquYTAegYGDQF51SIvvtqF
KmG5iSnhsTJe56h4KoWgbxqcNUHhMEdO7XV6jN1V5kAFkFB/3UaDt9Fc/Sgd1Zt8Bdvd6Zc4ZgXT
E1xNDpJz0SUbk1I7zU7SKIeoMzxjNqFB0kXgP5M4Xauxai8LGEXuY+WxSeRVvHF9SSNo+eigEEGL
KVol13SfSSJVFpFu3vDQdj+fhHNcIkBYpO2UsN9zmB858oOrsNgJxg+X7nhFF9OTfKV+JXr0lu1q
VcWH7ALuASvYTJk7qIF94j2bLB9Ea2BBiTMlMwbHiYKU7S1VHXqJ10hH6RNHQi7LiyszT4JJZQKk
7xTKyfkd6VKqIYpBVDjDZwOOq0XjaIVXv/cx0HHg/SWrtCuHtRV1l/Ju8lyOPLvyVwENHozADWVx
tJe+0UD+Z9nJi6YB/2Quvl+rpOiO2dEzb67fjXArudYRP/n79lSuGY9caDMl7G/qfbYq65YT9TBD
1RxlSlqLQfFw9pi08KfXa/HMpAKlUDZSq9KhOPHRr+MPNRpjVGxiwZsSspiuCE133tSX8my4UOJH
38DYpeZcmzx8H2sjkakEgKTrIOcwIwzsdj7FRNq8n+hCVEArzzIhyPuzmfZ/K96DEUKmBp1rScCh
ktGgitNWAwKfmEbafoHtvANXFD5XjKXOF9Umjqbye3AsMQK1ubuNjq/0gyBoigwyEgTfif4MYv6P
cNynJcVZT25LqZmkUT0lwcUavdP+r2yoFgSenco14ACyywTMCntOOC6YfsNSBPDLWktzXDqhp3PL
q6C+NXBMmQUM6R5HAYZm4h54E3ofpCfPsXUreaMWPfKHNrpCojbVOnYppks5rrSLt5rIxlRDWQIq
O+4n2Xz0EZlmPnz44eFUyMbprJBi0zl7vGKd9vuNqkVRvj9H5xxhSCTkpqZGwSbysaTC5i4Fn8RH
wFACXf6VwBu5hxIF7Apl0jdhLYt12+DKV8vaF3nZbX373aILNCRpvPXchCE2r3RpgbW7os0xfBfh
mdwta2F4IYZjyBXPM/G0/9h9O5RZ9oT3dvxDK5Wo/HTNJBePXiyuVo3q8wzuHhRmmXew3139revI
z2VdmtG3CDsV1VLFY7svWHNS+AJCGvOPSU4y7kkE3vNo7B+ETUnJr5uIaPAxeDbBAG6PGwFUTjj6
3JwseDpY/emf6VsFNu4y7QwTVS2mlaRGnyIssE61J+9EVd3JFCY0IKDXGagj5Ay75qSTMg7+pORL
2my5ZVBs9mo3mJVgxCInQByxyklL2AT2TCuKyaz8ijiresW8mgBjW8EW/OiLZkSVfbX1ltISyGZA
KY1fZQXR41Yadb9mM3EdBKqFQwF9idbqkug+LMV63fA2YmjOo/zW3QXaVa7DIFcXIDo5Avnf4RZa
X1tWlgpVYZLLfi8VZy7B9kvNkgWbAIMSUdknUEeVSPb9dJdiueoQ3J6XgmMvGMg0YjvrK4AO1OZc
HEm4vPTd422yqyYGDX4eab1VAr1IsuaXOQ/YYAPxz8W1c5stcaBSb72HY60ql3qZGybxslUaraLx
qIOcvwzJJT0apl4heZ8r45ZvUKqcv+D8OOiKtM3CZotTbgtmjOyjdKjid29dd2yLlBNnmtLlaTR6
eE4ApQunUCJr3UyBTn0kJEzsVHbWhCI0lPegVviJ1LFaq/85tiRONS721VxBp5B8vmXlf/7iunpr
4ndxryM+zVD5DoZt9K7jkdv4PHQ22/zYVHdzF98ZRQOwgS+egDTOOzSV6iaa1G8zNhkrDIga7tf/
Q43d6FQinQ3i2KcxSSTLHyKClMcZZlC8K2V1+bKAmrBaeADbURk+gk2YYZIJrHczkKspDzjHhguV
nT3pJf4C7eN8b1E2Q42y3Y4RoB7fihzx3MgeUl8Lmcyktk+Q6Pyt2x4fSnafmROh9K+JZ3LGSHlE
aNwQjeQmDKSZFPv8qDySkCozz/1Y4Lj9uMUihgnWkoPuNHUSZplNiohs2Qp0S19NPi35pyzsyVZ7
4dbEQSeVYXSTotpWq3V+YEhO++ysECUxMqCdB7A/fBVceDYCIY2pRxSPte02+GU0fakYGn/s8ggW
QnlJF+EK2+1xjkeOXC3orMKXL1BX91IWXI1a8YeIkh7xyoOwC8xAx8+xdC2syJTu9+5C3uoLSK4h
2XY7l1oqlzAqutUNhp1YMlcbzDax0iPO2/z/vuso5O7qeqm0e3lcciLRx/aNhMm5ELsaktFIbd5c
JuNGV6gh7/VpTHPCXAd35qwWf9JrOPbPjw4yioAvis93DLoSTOtU9a6dAVqMMyl2cizo8OZ1Sy0I
xn61ByAbEfIO0I4dFDb1Ne9tAfRcXuKe2wEKOTuM8Knic3slyvvgINldzLNERXfS/uRLt1KahOI6
vzxcI+d7Fy+N3OCfkzwAqiWTMUW+FWvVXzhjvdJGBZCpa5K6+DblVWJLSZ1i7SsIH9QJwdpt4Coe
QxHOPsCHqqSQpUzsSoGqZt1jieutHMS1TB/UEf34yE4RRdEO51QPnBKIu5VjYmjMGPEHuRk5nKIr
rY0ENEBE5tbEj+NZ27narno3Njmnd3bijt27QBwbioL5244aiT474KyhEB1CaIhraIid5XetqLUu
ImamKGlaxZ2zqdUK92i5QCg1wygXvONUqPDFOTAyv65LhZ8vf4pBBlGjpfxe0XSbGkiQkRML1eLU
9g3L9IYCFaHbdw4QSHH7pzFH73dTUcPMuvHC+ET55Y7Jg+ib36R2ZaIzvxT0hWkg/ADuHsYd5IPr
5pXhVAifcuO5my8vUqY+099wP4BFjxmtrBcvDA93HaZ7kvBDQQv7CJzXkR96wjhn039Lq88iC3Xl
Mgrg2WKQOWe7S28W0VFezBUqFyw0HjgMpB9xK8wotAOAr0M4QW//0+pi/gkGNmyvpswCRen3fLpz
ATFsgmuyui8Wd1H3o39/kO9JjyOlTYhxCdIFk+skSAj7IHbtlWqPfNL2zgTIjhhvaTFGUQbD+iBN
d+l63oPFkdhN3agCgduq4qoqz3A/W2PQqQD6YBpk3X0/tMkMP6JaAIE8AINMXiSUtaTYdDSU9W9R
sJQeiUQCPi+M3A6unwon0iyr9WyqE7wwNf3IoaYtc6wk3B1N5GZkslPBl4DcUBQFhdYmGA/D2ksu
B5rgcb8i7a2veQ2gTiApT7DssPGvUfYTGjGRPzMiP0bA/SoFiZaTK4b4dT43bL/TEHTamR3w2Q3M
7MgNLCjuOr80lKDKvdY9vHrjYKp+IHj4PRXn3gGZTunlGjlMwBTb06vbzNv4GnvLNp1sq24D7lfG
kDsWHiui/ivBB2XZjYTQSmNLerco8nqlu+MGGYD7eGzYfvbVxKDoKupc1rQMpRAIPXGJmbzoc85r
PvtuOZLdmWsC8URVUdMB07y9vQBysXKbjlQQeezE9H2sBkBwxJaLDRHlAzKLeK5k/Z16nrzlCYDq
Q2L1ycHCjs1PJRI7XzWc1K7RrRojebZfozLHWFHPyUIO1PDELa9UdWkOtIxMloV6BD+y8K0u3NoG
Kw4wRD+fT/xgN4bBJ3xfHY3YweJim4AB8MuVsGOJN68aKSOq0yxUebIcUwHc4Jly3avOuEFcf3gF
XG8+yyh8UZkMHgyO8+oTMZdZZBAiTwMeE3Y4kRrQPp8BAM+FAvLqYTt/hzetLIowEhmO10Br+LbM
1/qi8PGz3Jl1FweChSlMurAP101jlGg2tS9Fl8dmd/vGNW+ghPAQxIK+P+bQx0Izc/gbwJns7VuU
QBHpQQCBj1PXdhpDcYcWGL9GrajdsHPuvgXVw8WUF6C2W0yFzbco1J0ymzTEoAfK2CjPlKgRlUYx
LBp6dV74nlfeJy8jPj+Jixd7BWhp596VExlCXmFRpfVQsUXDbzzISy6HURatKct7so/vKXnTKZ7k
KemzPjVQUrJhb+lN4fKrzXwH2LiDGJZfMw9igPvmiaWGch0+poIYWQ+Px1RFpH0wISj11O+Bj6tm
6cRKH+nQVzw3OhGhhCnDPITTuP3fNS0qvAR0OYDA6/v3t15YoGIK310SRMnN0CkiPHoZ86dHM2e4
EwT5aEp/b05nZfhsRodQ2DZ6nEr8JPI5BJSBtuZ8NdPkcDEcrgxAdZnby1cgVCLVTcvhJcyOXT43
xGDGHJ9Zu7VBTTc0WT+SXNCZjwkwjnq+9cgBRGZDTgJowYvfcAbIpa5wDOSJfWLMC4I3X1c0nyMU
yYX0wXTt+RJXPCVDikD9UC+ZIAKaM+5TDBxkqh0xhU3cWAa7VHqwnBPSYae0D7WtvTCitp13O/qU
7afji4O+NZbsPlSUUFKR+T/Qm7BWuG0ZG+yMSIncYrrJODlljCsKfefUeC8AKl31oZWFD2ou6xUW
XGY67zhVXwP6YoCLURPiN6R2vgN105Hkci3jDVuipG2+23pzZmjlyjveWUSTIC2KEdxCVc1p2w/i
IoGv4hwIrp82vHoJf/aVE13ReoRCP8s2Zj69C7XUatG2ib+CYfghFyyc8lENy4WEmsxJLTsEkG9x
p3SmbFsC3zyWb8/irGSn3vMlcGjZcj6T+gzmVSV7ljemvLWCJsOaFCpDe1OCx3SCF1FbTsg6o8Qp
7wa0NSbuOtB5zA+GP9KegAnWjAV1/hC64uteEvEB85XP/ZwIM8gzYD7DshOo+ITtluPAcPX3tHQp
dvOHBcW0GLyrij7bMhPV+t0gthTbAGLL7GD+B06KfrdsDDovTLYvorcA/h+FHdDknHTQG+Tyoe41
bHhx4REJL+g2D0sCLIpof2bR3KNB2pki4fCSNSQVLTJqDTNu0k5ewjH+FnMDGj/3LL0avLY2UdMM
j+FJIIBSGGNDd6BcW2veJim2ehNgLTprTy/F90XVgE1bk4cNK4skzTrrZmLCfyZi+KqGvZZxODoI
joHOfQ58XwQpT3LjNKQcQhc4TrvIdCarTNcbJ+0TQZd7ybbTXFqFqEh6kyQjdHsQAVZatpky7Ukg
bE8WHS5YBw28OU77zOEI5alrXYiWzTrGtgH1Tg8bldyF5pUIFEJ3BlfCDbc4hdMwVF5wJpUzj3Zr
uhbAf4NifGb+/wUWh0djAWiv0C3OC4qTY4dDnjYHOqcugNXT6eDTKCdZJ+yL/aJinPsZXRWXyMSZ
/z4mv5EzBffS3TFN4Qarm8jUCMuOyD6G9g5iIU9f3hpwItXIGwN5kNmjzXbEQG7/IFR3T0VaLMut
KMu0r3aCFvgCRzxBXlZC+wMGrLLduYcuSnIzZmZZOBcEVlcG59QMv3OF6vuagp+CLqvglLvuyeEt
EM8dCg609TTq20iBO2BP4ibbRY7uBwW4aHmVKm8IWvKucKdym1yxda+5eiq6ddjnKDV6q0TTTmml
hoVMDY8VHzwf1MbXJF3PgDFK3u1e/X5nFGiSTQHGEGqujR7FDiqr9T0Eu9MaaC3zEud+9FXnBd6W
uxo0r+gbAIKmnZXFfDnVi18awqih1/x3rxwvXTL8Ep3b89vj4Id2/YrNSpb7fp37dribMS+Tymah
Tc4cnd7UPrJMi7WtcPH4V0mswF7giRxc/K3eRjEzMhqS0JcFm5D7TvNL0hAnlhG7Cq9W2IupaNpg
y+Bu9UyilogYp8R/3Sd/EcqYWDNXFTfcJ1ZgbU1g0KtGE6ZKSEhbqFgWn8bgSt/L3HxSlv0YFMiI
gqyJoqy+e4EPmteLrGRjmb5ORsE0smpi6HSRV2eIPsmVMHeUinqDeXDMGaMNzetzohRtRfGkSb6+
oFhniUCteALc033Vdz+6JtV5B3pFbOuXd/e9PUYwvIBUeKHXoUcf6D1K9UefqD+rBKxv9YYZmV79
5D+gQHJUWlwC0UQfSCqA9Q0MyFw7kA79mTU57AtXSipvg7uPDQBnKROwARrt1X9nwJTgWhwBzBDA
sClJha3+HalbvthUOe+tEccJXdR69/ddOQySRNprrxbmPYfXlUVcQ2HwJtTDeuTTDymiQe7fc0SJ
nVLgcqre7GkMITm8p+2JxwnjEkKwq43pPjsdZNGOHO8qCDScDKINj4Nj6LVzSBro3uk5uPIHPzVw
1pNTyeylINx910OLqldYIcg46WvRyk+Ag2gMB0FDxyB2IO4rRh2MdfigN2RP3+aTrBYphdDLFymK
EEOt0I7XuWYmXwp6kswl6nD4DSqFVYw6vjBqlAf8vLSAymlGYAsgOtBXGtq7pV4GOr2T97S3/9Lr
6pvvtSqAnPV6wj2Bql4NsWDwjK/r/YQimVC4BBK81NzSPn5F7hhYCjGyynMKU+yZUlDwVMeG19y7
xYJHLw2DCzigGMVhsYoOEeUPe09q4xHpisTIz1PdKySyXxJVvpHPqa9CEHCvg7D3xi/2jUvJGj/U
9EU2KsFlX4+5UI1HHtol23GmstZ61vkruhU5lg7jZN+utyz0WCh472G1LphhUAJXrWvEoTsQEDlf
4x91M040g+10mwzEJKX9yz4xrAlMyH8hZUg0acpjxzt9bktVKMADB7dxJkxslXgFjuFktbmM8IdY
ZPt2cDqJvC4bburWGf/WwOCHgBgM5pucvPzgs9Cq7rYTww9bQWEPpxGVsU6FUtGgnwR/Uw8l6FHf
jSbyaNeTyO6SbqU2pmZqQ8iTq17bnM/vcFcv2f1uZwR+pz+umFmQHRRuWvJODiAfnwUCLyreq7Wc
PpidnqceOcBElBi4qmmYAzg25U/aDqhxwjciEVO+gQ2iv+tzCkkeO2vNWDv1KgxJiuKAFesmiJuM
NeECrcB83lXLRY4pmXssRQOMzHnir737JgxiDe2fDzJMTFxDfcagJnqR9vXzI3Nfi6DeBKqiAz8c
YKYBjGtl1NpP9aW0r45LBDKp41yyUMUprtAL+pij7TfZV+m+HHR77O2aeh/pTDnLicMO/DLJCH1c
aKRTJibuP+2ry2FTH5M5pZxS4Q/7v84Dei6bEPSVOBX/pdw0jWSR4DQnCbJz7YGXAAktfuPzl1r5
uehHRAxZqO9er0p9AuZNMSBO6BU6DBw8nBZ8ImEBc+uwrqQE2DFWP2ZBQUic1xvE2jg0jkz5nToL
9Q8pfA0e1CP5oH21WUpOGptFBJ4Fgj0pGMPEs29KLP5cgrGBV5MuiRRXxzjuKtBo0DlW2MN3WGir
dZRj4eZ4hOjcL3Wn9tfopakiQr75Rfq7NXlgXWSBzb4IkPrmOufw/M4j1KphCY4JB5rigL5RYHE0
v3b9f/U0AV1YV3mEP/D9dsjOIvbGQhn2iJzPvWCYI6yOemxRUIE23hLRg4oTessrpA3B2VkuiyqH
HJG0Z6X195wxWNNV1+TI4nQlt5Tdp0Kdi/MrRuoIe13JF7ozSo6TfUsbi0ftJkyyWWywPtFY7jX4
P6CDr+gs/21fk4BCTXXyDoutZJyu/iKJYI7gPeCkb7Kqe1IuGCMIIF/ENljEe6xNGUJqe1gTR05z
cvkGXa12Bsu1SzaTv5mOTHUJbVi9b8juP+c5yCjMIwAJwBZgRQOx74SkVYct4d6St5a7J7Fz91qx
E0wHXIqpYDUnp3nIUdRHL/6HiPhiUL2Ch2DPmXQAXrlHwKrLViFoZ4auzWgp+HrY9PhTdZRmcztB
o1b3/sLn3lka2936i6QPIvhoMLwUAItC0zDroTk4yPgJIaArkN3+d9v9F4la2XCbde86Aa6OtPX8
9xoWgzcL1nC6x5di0fYqT8aAvFOEbKENjLb+YiFGAWbvKUBDZNWk2SbFw3AVlbSCJrd4Iiu1isJ2
I5riqz8p5+9Rp/9LAc4vdtZQmTmqnlHI/SBrVtXzHGJQTc8j52QsSs6QrnLk0GCGR3lSdY277oLm
bj0CRpwe4dkwIyn6gpEXtNG8tuvJ//fv2JUKr4hy+GLrDDamMPT9mDhVFwZJn7BxQJbE+YeiPWL4
2wim2Ad7/GRXfNhK4CrzHJBrArz+v+X5U4By+UqXI/l+LUw9zG6X/uVw2+9dp0WTJudw4yZipxJk
qpeAghWCXoR0Jt/Twvua+0bbhTC/KJo/AYsiAVXi9aJWkZAHxGYnSWSnUH3otdjLFL0VSSDqoybU
YsG6zm6yjw8LnJsDpGZwmajLLhwTDZOUseUcg83xNnIHeTdfT8qL/BE2gcKui8K/9U4Eka77hUQC
lxihyWCNOqyo1e5i8AemkrVxyBGoW+kS8tU3NByARLoSvNymv3mPe4Jd54msT4D5smzggEpdtygs
6Pq4rr78zHvmW5gTs6GqqCoU513aEz/b1uUDYM/6eCw1Opzx6mtqs2JX8lysPfm644JA9GkE7uxV
PEcBBLZeEhE0YwVIlHormfrzwx/d8mmk1HL6TJohnzVUGhVLDUQndF3HK34bAkW58ifXaQ/o689N
Ajz0oz5XArVKiAf8taNCZVij1fVYXKditVhi47WSf9eeY8l4V2t/dEPhJS7eFKjUGRASEp3UEazz
zfkyXrmA+RUHXFgT5MRSifxzqiBrz3255L99u/y5cOIdvw7+I7sjOfNxXZl622NGjd5Cqqs42FRa
p9CMvVc30gCe46HMe5RUl6JaTdgLnvXNpW9r9zWlkZu9AQj3iPTqBfuALMXdqcKxWCOH3amgbhyJ
F/Iu5dtvlmeY2QKpc0kg5bXHwhQEOwTRmG8bWRMDceHmxeLGAh+Ygc3fBwj0CCIWBPZ7zNtuEcBf
SmIQBReU1jfS49udYP0ttX3vwI/B5qMzG6nFFfvePfJ7s3wcIlJgdQdC90wwN7ZkAzmFlTgWlBxQ
EPPiU+WPi5H9AN9pV03U5lmuqpgvEb7fgPNTHcMDrucPASmLejecQorfI5o2XqbKx+You6QapMeo
13Oo/xc6SceuTuerIVFuOMX/7geIya9qfPhQHtVBB9HyNYgp2/hAP5nQSqZp6rnndxlvbeq8khjg
E21ndAXfGZnE2GmGBJAfOrTE/Y/luaPOxMziwQbfiGGAZqYMvzkr+YO3xd8KMrvQrtTveXqmMI/9
rtmLAGS7dwghUrIvNNMirvLZEZWNKGIBpftKm1PZl1zZ5BUwEwCOMy+sRx3fvivdxZrlehRfUOHg
6WJ/9LTTvcmMvX6UJL0vnJJSIJS11IWvdKbPnDZox+06qvUja36ZAPYTaOVqHiD3z+bl5ExMToGX
wJs47jdV6JWBKSKOSfXpB/O2KQ3US0osXVIV2yPIN7LA3R9967XMcq75NaLlawS34JLBc4Zm3Vim
8Yde9ZL7CwLGhgMoFaSbDYf1z/Sf0olKMAqV09IFgyB4dGPwtbekAR8UEXlK0ZBgu+NsX9vOiv10
49r/EdB7c+UFeoxAFWwSEdFKI47IJqQ9xIfeCNmSupjgb6hXt1XLT4LzhId89/zKHcCTQ2vLfsFp
L6hKzv3Lk9oRWatN58wh6drl0EoyboZno+1KLRqSs1Jibhgbbg+gAYZ3x2keS6/VIFkmL32J/LCe
t9IvZDefj2KbvoFzh+xbF3ZZjpXn1pL5Cr4Ugmb9MhLGRehTwRCsh9aRkEwx1dW90y9fnjyaVRN6
qruvV+t3GS1dU9boFFpH/FDXW5iYag5KL128yHSIlPwbitRjeHm0CVgBt+Ss7cYyW4RVrSnMcfr9
3BH/3zYmaZb2tubyGSieTfQydJDLCeOQd3LsBpynvFz0/0j0uz15NG82C+GmNQz0/hdt7SDqTVYc
29UQmfWrTnsaeiA1otSoYP7DlvMGDKmJZRkRMjNMtyNpfj3+CysQ6EL6+jSBcO4a5DgjLZhvsMlj
GI54rLnA1qGEa1Gsnbun5/hv3eFBSoQ7+Koz9wKkkGo0gD5kd4krrbq58Nb+pH0Eg2gxGGhTHMIF
9VFK6WZlDCyVtA370/tsTli+ljbQ6V54UsG6ri3vM2xX1Rtx9SNdnEcI27fNEk/IF3DbmUzl/XE5
z600gnVoPMrWjk3iGHzzDCjojq5hquu1+pYovkB03OidOi5coak4Fd+jflSQDlJsrw5SAnvW2FWu
k/NsVj5qTCgcYSJNfeoMx0GL9bLw6eDTkTXqob1R8687ZAPqnkMFhvGY+3dbPzBB6JJMtk09vl54
PTWxRQF2YIUAC6PBFq1ghAPbin/fROvYQOK/2E7pCsM9iCx/DeSQ87+UmzVbNMVySRZTWpKVunjl
Fvd5PonBb1QWD9HoyfnFTXRaCi5xadC08GUFXCUGn8iotBfyLsTHUp9NHy1dq808WyNRUgAVB3Gx
G64TyUC0rb7sb1Oy9W5cAcnC2za47jp35UUkSmkP6XiUQz8QcY6RlfhyzdXf10A4RjwtPRQ5y5AG
XRhnB+CewDLMa6ToaeLYz4BxpudlkSaBYj2Co+VSMrddHqKcBaWzR+0ZFan8wWr6AeOhhJok7BFl
3q2EDP/MLWUjsIb22hh2NA0GWlHgUjwv5Fzizdlrgn221NkjlmTe1Vq1wrtq6c3PKBN4c1HbCVYN
q8A2JJATe/OOcMqGdYFVLIbiUrFcRcDc4AiqNM1lDw951C3REKG9n4SlvswHjqfkOST+Rtfda6PG
t7i1OL3ZjcV21EiWAV4X3L95vXZEXwcyxeRb9qxW2XynioYOVk4UzTQgicEnB0w38iu4fCNVpgu8
2+JB94AiS/bhULU6xgF5ltky2Ma5jnExTdPW5h4xLMPnoZYtZ9TA1kTuHYlEMBZpRZS+tVQug8eO
XmRX/KJgMZLiMPIfLiqr5vk9vEV+F4JP8Y3f3ZmjAaW52iCl1jVlKKfZ6i7U6KgSr7Fhhq4u7zix
TqsjFXYJ4g9etxja/RGzf0oT7o2l8jEAqVrZo3N+gx5UK40vR1QIgwdrzH3Vr1RZz73sUIP5xoQF
PHubR6eSgZd4TfYxJuKpN8KJHhQrJfYZbKm0iSCqxbJ31Zd6NWa5ICtYsK4qRp1yzL2QTrpvJvSj
qI1II+G+ShFZ1pmX5BcY+JD3J53pfdgmg1+cw8h5f/zo0KSZhVXEgtbA6OIo3ZZitNSguWocRVEy
7IvoVG6emnlwqHd/WgNzEfHv0e/e8ePV3yOlDgo4o7Q2O6pkWiXQRdObq6UeEk1440bcz2PGjzFa
jwW7WoA0hGTT4wPrGa2KxM7Sb/bqVctN9PC7+kDv995WrAV6vr75k1+VOf+2Z7k+yxQep7ECFPvh
AFGCnfd3f5XMVulh4EIkZxphwCZ5XVxtvzRxTo3v582k+t1nDfjYkI1OOt9xGyqFdMN7kvAe4vF0
lE/NWiLjzvofCkwPtl+/VVp0NYRtWJKsLEuAeTU8aZ1pZfWZBOi/NprkxHoLXhsIM7DPT2RzBG0F
/U/LyOzupYH9evhjW1ifFgBSj+Z0k2E5B9+Xp1Ibu8cmsPG27gq00ziAi7Z/zygFTUd2NcL40vbO
mMj0q8fBAvWy0vCnc8ynJ/ZlO8K8flM1oESIalraeGwPOaNthDmyT92kIu4xX4p3Lzv+RDrI96Hr
wh5sm3wChnhtz7l7N5/hMsYViPfGP5B8QSQZMcgwKozHXqnvhf/sWHe8jpyKyq20SpQp7B3cHcPE
F3LvjYwUQ7EmR85g34yFyg2mn6y3OweXk3Z9V98QPw73qSGZTSkmuIpaI4pDjEXDqw+GMCzGD6Kd
Ws4DSWzeYU+3Q/V24AsM1xGlB1T3GrLgPWGA2LngLmpNKZRdee5vhq57ZB9xcxzQxR/RTggo5zuF
vyR7SzZwnm3LbJALHJRheMt34k+OOg81uUa6Ddo06u58TSm2WYPJ39Fs1Z3B6XCBM+UiHIxoQits
04lDm11KvkrwvtYWKy6ZErX0oUTuD1Fg6FVWA8OdwOEWEQ5liq4zzK5Qad7LygOg54qRhQabdPSN
aYwKZmZI7koVB1+5QusjfB437HTVXkTNMF+SnkL7zbcAU+gRiE8LuBcKFRkuDjhFs+Ffa9mFN/QJ
e7itoRnsO2yHLnoBtlfkU/tUuje/QyouFGQ/Hly4YWqEfYCL8721lvPqLbS1He0V+rPUAT8Kq1/+
o2oZslOEp+uU1EfdLBeOugCVVpzbbcxUEA/qJb1PCYeTDN/9oSv9ljguj8xYcfdptOM7JPaHMgbS
8i0P/Bq4gx4Ol2xpB3gsVC4sZqBw6gTOsyTZrEZGFBg3viMWvD+A9XAOV/dyTT19fTjz3A82dTvV
yXbyACEOu89g/hQEVVEDxOwt5XIfyhJU95DAsMT8/KTL2HJIK37wG/xzHSoQGSPqmkGJtsnicj6w
pENvqKLtWKeIQrjLVn/SW+cXkLSqXanfUNr7si4/MJYQ0MP3+vZH9tecrw7m9HTWXw40qHqq02sC
9/jqJ4YwMt7YQl8tJbTvvE8D3ZHMCfZs+3kkA/rkPUAygOhO99Mc10ixIThVn9b/aRMaQFlN6O+V
C6rPUKCQecjGl87+e5zkAjRQen5zXxongwBb2dtnJgJVBoDbg3YZewK8zyWJefAAWkRYqD/69huy
1VFD0JCotrKHKxBEgvV5KikSu91tRDTOoGBuWyGcydfFB2bc7rpPg5fe6epbGIGihFIKvkmZQV5f
uztmlMQNNjtsEXRl2u0/1Xi12VYZEDJ8yUKVduM6nkbb1xbk8I+obX+N1uDwnQ/sY5uKrMIaanCK
rLgO4ACqyl3CGxr8j9n6O3KPzAH/heeHwV101m+afGYKxgzMTm/RA0MiW05Fi8BfLXNAx3jjZxI/
0w9cqwSbICPX5dy6D/ThrVjlv5gkopMFgK7+z4I4q/r1USjcpVna+F8h6TETQVW92xonuWMCOdtz
FtvdLDTH+GAJZe6QHa2z2HNBTe1YWLERaGNxlRV45eaRFwmOufPCjPM+o8PFWgZ4LR6/94RaslVG
h+OdwWzD2c9ODn8ianu3FrrJFkQXvYm+JjLY5YaTAWR3qtUl2jok1HafgJ+gyl5H0HJB8myVMT62
p0ZcBOivUgk6GEuQ9BgAluSanHdboiYJ2B3a3qZs0kuHEHRp1zbNZ2JQmUb0r043YWQWxH2TizXW
qUqG9e5n/gR7jKzkdSiq2Cow4CDCydRt7zeCgkRuuK9TRhp/0jDvGoo3LWHanXOnQOGjc4hMCXr1
WWBr2YfGSKiEzitSjTqItAwNV/hruW1nXy8UMvPPGl68oZSbD4QNbpaV7+HoAVVvprW5S+30hUvU
xqbUY2yWKvsGS70SCPuRzz1C5aCFIom2BqUrIgUUM1ZDVGp82pXcH8LOYl/KiiSpMj1xqc4eskZQ
yF2E/BKjxpphqqCeTU27cLtGDJ0OMPQuo6vc4q3k/mIAcDzAhZls02P7ZzBHmW1l/JHLxMA/tVYg
dN0Ui3YCYvdld1HFJ69jSdmePtS7TWqWoafzh5enDS1TRuM1K1gvBZy3JOcn6olgb/A1bzBub3yS
rjAnOgXHJak+LGJVqcZGmhJJOP4oIK9w9JG4vV4FnQ7YDvoarpZplXAPBJhjP4YAWAFPBJJVZgHB
KyXYDCvTKjAZJOrbnTmyOPolIgZ12/kqmJzCdb1tTymkcWGOsHT53VoQGSKEaUp1zMaViaoFzK8Z
/6MbBcmh3QpF8moTkIY+eKz9wX4unTzDyWGh/uNg05fbnfjhPwCnASMiQMAdnJuaVZL/G22Ggy2F
O3AKx2tThpj2KLx2p7m9B8bXExQkrhRP440mLIaknnUKXMrryO9kCdD9XkU1z4tRDIAl1LoNIGg3
EL3hRaLLfjF+Q1B1n1D54IYSD8jAF7AQr3xkbRJiNjOn0b8Uhc6U+O2kZjtsmxYfR9oxJFSzk1yB
+BTcCq88pvJ3FNGpSQQkAKELQ/FjW2zapFnABZf5uub/jDAbyu4nW1wd1iwTZgYQodjOtvS8Bjb1
rbVUJ0ulDp47BEINxX14uE70GDa/dUOBnlPGpEJgcFEGKj5sUGNWrVs5xMqHU/NFce0B8zHM8G5J
5xX7kidr1YJVodDSFN4CcgbwlQE2GzHAJX6RSyOECZrxKRh5ztiolF9NhFzrmWibxufLN+TQEh4t
+GBFsfpkaiT7gFj0hUcCc07LSOoKL5h701Ch/0PJmKeiIuxOqfw5toTYGkIjljVBE9cYbzO3s2RZ
MuPxnusx8uuZN8aU7ttKjDfUVxwKLrwW1GmE0Vf2vIafbcLPffMVb+6HfyNsU6FCdrpqR4Jq1EcC
9NV5FU+XIM/aqZEj8DUff6X9kl4QjbPSLWdzm8vum0c+7ob2dJxbHaIZJOMdX509KbHtFPojpM1D
DzSpmQvtuGmIEY5kY5XnssRnyA3reHM4XCHEVXqJ6CsBXGG98sYugrF+sbjH8q5joNdqmbn1yNGe
N6wEK0J0RUM+aECAyXKRKQYi5d3c6topCkrR6in3QkcR9tpmYkBNiFHyNK4FEovNG4uE0llcmJ/u
Qe7mIdTbqlA/4yu5kFjHi26AMR1Ysfj0Xu93ANb44IMw1dpqIN0n8Z6cIn9nzlnvXiKslYkJZ6Tu
iR/Yrkcst4aEe2eAwVtii5Ocbrjn5EgZRC480oCDfwdkH8BA2Ewt+cuYUhjsUps4PALsdhJy5a8w
3sBA/kXnO4z2asYFcb2K3FC8M6N8/9mZOpEKbW9CKBkJm1i6WZSYBhD4EYwZmauVz78wHUjGC8S8
Oxtaz2Nant4yT3U7bYiimOgh0eV/axI5oRJjHK0r60OdbK7B8f+nbMiXIeMQUiG85pqoNn8j9USw
hCEFUcUz2jpkHVlWjWLoULsJWe/GR4jmoBHg+mlwMoVfzd3FuDpsb4biDK9/7hwS/3ZetpW8r1XP
EAcaDmFlrbrsdxAfo3T6p0LoOtOCs/Ol+TddQMxooNaTalUetKsPe9i5yjXvTdlNc9fyqUVnT6ay
aHM9V7mseRbHUqD7lKJn97HTcHlgJkER3RCv3J3r7xSd4MXvEnia0hcpatx9uiPUNq/Sn0fz2QhN
2fOS2v+jJaQDdDni3w/rqvJKmH75S5+RsuDlQj2iMFFDwFMRQd65cUqLxmdhND11Pkr6Ij6OeLyE
Yn9ibP0bAiIpcPYBEhjCbnwjC6GQeU2EETv2Uv4V55bkALXP9Rm3j7GvpP3DgxB+8b6YJI27EDCa
+SOfRwyTGah7yYxBJ/DWeZR9r+sVdTbLzT/9jYBWT5t4GQQXgAnGX1nbBOG15gChOl3venvx8ZKJ
CLN952ZjcQJxX1Jxm9kKtxUDOMredCE5+O3UvbjGwxbZZg0Vpp942kqETB6AVaoBx32cdR8lUL1+
k4DFXyHqiFB1yR6E0yL00hyJjd2lMfwhQxwBJYGNRdELGNQuTsU9qCmCCt6rIDIWu3MvI11ovvyh
LCFXA68ihl1HRwmsbpb5gcIQG02S7LcekTWowBYXEj5thQUOWIsvJXJo9SOmxGL45zdVC7LAmstg
fqQWqFgsGoakG/O33jBwhykGd38qbuVyw+W9p6iWohIV35pPTffLgYd9sv3nGu4NJdc8nWutJ42/
+rQD+YCvwOJXEFL0bI7yrhkMC4cXj526XY/o22lLPBa8GrgwWmlW7/EkuJZrcc8cvOwlABKg4DjA
Xfy1Cve5eW0dB3Sg7qSpXGdZdXfiRYdAVLw6k9oKXzX8Zz1didO1RiVDklYgOvKCfI8n8g2kvM2M
PtKRs2k2RvUy7gQmiSE2izyjgbaUuCDVD5x32B5pK1rZFWBTyC5gTwLzrSv9KGnNDHlCH23E0Xm1
I+BZ7TEER3qjsyQ08RBCcifsTUhjCEnLWNvRfytV+Hk5xDEeH23sI9IXvakN/h5NEA8iNzXGUnTj
cwcu7ionDen68Ws+pqjvxLhrSeCIVEr3zJiR4iC+nez87PrDI3YGdcLrgZusTXWldpndV+pWyYDq
07qTMvomvas86kiouhFW5wQcl/mPuA8KVKV/ryf2T+TsIvxFU+T7KbwTStYWOmW1K2B8eqNBe7CD
hZ2NaQ0mngElBkxieyM+AXu97ec2IFRzVDChE12HpBGy72uSEkkVYjWXJXmazqkgP3D/EKfK3+qN
GWJyJOEJw0zLChMrLKn5zNs4iC5mlkkE04ZHdiro0wpDPkoMOL/dova3afBpAoMX5cZGr2DVR2AO
WUZpV4m6e+OGRDOF0pbb1TUwzG2etHYWeoIdVIwZlUE5425BYuCn5L7vyPFif6lW4Xm4CHcs1UHM
LM7iahotkLwjfKYwH8MGXZdV3Cl9NmnW8JICoUM7+O+yBKQQ6olr9n9hvYZHxDJKgKOjOFmPIMgx
xbJRseMKXuVlvgANTxRBodSUXEi3VigRPSJasNz1AZIuq4f+wrx3pnTe4nKDHhiRlkMWApZE3GZp
JrsPu/ACubfZSQTTBM8vzksVHj8zx5Nj0y7fY3lzZtGAtCm9BlCBI+WNTyYIY2ujYVCMkWoqqvTv
/ZIVS/mgylLUdskHyYNgQk/O/WJyNdneNsT/mqc/OMnTY0wNMNqgDIMe6hHS/AkFzdz3AHIpYIDX
NVqncWC4x4eCqdWcd80xLma5ypOYBzESFljFG06vMN4qQLNdYzfRLqAASg5Sr/n0WWqlXHXFsDbt
Dmu5F7dolI1eaxx4ohU2rIg5m3FLzhmmd8lim766ubw7+rOPJ39DriA2oe5nRTyR8NP0HpHqv9kN
CqpyCcF5xEHuGXHYhBDHpNBEg8CBNIYLYlWRCkBxucpf6Z+hI2otUlSCEGDBIZJKMLMbYNsofy+X
fu0702az6KIKLC0rBNs76CmyfcnbwoRX0Ae18/Sgi1XcuE+vCxdAroYE8H/cjxbL3bPeNsTE1h/7
QqBYQPkNFhADeIhEZUzepziOI/1HTAD86lA8sz88IFxYkuaP9lwyWnc+XftDF8+iDlQILVW9WSa5
t/8zdvruS4SDNNbyasKLZPNRUypTZ2ihvhPfmwW2v7MC+gGPDYbsD8JsfTCQbnaF2/WVgYdC3zBq
zDZgNAuD8Kut2KAs8cTtogcRc7SA9IVpW0vpqm1XO+8kWyh6fiDCTWGrNsSw+hY/FlMSUhkuudX/
WJtn8BaNdAWk3hohX5NSCVUHr1q9TnnYsikdAo5jvJhgnU38IsPU022bM/BP+jn2C+oZvLgvaCkF
xHHY6KxDPFV8IOxpSYeBMs+TAysAl5Xhuz2WqYPenqRQXb4fSje74rDVIrCIdk9TSWmLjPIjHUaP
JDO72A72AXC89FXfnnGSg9UNg7QSsd1EoecdmQIjyZOKf33vq5bwqs7TTGl3vaCgYgwyBAQuy3io
Cne5JbRbqfqhKeHqhiGx3NljTGK4Md3FWufgK5OB45nTdRaFkAdifrny/cMiT6d4wiFaQinS+bdM
mZLVjxHuvg98IB8k039HtGDviOCaJnXIB9h01lGFG6AzSvDp6qaajgXgjR+XzXM2Nuu12FcZQgl9
LmJkqdAsgOTAxddhZ4pQVwENtPwyQWMcUOTlkqw0wXkwHbyI+XfwNRZvAjM03aXNdISzQvIOZrW6
J6l8/XFkY5CAtIlcPv8u8/mLwUJT9O6RwlBcDIDEL1sNWIFnnmE2wKvn2F+n23XBfQoHUVi1ce3K
0/MKLLPwIix8eSpY+mn8/by4TUCUOYwTL7QcgFmF5pfbbhOCcvEPO5oSxr/mNiXLZRkY2k7qK/Um
YyGJ4n+yESai50seUvzJK/3gnu4f9W22EvAx5gzNuVb+R3ESniw7eFTtV+B1pkCDJRC77Byme158
+EhJ336G6N+RkuRuie9SWtXvbemuLn4ttOMpiemEpFow9GWdiZky6zAiAw2JZuG5z75jcd4ysdxX
WMO4BNkJXRHq37ZWt1loAHxbjemD1bah9wC8i4WlOuiBYuA4eVOIY1tS/iSPAmFJcvWkyKKH0I28
IkrkHWRvMt/VxIYST2YDVXK7YpqZw6+t8HwPuyOmIbWev6XCSEmIHuzq/20oNOtI/bQjh8pq/8dP
xNSKKSx991zOzcqBqyn49gI84t9Y6OUjD5ts7D5HDmIQgYZav0nxCxzOVsIIgIMK75PqPHQCriwG
2ton8/tzwAvRrk2yetJzN5FLQaUlbKJ1PSVkm+/YyqpnvcN4s7MOoJvBacU1FM+UZcqQ+4ck/Xxr
NEt3O1C9kxyJxGiEKVUmtK3j5I/JYS/g8jgQmhkOhqnuZQcm2SZ4d54NI1d4LA3A13UuYzoCusfJ
6bB4Ofummze5CwG+tCy73VOMn3IzQY3DhJnfG5pk5vygdtER/buJlWZMXSDtmOfaQ+MhHqKnyfTu
z/RggdvIAHWzdeH/XhdNU9xNzlpaPEb3BMuDr45mIQkdAzFHwq9/bQtuSIMdJtmEn3h03RnIsaF0
H5inP+2619zaJ2n1W3M2ZF0cPbtr8eZlMcQvb/H+CY4Zw45HrDOWEcI8HjF4mOPoHBsMujgoyuse
d59No+D13JfJ9zYoejdgjpN8n5zuyukWgzRbPdwBAPzTxFG2OrWM6IMp0veSUSsyURFUFl0L0tNg
qbggJ9kTsx9vPLRal4LYc6cgA3XDaCsUDqNBMaUgjlzplQyMF7XKoSovkwbedxMiG+RpsDcpgGyl
FjunH3BQ/wYcI9AP8MqbLtb26YBbqiJ2uZfmojClVJwT45Rw59GHJMZoYIRdG8YeTJRnOURNLNpv
shW8/erv9RvmySgGXzuHXlxasd4fThOupXCKuAPMWdz/dLZ1+nAYGfkU+f6b4V9dSCb6JsfU1BeQ
XYFDvgq2YcZDYqkIzyxBOCTiOF5pDYc6oCo1qFnayJjTQRCV4bjdDSagGzVzPm1G49sEkODMb/PT
KCiDCf8Jc/R/fKzXlYgVT/xKcOJk0Y+T8LeqfiZEYHRY64imgeduM7tm11xu58cuPJ1ppy/pqcDI
9ogy3j6Y+ek9J2mKwBf90UA5ge4bAJ/kFfVyWggftceNcKdKZ9AztQNqgix/8nIV0sAvqLzPIZVx
2naVZwRA902A+9Dee1T6pjGZrOdvR8T+RGNsexR70dgODztJ5qor7QLADtEj78D+kNGcCdIWw+b/
t1w/rkNefXqmHkkwckuixnyZS+9XIxOcX7QukOo2WnNQfKyO10ZWJGZ8e6CXb79j6Q8CXK3IJYaX
tuklRrcYWIQtdeeLh216a1BVuW1GUI3V6GPo26Rd1g20yWKGRnQAu+0iBNMC9upjw4cDSW7wihp1
ouFhS8Ttml56CITglaacS/Z5g4YMBtNNKRTac88pAIv3y+iAKDqaWmH6Zez3GLK07mBR1CMryVjr
gDiBUJZAqiAp8542Shvb+hK25T4Qngn1KisltsNd9FlSlc5IfuudF6HjkiH/RssIe5Z6RweGzbGk
W6KwxiDQl6PASGrmwErHNkVYd0XtU14uHYlp/W/5CYyYYlI18XRjhACjYofTEmnCWrTs9oPq18LT
bjoLpYG4DiK4pOr1yn+ln1LQXBC/4ncaFIlTtVEwV6ER1h+3JHBdncjM6r/RpS6ZNF+K79NLS9GC
ohhHM75tjXvEao0vIp/vd66nUwIDg5UAFDc9TAbj/fs1zcLC0J8zuoRITctPrvAYPdyL1BStlwaV
hS/cJfAFPRxkYWAMEz0kzBm/s8bxUNmJvNsqs0mASOzeJBifltxWWY/jZ1wXUpxnLAsSEtMQqlUs
0rNqhPT9MLQ7XUsKBJJKpT322vHlQp9Zq3qeabcLvfcLZCLMm4HgWpSHGTeBMKcY40jdvMgZ6Xw3
b0kCCJzZjj2nfNZpiE82mUiEQDw1hYvD24S0I9tfEPZG6itp7/ccd/TDjDjuzPMUncP6ASPnquBr
z2TT8msB+pXNplLry11efWSSsHRGpjYE7tHc85Zl96dXBJlmsYI6roYsoBw08fAWpmYl4mH6g/xx
xzJiKFC94Ql7k+HQyrS9VD14+WAUMtlEakGKdGPhbDF7AqR248MP7PHrcrQg93ZhoXhUDMOk5NL7
oetzJ2iqc4HYA5MB5B9RW0walRinYmoRb697mdVAyc3W34rPA9AlBVtmtvzqAIw4mGAOb3E0wOor
ZxHYOm7xQIzRvw35FTat1aW2c9FCxx9S1OOXxJXoqrNU6X5FC/W0GvcXjmFaqzs26nyrHkBwA55t
S08dTuaYC0PDWRqtMvYyzVrMy2dYFXykcrRw2PDohlv3+gLJBwFIO2NmTVuqQLK4W3I7bJKcp0Tq
LpRsPabMF5sUNrh2KpzWwyzLUZNHjf1DeeWxww5n4ooy48V+F0tE6Hq5SXvnSyZp1VWB376zJdCQ
FecCXbDaVI4RfpJPwaGSYlaqRCC2dS+dCgx6oiCbOrz6yQMjQpHxMkmiyxXg+KQJzmSNxGjl80Bh
O5oQ6ipjr/J7MAdCPM9Nk7srb5eqAovWrOFUhccgA2Sgqaj0nkgwQT2RqKG80mrRVztgpeVB+FmY
uYiRQgETiJbH9IrhK4ny2CI99MD4EMqWPHpHkmIHY79bvc9yiyeoUWlFPaKSES9weShP2DMPRug7
NlmMNWDm71KBgHJylh5pBg+GwsDCORhTDHjyaEVx0/LNVVHWSbJAXNREUwoUwIGxLAD50Kf5NqpE
hpHUusba4AmhNjSIHvISp8q597XvlTNxQhaz7GjSKCUsDxm6d6j2enTQNDyRvMrV0Bq3nYfJlqE6
AZnZIwxdiatFJRU/MKh0i7YTdnBb6F7Ql/qlgXRFC//RQsXRA38JxeZO+6Jh6RDpAmWbiu6Sv4if
VS1HF5yd2LkgmeqALpmMHXNB4bRo1U+grI+1aQ+9iMqsuzXgwTIrTJHTAVcc2qYw8c7JHTAm6xWB
/YqxYpMtUDEQOKJromw9GQ+ZlR+xDiwi5xx7RIiv8iiOqNTUdVjJ2uXwFI1CfXNiWoYxPdLbvS55
9iw04QUSbGQVpHQQso0SmYhwB0bmLoyDZ/TGq3B/TUjuGH3axHxeqEjZ89AK8JLXY/0fGmckC6lz
Y2xqtIKc5YQMUbO5y5RAz6wmTGrXFf+pQVzSFwpfQdiASBdinSyrDzQZx6p9ab3tOa5Jjme3nmZg
gVoZMuy6+94fvSp9F/2K1/SoXZEU1/zSr4gILMahqBg0AypZeHu+FuvGN8aDPY3Wbqk1trywl4fh
XlALJbop7iQ/h8NzIRwJ3G5vaU0UsXluBemT4V3yY3efYFgQIOMprmwdwJuyJhPvdHDDWmA/aThn
Au2LC5zmlQX9oOqmz6NujP0kwH24+cLhfQ0Ix4GqHS3FZiiNyJjJ2mdZPnlTlrISEbMyGxqDe0H8
ZrjH7WC+Ll811iBz8+TX+19wkKGZp8KoIRW46ojDh9nSw3+ZMkN9dCnJ9RbPi/UYmM0ll3aA8FQl
CXCCxZUmbtvO3/aQJGA3AFrsuPEA6fzpPhMiCybHmpAFcSqUqx8jIa2fuDDK51QlTdtxfmqAMpnz
FMeyFbpw96gtMhZhPB1QtjfpSdrdquXHqZrp9ElMGqSjwQoWFtHAolgdo85cgbzwNLAnvPPUa4dT
Fqj3H8W+6PnWaiDgUV3A87JV/Rx3HiosT0q03Ou+cFXe2Ilf0ecCN3xCn+ARQ1mPx3dwhpCioGdD
bLaYTWpFBz76EHlwqqdHdGEu9HKqr4N6cpA7bpKWRtsyje+Q24KxHql4B+1iKJMwLwiJJWeCxIfE
6/XKMdmLtP9Yq6Xlc0JCd3uh760TVslvsZlvgFi1DSZxwI4jXYr4OZrEAjsHtzFQ3J5IxObCuV95
Z2uQrKFH81jibndFvy7DiLuyF37HIkRP6wJOEDluYh+yQjd0r34qXAB9rpZ1ervQPEBhyll4Vs3R
BAvtsQ4CfCnFXfpHZggBwZWdRe1ghyN2urFYDPWvcflzi8IH8FnwRfsUnw7ag6BgtUSNGkiyHvQm
VfPuha5RVS7Y4/F9BVYy5FQiRfHZ3NUrEvC/A/cJGM0ATxtAk/HGfHlwEdHtyBm7YXmmfooIHNWu
i9zAxRqSNaB9XCqpMfZ8DFGq6wAxNZ/IVB7l4moe70PBzEsZmQB7bLs3Y3icbVGf6PNeCpBFuQ9T
2hlEL8yt63XcMs56OtUHGaIred0pe5c0yXcVwZqvnoRqoNRHRaoTNJu14oPuBX+gawhxyGx4Q/nQ
BcUlhIWLBYSrT3wCtvme1hjFJKdZYv/jSDp8Tj4hPfhqU95sCCM13u21/DKQX/UL0hhOxAgdAfU1
60NC0N560U/SPMx23D6WTGGuBwandpttlxYVTzDwGM05A5+5kP0n46hnWFP2Z6IUeRzuRxO5VlVq
GjsPJ0aLYI1ELZFqn4G7sv/yvxUzXPfrdQk+bZFfD9E/toUjk83QYAmQ9XhbAPLP2jzLEt0nqyAg
rzvmaZbUp7WEX1cC75cxBpxjz7XhuEUGUGhNMf/LEyvjf74jH7t+KABZnyhtB4jufvW1gHTFdrvR
pyy6lHWPc3iTsAL0e0Pz2hLl8emtKHuOMakidQp2tKY9Mw7NlQXEB5RRwMQvStagwSN7/Nfljxre
58eWMJ3jBW+0KVQyHRprtiqtDno590ULOqdmqgClf7XzQeq8hNqDzMirYd4+UcHU9tzdAqUgA0V7
whnVv2Im8ggz7QF13AF10agY6nWnPEvf72YzcFePNblfzJQ6ageD+13o1NEUz7kd4TCrfNRuE/yN
4iN7UpCQjVTIKT/OTNEdy0qixQixiiVltuwAJcXNpqzKzJxPvCQHQeArOeYEC2qlf/YcvD2ZB6g/
nimwo6fCaB/ADCmqZJ0rqwb0wXwF7QobE24NMbnJncpULnuL2FnupXO679bCf1usOUeIMX6pp4d/
RGxDMigimCNU3+HeUxYuA8f3XayPklm/rkyTZR3d1aIe4jOzJM0SouKWoChi7etHrurs3OgIR785
YjTRHn+3nnqMPy4UN/XkgCHkElWl40QRxhW3shQ2ujfZazrd07qFKQ/2vBXHqD0cWMuHiNy+1gJ2
eiYncUQIdyT5SQYcm7/NxxpwzOC+igOe3ZekIYNasyAZMF7i8cbSjL58B5/I5GhMHwNp20Hlj1W9
xbJAMy9/5p3Y+zaiUUOoOLD7sl3VnRMTbIynMeUkdLoHe00AYuVXda536qxvZ/NQ3SSKocCgftXI
9STfm3F04EiMS0k0mLujNeAWH5F85s8t4GRT/pIkmSudmNWQC9DdWRa2KTYI7PUm05022e2EK1mR
kQzG4mXB92B3e3Z3RMVRP0uvQ1GkJrndrMIYduwyO37w6WbBc+HB3h7IX6EnRM8S3od6v3EG5Zc4
zgVgdFfYOTo+kkqGKuOpKUUL5BSkwF7uY8RnosoJwkS3i2DAQX1oDwhWEeSugCbI82hyMSh2ysV9
Ozz8c7knKwNcv+YFrI4KTfn3t4uj0IV1oK+hGnRSSTN6o8i+GUJqPKIo4+4oORtQDtZEECQJBVVN
1YgpZfrSBAmsXrAj0/Cqjq+vwd5QjdDKGnPE00VW9OzST9/kRadcniwCHc62t6U599FKBybxGCnd
j0T0PL85e6bnh+eEOT329PyrgUxbG+3hahZ+ARhJWfHrng6wYAE9LszARa7fXyY3O6v9D3CbwReM
nfZ+D6fCZwGQgd7Nd30NCCvYaz365cuq8uN3dNzSYzinNVY80kG4KgvSlto6aYzmyxNIKMq45dJv
0G126GDUAHLT50zfI69Svz6WKRb06oFFcLi1sBYql1h1l3DqLd/yJzuD6og051jrwgBkVLf57lXG
aBonPszzwsZ/o4GOxtz1KrxxIbvn/K1Qxs+c8vybJNqVg3KGlotYIwqciazT1oUlNqiuhBnS11kK
SvywVHfQVHhhhdt40w7t1O2q6sXKJJ/AZ+1vahz7d7sGVGXL0Yar2GJOZ/PopzzcU9gE5UgqMBqk
99yrBdTqbFbZ5fyrdxZT+MBzYLwfzIhYYRVm99Yed/tVIuvv7pmn2+OHPva46nXHuaSnpvcUC7uc
nsy8dudRAUQ3na9kIqKWrnOfl7RTy7ZXNS++rNIDMUP1jABmWmr9VwOC1IW99UDb4e8+/LEJ0Y2o
6C1bk83FtV/xzbMFgc3ifaGxb3o4b6lreyKpOlh6Gct9CI3DDa9iPGeSc8UEA66Jcu2V+xPmefJE
bLxSrULNXR3KuI6CKF0nuQOYqvZsZOcoi/c5RnPqeEG1wLVoVGDceuj7O2Qjd3Aydh3fUa3Zy4cD
TZyKU7R4q7fqr1UsCgwdV3mM8e9k+MunZaflYbQV/FKMPg2KYWHaU32S7S3j9emoPD9Es/saCWCe
8+DKuaBopOa+auBWY1f4+hF7fIR/mLgNfOtSWS8su/1hI9HSKVqAUeApGg2eMmuY5OFzRhgIrKza
KkiSdIyoRPcyQQflnZRn93fBeXCZF++9LL0mPvTlrMx/iihZQu7ebNbPwN7JhYOmnTWOc9je59xL
IRDw66ly/4zrqTjqa+XqSy/jYC9eK2KrqPFVvT2QJcYpjy66gUDP3dgtmzhJ7gqwiWLe24Fs3mpA
kcJD4SdIEjug2Gw7gOd9CDmn5vnxXVNJ94uqVFdl8NlGccrC84ZZ5Bpda6COQKmY2/fvx4MZHrH0
MbcUaIBadiacxh3lsn8CvhsJ0i/50icuVnc5XwvxOhp/4PYmn5V8CjEcWhgOzM6HXkMZCOGIuxZM
h1v2QGe/rL8rWN5b3pgAn8wQdoy4ZEhAl0cNpaA0MQplpfoHyCl2WEvlGFQQneA4n468uPtTGVD1
tl/Ivu6XyzCRKjDxvyNaNIYPflF9C4SY/xSXoJbylFLIRXs080+61br/7/Mev6fiL3djCWrkjKcR
sdEwc1/MyY9pWxgDicTur1nbaiydH/ANUcXslUuP4XOlb2sN6uKLDVHztYci9mh+MuhrzsjaZ0lK
TSQzLwpF5PpVK3TIap/54Iw755Sji33cYvBfthc9v194TzOKjng4aBBTC7puJGBOj8rf3VdU7hC8
gP0Ckxsrf7QozjFmG8L81eUvNri32EBZqE2YGK+CNNtQiDnUceE7lVv+mQ0fsY9LbPzIXvxec9mD
tlb1c3FkC1wJozu9zP6qWXgLNrDxpXruYWZdg9vgYCC06aWLfyIxnQnLCkwtGWdiKxnuR1i+wDL2
d4kMa/OITJzFdnVyOKWRJayse/vVfysRLPSZx4+vxCbB/IrmvwjQ5Oychlfs/wTaji1GS7rvFjok
vn+y7Dq2FMTF76srmexipiCn4GrnrlKcj2iS0cnQdPNeSk/m8DKYazaEABQjouJA0JU/CH5yvl/2
W8h1C9GLhHj1bAtkEhwhyBgnyukG2SWa4rUCjnqgTiNfHRq+Kf7cy62b00MOabmwo7PjL+V8/1sH
1f01O4faClMCvhQ2YbV5r+rkR1LOp+zboqTqlNioD/6O5hY60NIcKQRGAODCl8/bWpxaHHVI5bku
HppxM3BrHpYaooyBWNgsY91jLjaMouoWOZl9YgXiFBN2Znx1JVlW34P0JX9ESzI80Yie+QFzzAa/
NrqHT1O370YmfsdP/v9RclGaLhcVCawvQLrIMgVIm6wo+ZjDDKmoPM0sIVOGMSczbYJRQHThDzaP
GrFe5RE9XUubo530TFFsCM8BVtF5mQFYAOu7ch/EVu7p568HfBUcIZJCrfHkRRd3izAyI1IOhBt/
isCcyTAM44Tgd5skZ3g5ButSUqDe0f2wQEhPdGmojR7oid98I/vn6XQLkDNcTsPMZqtH4T/mVpAA
gb7ibYXZEu7QXZKaSg36lMlIW4GXZwHFdeTxH8OfpnP0z9E3IoTaodS0+Y+0YL7KJbHztzcPilCh
e3lLjSQX9NumozuRvzViv4LcDmCzOPzBPIYktfTyJfN2aU34wE3sieTeYvNC5cyMuoOM7KioKShD
QgdgCjY3n0RHl0Y2hHjtr197CdyTv+aK1DtAuOouG590eM9lDdOm3/xhHIjtmaOwNS6KjMh7XUab
WPGeyHQdFtJ2tHC3qaVMwcKzJGPkJu70keqKgd2UVn66NHwJhl4PrGKJoHbEyD+T3FS6xA3513tq
2ZqF2rDQKjQB4Hvc/oWEoE4JsJW3X03kc4htDkVvDZjWg61M5VhKXWYhO0CE5OMV7rKs3zPPPWLV
a5CbZaveFLe+ishy7Bj4pLlraBGPO4/ceHjJlfv3G/Awsfvzp88wWjmyfLmk02rvut4QJgjQsiAG
B9ZsAS6Bth3qHQx+FgueWf9ngtWtDFdXux1tvVxtb8Gxty05TGfyhJJ0DAR+A3Dy36VWnh5A/+Gm
KU4zHSxdJ20RyCVHPtUYwzc0OH2IwuUMtpwajVj69Yq7tvI9GIW03YE1OwZtUTKT/mc/McpVMiXx
ecPaZVP9rL0ke4eZ9jTYGEENg+LsEyU5rJ8thQwJqaMF13MH16vqnT+4v7v1L4sG8nQXK5NtUu7R
+RiUhMKeUdXAwDsOv8eS2EjtGFQS28VU/Y+70nAnYHfumuk6FuKeBWQvKAIpwv7vT+MOOZVDP2AB
IjqMMS4QuQ4lS2hmL9a6BYKlZUSlUfwb5QfGIxCmvE+pBfQXl5fwvOCH2klhRH8jF+098zEdPnMf
SwB2LBXGxQkbqaoUY3Y/zDnFM0DSp36wO0V364CmNM1d7FZGXJscjZ9xuAzc4aiCxWtIn4bYRGeO
4i6U9xqvZVbKhIF6X0GcEHT/1NLFMd4V1HuITbEFrc6j2Vc3L/riSfBL0nVunYroUxqrrft4DzGK
xq6XyvovfsWjTmO+lUdaCFFvU/yMQFMRoPxpapiQCU4Epu5A+vKRHb3ZagGeKOj00ZKED5Fx/IB1
Ti2j/Dbc5B6pgyrnhbsqD5IKA9cofiMcdnYMyBlYVppFgLO8/8li+i5xQRpyUmSIIrnJbCNuZeyt
K3vpAU7RBU5OsMqEY1W49d+cGujRzHLtUVg4z2UDYYcRMiG3soW73Vu3W76KowsaVq7q5wsSnna5
nQ6wBYJO+dZUDOGotqZUjj+EMv9o90BCkOAs4lBJxI7WdDdWCj2qxKJw3xHPaNsnpciDhfLAFgfm
Z4vwZbxM4zk3rcY6lg7ITW1fpmmIuqeISSaMw1cTU5OKuPRYqeX+cl6FyUYbTJdrSk0+/st3P4gk
AcTG/Xgc7yyPHfS+gbMZKAJpEVj8JHLmT9MVh7SkcYqMxt/4+rsR+DUDcDJtxxSZDJfIPONGfNX/
a1t3llBw7DoziRx4UQtcR3LpW//EuhbWdZKTUWbUxSKP03S+DhM4hIOSuzWX0DccAgcdeTgHelel
QRuL3Z0sAKmGyy4+YdwHf5e/P9xv590215MGpRYhBT0+S/2ua952GO3v8T8O/hAyerbyELhGH7e3
bihPoOtmiCT4L6H+8i4IctYLh4u6aZSTkTi+5dgh5BSrbGsjc2lre8zbNsjC8/it47BIImeDvXEh
LRny2vYCYqAqFADcd5qpEonJQOnbwVXqlCG1VJKD6YTgQF+uwuHnKRFJ92G1gGgb9upFEiHWHBo6
or2kI3G1NEjJJ9Ja32e+VVFqerHm/S+dEcaJEOUrDAy4Ft9fCCxUM8lpfw1+R0QEeaPbvHafBgIs
Y/KvM/BEYQNaX8AoEjRCB+J0Qq1cPFF4S/oiP3Em+JM3jOgo2WemtfFFv1vpZQDuEg27XES3238c
MCy33QSKRt2DTsjtwQiPMZ1VrZ28rBqU40E5pPeRd6mq98fNANJKlfSwO3t/erPqZnxHmIbTFXh2
oF2N0SGkGgpGUxnxmcW/nYhrothkDuN7bczhXOwuO2A+LQVmWHBL4P7Mfx3cvf/D2NTgid0QP5kz
mvfkA8K5xxoeVw/I35AhOyIoRaTIq0vMelv2hN91rS4H+QbAgWwKK2X0zlhJl0jDPjEHf7PJxAf8
M0x67nMbJ5mth0ZlW4ZhvsriJvQZQloxnBtuSmEMIjbxeUZ4iMU7YIdFRzufWMT737Yd/f55lPUp
uLO6aPhuqHyroh1w6FtgwJ0bhGDkv98J3tqTo5FP6mC54IFUep2I2tia1mDNUG29a1s/g7hPU7u5
ZggdjASgNNSGtbGXsVXk6lgerR3Z6lLgGTlCIHzUreAsuP3lcKZxQdeB1vBxWsyinsop+0PhFo5t
nBVKB4stIRihp4U+L05k2B2RfQ/G3cUvEw3pWYlab7RVGNE+QG6vBYnnzn8lintI6LXL1tpx7u/P
KE/CX7T9+iEy0s78zL4J57umJm+WEKw45i4JNsv5lknL+02OvSQ1oM5940pbf5D4bcLTdgGOOHQa
EedVjfTwxbYBy1R95xRUCjAsJECgdLAsKUWVRT2nThGioh1CwIoVKKQYronuwdj+bcD0lNH9hg9v
hfk0IeBZQ0+GKvJdBCg0a/m8vQ+xbxJ3SCnwPnbgfVqcqcS8dZPGP2tuo+p2jmunKCowEayh1tE8
98nDFjP/gpSZ97ucNuw1OzFU6FUNoBTuyZUEybaMwCRU/AsioSCNNszPlhGJncTIdvIXWF7sxVcW
ZsfqZFaJ4AsT+ESOboCwPL+wzO6tItkPunfPWiXmuNr8LYu8B+AYFM6uNkHBPQSMD1nVSgCZhNrY
wXsYtEjqSV234IL0wI95Zf0Qv4+4AGy61qRhWYwLaz6/dhVKCYFMHgUtigyb5f/+zb7C/W7KDm99
gIn2K5kmyQEVPUQus5jo5P76G50M69iPKot2RMxITvGzaSXGx6SlRpFM2Tx0ztMNHScKJKfQcHmK
L+AuXti1vQNJra1WV2OyrDthoqKddL3NIwMXBFxLlWICySbhYzagA5viwXiGejPknISfvIeAlY6I
QkZ77x7z7nHWlsZI5j/kIEwveR5D6YJd7GASiFgG5Kow6Yjk5S4v8co6xNXCAURNkf9vzP2nVosq
mXV+hsQK23uTNAjCQUnz7LAa80Hpv48uuzzpfeVRWNxB64r+BfhO4oNl1+WPeGUCPn+qalaTH9oq
NjT4gOqBhpYasjtLXSMx+GVo7dhwPcBjK+F7cbhE92wjiteWJ2P9pjJMi4m1WLTf3dmyCbeoDceJ
nZ5SSVt+6K02XN+BEBhotbaNoeI3vad/Om1M1Z9tVygBChiEU5TtAFZs3bMQ/15XwMDq7AleDhLa
higyQ6vqKFDWyu3OmkUlMk1phL5/DU7qE/4za6YZwS/B5iKPAG8tAF7A1yYQsQKgKDpOPtnNMLx0
FdzyLjTaU+ddCyhwCCQqNQxpZ4qwq6NI/PyF5HgD4Hxpn6aATT3NxQtfUpDXN1UuqJTTN3eh6Jnq
7R1MsvREycp9Qe/WoDOI5J1e8Fj07gR0UGnDylTFapISQYIzrTS2eLhv4pytWOIiuf+UPsAf1SlH
cgUwBC3iTn/aeVAbJNH7ItR0vCoyyit3MciAhUgEu/Dcg+ca4YfGDHGzEo5th/H90kVs5wKmCLaO
PI5zUHaXEex515Jht8XUkBQNd74vHwPSZZ5jOm5SO8eCM0UpXU5/TTusV7zaEUmKldpZUPTtPKOP
0gopW3nHbXxaamclyYJ2nRF7zN3hJ3n6ql8FOsDoTzaQfajScJ4N2yatulCAARUSLTJUa1f3rn/2
Fagzfe96OHlcmdYIhVFhfPS888F0+nW4OiB+AbOuJJCQefDMx5hqY7UMET6SDvLGDj2G18TaIrsc
Ybg7Dn6SHnSRX4LsbFaHRtAvRW4yNQuYRea0lS9+9YSAeIqURChkJY6plTRRnQ1pkY5DTZHWXv89
VCGolFWCciT8MvKQNPBITybEMCppQzPiOrt/7kVsUsooamsLJ4i4faLDvdl23hfC3Q8QwgFsWact
5kKtSSxov+cwDjVXig2uyyUnlsnx6i7EQSTnaCdMlCs1liNmi8pX3SRih0ldlK2GEvahkH4AaYNJ
VZiWr5ZSsQ7jIk3UJc7y+MGL8rS/fhIj4webzc9cAADzt5hMKk+cjFAisrVZ5+6Y/ByQ4TIxT+aq
y4l/dv6V7WBQFRbo3gmlCxqBQhuhZxZxmAj20MjWA/HPN77bIHjo6vSUSkZ9Sw6i+FzofV+MPKJ0
ao8sAFluU0fXb0I3Fmg+1w7SWFJ+rolaZLkoZthk/KHVEx4l+gyXjF7+H9/fnu98Lu+4Fub6QBEw
mxkYpLjbeAeNnvhX9PAtHOdUf6c2vd+ygPX0UOnxgPqjOJq5gH3W0dlYXj7FM1NvMg0DiS/NyxiA
v98woLxAIiLGAOPueqFB8yV61BWJRyVeAxUNwU7dOVg7UiCFurDl0QPZxYkMj6NBqib88IMFxDU4
wmw7eFfAi/Fn0Vlukd8M35CuFrHvqI2NsSZb3XH6NBnoFbAlthdgqX10t3jCVLRJ+Ou5Fh4ImFuB
RYsdWrJB1TCz6XkDeeTLwulCp8XnXcQ9S07i7MWYWLnwLSvN9delfd082C4mJfEPThjwmyZwuyKF
WFH0Hrp/clIFx5c1JXwk3aCw+19FrMJWlpLvmePeN4yiD9st3yAwrPQVV8teNVzUx9n9RWVo3TxW
cF3OQqyjXp90TzdJsOt0sdfXaSf4SmZmrNuiciaSCsYmEm3Bj3r55YmzAtfYEsbtwoOW37TvVtzY
+A5bAukvJEhyC8g2PM7vP6KKW7uk/YIojIvr5f187nuxbx7ogxLPcaBd36zUebVxVTqcbb5pSC+A
KBHQD6oXJvKonSp9Ak5ZHzXZn7KOfqdHgnmdxIdkr0ZWZ9twE5KcBnKEuBEwzUdOjMxkS7laZSRQ
hPQZ55QRvbIgh062ZPyGJb+tueNDPTI1uIO2U1wNRg/JNiZiHbCtS8eoZC6OzvGHLvy2GSu7/WbI
4oloUSINVBCcTv2RUy1H0cwf94ggreYpSxUKSuRYlhCRpCJvv6suLxkGwepyujhdTy9XqGt4rbX4
Dd6+sxTBbohAEarfS76XmhOLnbb6+JoDd8FZ44Hmh3hw1CMrFkWhjxk27l1wqw/gxm5HqmtqSdMR
TnXe5fkG7w+ZX7BTgNkPexku0wT1ivyDsajDek6yQbwwy3HfKaJGcvVtsgCrat4ZMivjZ1AIA3eq
/xmKO7WVEsudaJ3lLjHJco2yTheZ8yx1AdrROT8zruum5Aj9OTuKNyj35kbfdD5kpUCiBgAOjqRd
C2yqiCg2OnNEYYYyR8Hd6htmv/c08W8eA0bNr0i3eVrvn5AL+MxbonXwyXdSVO2O8Woivyh+eQBE
5ZjIa1B5aOFw7LFdAYmop5U/AOlb365SN+W3MkOWR3MTmhuWFsQ89QXoO/b1TuOe1OON0by2gpoR
kgs5cXeisriMtYfSUCYgUMdbCtn5MFFmknR/9FwtbnHF+rEmTrYeliYwbPhLuSGEi7ySVqcdbWXR
XJoLau8sccRSMUwocM6cXegugU004Ao2kYETPnu55uLZKo8uhr53EGZIGc2lijO0K4R6/vBtTDgX
JPpi/Ek0HkTajR36cWI9XXEklFzG/IijeHhe6LYNLcE9owW53lfP7+MkNt8KazuBgjqt03F7N2zL
Ww8fWX6LKw4BcACl8WEoy97zNL8X7SLDNp7upa9MMg9IXCi8w9Btkf+a6TcRWS9ppaX4/rX2RWqK
XczLwKbHTV2iyGEl0+wfhtM2jrSirZ3c5U7NlAeESWm7r8kkB8v4jPgoooFErx+KITEQgvz5h4Jq
wMRoifvNY8iK7de4YQ1ePMBu04+1YbY3JeaCADtovYcli1YBYvc3Ci88DJFEynAh1NglvHRlvnLK
0Io/P/+r2T/Hmr5x+sCy33+WIVuszq8LOlOun97fw0USAB0nKAypZy7yvbbyrtZlamoCrae6TPPh
oF3O7asEcdlMfecTCeh0MM47bByLMmZXfW2igXZaCSjvRDSNZw+/dZljr1C2TEcZsU/dBpHS9jI1
RPYS5hMAsN1YYyYmHuK7WITlGgrVma9J4BEI6tG+zQFW+DLEkmSdyE29qCh69qFIQMA4w2tIgQA+
MM0E09OftXsIK2jmyoBbUMlYKvpyBK12p+BaMpo3COB0biYWUFZLWhlU05am1zfoVlKBeEK3+7l/
FD0/d+6fG+XezlTp08EJB31ofHFU0aFicazeo9X3JFffmlhHbJYx/Do/p8gDDWtc8zeX/aAI0u02
PJW24s3dudnhuBRFLeEqwwc6FFbBruNWp42a4n8ELRKpVGhjLpJHz4WbALADmEejOIo4EHog2oER
tlt6xYslBaypYc60qEOO5/xY74M8a+h0G85W22xeQ30TqYT0kF+mA1EjRF6dHb/gN/jGWLexIUv5
oE/2ta6JwQFTJ/Wq3ODBXEvHMfgR13yejuFqvZDpWzG30tCl1jdsLE2xl+WpHMwWw3cj5jNTBQRU
AT7+MdXu2kiZdQhuf2FEHQOaHwT6q/q/PRXYvicIDQPBwivCFtSRpQANxkgB//wWxR+nM5CDwm8g
uBfL238FqJnSh9b1Pm+OCsQUBtrGD31tm/B+ob6u1kxGSHrUM3B8pBn937BYQ6nZ+jCNxSlrwmJW
BKpK1PfQsCy2M9P8AyoBc/pU+AtsnwqmQUVJtrOoKeX9wxVUhauPztX3nocgpgjU0E3fVjVOJ91s
6heBDuwzN76SlcNlapDBnmNZO+qZi7gWJmGgqvqn4AVPZvB4utnBzSUDcvXg69wJ+o4h1WOhkKmH
tGNtFqxi+e9k/TWmuyOkTIXe+4FFr0WUCAPJzkyvcFLHWw73VX8gF8/o8fche1C+8SSRfsI6RHcu
xVeC3JU670RO+rtYJFfF5TV5n+AsnWjTFY7EFJHoAaJVxLHtBdxc6wlKe2bvyO5/xqKRvWQkJqRs
eTCw7Ah78LL2Q4IHch+F/M18Uc0ori8KGAq5QYQPbVm2yIoXaYFgIlljmj+DRXxJBoZw4902tYG4
f+Jm26KJhD74TEESWnK+wA0UlXQt2Ur8grkvZbOQUhsaCMLN9RNHEN0RDZ/H/A/vPG5LNBC91pad
bGAYAY1CK+C73vUY0j5AmpHGcQjmggyXVMLa/z4ec1MLnIfbmvve7gZhTGiY8GGWPd33Fr9F6lwX
PSylzNVTMB8Srkzp5flVd7rYwLjDRXoww0o/6ky/7eLEEHbMr4Hk3MYybUVos/Pz3XCb82gx4anH
Phy6R45YBtoJzAuyGeV9DmIjnh3/f2FBZkQhaR44ZSE0kgVAlzetUd9wSJgSPTkUF5UW/WqfoX/A
OQ/wCyfe8cNH/mFMDHS9dGYzWBCD2d9WKEQtlBDvfWfA/xHXpAaNADeG52Ha3ZmdY855gQu9XjxF
fOv4ETlNIQ+EMaCGJZ7NZIkxChgc2SR55JrYOjctPRyag6k6RY5cKsaeNWq3WcQu2nHLvyocOuQH
+o6LjAJ7wcyKw7OzlQ+XA59cyfgJ+V+0CUQ8JwchhJQThyD0Io58/VpdC0ez6KKBMkqub0KpNUys
7MdBLCZQJj4nD3rQxGhClKg/9LHHLjrGikhJlusOBkngRMgJsi0ivxcD4Q+XwoVDOfREczXov5UZ
OyUHA4YJu+APjnJjPQ11Dq7INX6WfRwMCAV7z2m9oCr7tkIdFi1XxirkDZUyUBtTdwu+yUSlX4rW
S2xCUcr74EO+eLvh470Jz2tlv8WC+mFrcsKm7pFTXRUKfoXFAZ7CYp4fcvXI49qEfynWEsS/6J1S
0PjVlSZDREuCi/KTmwtSzIMVRvYFKDvqsokEP8Qi5rG6gBCU0NMdx7bDFAyQlZ+RA4ddGdO0iJBC
rsxZ+oHOt0CM3d+iCaAEZ8HhWW/XkheXbG+8EzxlP6mguDOtfmUpBNEzyCulj4nCBqp9CzcjpYZa
2HpP1/NThTzxI2OPAkHsJoNWgdWArg7EPxHrv+fsPZXR3isnkZJya7hvQIgQhvEsokX8I7yU5Y/j
FmX5yKf8ujF/Q9l2IIK5f3JHG/r4Cn1yU05WJ8PYC7o/KhHnw0wL4NUPENerpm1dsrfv7cOnIUwo
h5Cg4T84mI2UzV5hCgw1mvI8y/Pl4cPgl7BFB7hN9o4Qw0PmPMm1XMmYG4qSJ5fZZwAOB+FXKwuQ
U9CVcot8G1u3H5e9CIJj/5POz8Q2Ojcue/QkHp8Cna/YCLINxRRViCDFsVjBNsF2q0g7PAA/U6Lm
CX7MDC01wfW/pC2Y92HQaYBeT0mj3aZ2HaIGYgrWfWTGQvTpHIggVIi2xB97vLEN7Yux83cDb7vq
JVoxc8D/nf8RfmxP0OgP31a0wWqUNLZ0Q3yEnyidnJAPElFtFQbCEXGI+LLQ3U/mwIl2EfIatPCL
3HfgpKDrmCxIkvT7yXH15Z1ppzBstl6oXjFZVOaJ3yoqphwMJG1loVMm6qflHw64kngCAvba1TCU
FhdqvkCfZ6/YZANmzrn4tPJoTKgq/beICejfdA3RJAtTpA9VTrJKUszXirEDhJ2hLpwkSK3r4EGN
TUFIc2DAHxJiyqcgGS8MHfMBhHOHPEl9l4+MSE5klISJrh7TtBUbgXVVG6eHVqxEcSCETsrAJ0ct
Q9yk0qYGmPZ8grhose2GZ0vLcCZmniLRbtz28ppf6laUXFzf8R7ygIO9taPzCIGIKgR+xAaOyVc1
+jxbSJT1XRNF8KAS/6YLM4Cp/I2U+opm3oBh73w8p9WwPna2w6cIUkRWMkF5/gIe4QXjJ+YQS+NQ
/+YOPfu7hFA1e5rXJroEL7nXBScmR/JgjV517fIfKAlINAKhx2AQPmK4b0ficqU2TqlDREoQ00yC
c7QHQBi1mTQk+m9Rhr+MjbiBGKq0v5raswX0MeP64Iq6vJNMxSjLuCwVzc19XgjB6dW0XC55RQwu
GrciIY4eG8+lwyMkJODwfGLy1I/D87JAedIlAVOqRY/nxgDSMiyULbS1d6FVdoJvd+zt5ffj1Muc
aX3/bd33p0QBhoBur6YydfbCB0CSVtc8y1Lsm68IIeKR93nzp95wW7ZrDj3WTNzCXAjFYpOmYIad
aug1xJTYRCIRqzZv3f1y6OvLb28OKiIFeXw3gVg2iZZagdMiWHPZSBEMkEG7uURoU9j6pqrQB0vF
rnb80+aTiyJDoQeazCTMDH0GixfNXSyv13lHSKx3NPunckSpfO1I4Fe+2kS5OzWzsv5oeD3+vWMR
GNBYtitMmnx6a+KWUOq6JmPKnpCoh0m7zF/PQOQ6UwUFQFG4xUeJBPaaUOnQfSlcb30anp4vS5oK
qIln4v3MgY7BOpvIu+/mVhgF9Tl2zs6/rwL0yaM7XPLLcciKNFW7u9LtmckIM/mKgpkYUTuLJLft
nBzuBqQ+vczEdGdExmvdPA51qqnZwl22jKoH86wcJ2g+0V6qlqWYkzstvN3LhOuryoDIBWSfmZJw
bvf8FOWUh2Nq9pI4sZOFexcrZfno2gEInbV4e26qh5PONsgA/L5g0KhosUe0x9C3SYvdGy1Qf5S4
txcbrmRJ12+zsSjuzPxfJ1L5p5bgK7SbRTJkTWukwK6+POBApXTtG3KHHTOGZfVBfsR+9GH6r467
FafhuNLxp86AoTGnwEqu9hBsWF3hKVOBDrCynS0H+vBm7fWbTYC+4QlPR7UKfMtvlpw3tPZaLLHA
822/ArwMXfk5GWZ+fiyYkG5iWRUsrk1y24yTwRV2OIqpZtpigq7JGTQVnmDVptalglASxHzBVZlC
UItBxl6woXMRv2PI0yj5+PCOllLxHwBCHV6/+UejnjAIvJcjjANqXrw0AG0r7KnyDJfSFgEvfK6T
xhydKLUuD83rSy757yOhfo6/wGWcFP9V17xTMveEG0K7ui/Zp63nYzujslGf5UbFvQVfa0BGoWzB
ytnZHQDLXHOaIAO3X9RyfOIv5D4dPfVMqu45TREkbqnUm3XV2+hEY2tC+wLe6f0lL/5CHSJkaGxz
lq0z+X6PSi0lwFgTj5CFB+sOygWSa3q6HZRR9XaWYQW/iTyFq1JiM+gFVyr3YOXLBOJRoW46knot
NsUAtX/jyVCWLvgKuwJBb2nO2UiL3/BREF93bqIZ2CZ2uGt1FhZrs9jGGmSWSrJSjRpNCyQtCVSV
WOYDWCoSFH2565t4PJrQALu3f04gpwTQblTlRz7xHpFPGz0vFTINJB+wqEw3HJGH56oz3TxxfvuC
knuqZ2jvuH+T9mcSmKHsaN9XOa/CI3FZQGtrtIf9qCjcBh37h/qgnqbz0oCtMAvaecNcDT748LPo
NI8nDlnsdxfsFdmmvG0/4yRKfgHNaXTVQ5xwvN5zKSnGxeyDtQJn5Edlhe7eXsehyFaqrN4PtrMY
vxpVsemLyGBGjvn2Xv89TuWwYnLnNgCsBu+pOXw4ULrBVXzBjmoTZS9YtjFRHrrUpcvluZuavWOt
/v1CQiW8GuLIDm6WVxJluLIecmlorZyTxIpiOdGFDp+sYb3O4MLPiXIp2tpn5oki4xr/eN4vBz4M
HvLx6oDjqkQQA7HrcBMZSKpM80idcPbQxDg1cQ2oEzWI4aKqOWs7GVErdzgvwJWeS+E/Rz0F5ItI
1emI2YJvWaMG4YzIbJCPzASRPul0TaGnEVzbucXmoXArhEb2R1xS0nUe7qEPgfGXJb+1xAp7cE+g
elR6DnSySHrvn6UKt9hpsxw89wX1nwXkDzMrRf/L6nCWiRtZVIVRE7N1mvDqC7wVlHif9UNkJqEV
t2a72OIMfJTPB+aV7/zFhvznhHLF1fWIc1fmDEHvOjhWc7dBW311v9oPqpaCGsgc/zsHu+3GJhl9
a4O4V+b+PfqJ24hNo/19Lm+4PDjY6fTOkdzOQLYLKNarDXrI345/E1u9lTvzDRJdDgoMFfJrJcBB
i4jSuREy2HkCARVVJW1EXymQCIsiIua82y7qNrZ4Xa+zubP4+walQUcRv20b/lKV/VZl9z7L9/2i
sxlspaY7QqABJbMSKIzMtd4ii/1ROYEHatwvuhgboGmc1SY5LaS7gWE4O6EvnIDgJpqyAp9NmFvn
y130IzAvUdHIpJT3yNDIWflJpGvcV6lNYe12WDARiL2XRKhAOe1zYGOQrr4OPMEiQxUPPT7/dWqI
dU31miM5dd/ehcj2MNPKVxKJPzlNvQlrV1UowWS3vGOiRTh3Q/2+PmzU01KKI1Zy+AbrMVzxR6Pe
qvDgA4DnsKLF2x0DtgCB7VDWfzLyhFOUaPKZ6vGWxFknsRlKLsi0sHy3p9nQ84lMmZ7orB93Neot
U4DjO86EPbeUm6xlsjf5X+ALL2yJQ+cIqeQkbWy/JAT3KR6d26x8mbNzqvSm0eCQh02ahMXJnMpr
mVAZmnvB7PQar2vPPptN7F5KTB24EbDHwf5GWH+3myn672RfuYB9U7i5TgNceZN9qCZhPhMgOGIO
rmhKCE0ZXdJmwntLqBrFm05lXgWUZh3heuzs/k9NrcHw6EcsgMth3yQ9QYRL0Yh23aeDOwLZf1eE
Ic3hWWkThJergnlIwgtI4j2rcLPWE+IQgE6l3jlIJULl4YJV2DNQYthyWQ6Xf5rMCjzTKvxoKbfR
dtPu7B2N3dkBWU1burnPl7sxTZ2cCi2hhvGI+VH4zaCyhlwMSg6u1IuB565xN3oD2gdYt2lv+S+R
r89qc/EiJLhmP6dvdca0xXj0ELqyGJ9Ti3DvGR/8rRvHag8dtRgIbJy6F/811MoO08bBz0Pu9Ara
rSPRJ1PIVWfDfKLBKAhRhcVwyonNNbI71/nuawpe6eC07gePWZNv3s8RsyO8B5SjVtA9mEBGGrZA
i0fJk7T9n8vSQ57qVIkRy/h4r6cjDyKrUXC9VGvegpwuNqtBTU11GrmpIrfD1wCBQAT7EDu5dmcM
tdgDTjl9ZtAJj6lIwMoHjFNjou43Naap7RHU2tIYvXGqNG+tbuo3xnFu9WEd42coT8ZZtR6EqIAi
D1P3ou9bfYJdDpFFu0CyfRF9H9pSYLtezllSpl1/4ryipHzDgNYThFQJ1cyGIHfVyzmlBS4yFStj
hQjrNWHzcHBVZoUXXnlA1Jyqcd6VdQyhR5eqVhsAf3aC4cugIYrwS8rJFzzBmNGdmxwxCPLmGNRG
3ZTcqfbzorr4fjJrhPE/YyVuLUqNkPEOwRnLLsvkesrHYsmVsm+m3HCoXnNcsqHsvZc3xYA4/GDD
vf5UxGLpigWRXUjKV+H4q5mjtuLMU/2JsXZ8OvzmgEtqJ4D8BQiIGHHg9WJYCdRiIDCtYYcK4kKe
JCoN1JpKONuECF7OF/InXtLJ58q3qGowjfcDRloZ5iPWj8IlwLspUrYIOWYdluI2QWG9mE+cW3Fd
u+sc0vhwAry61Rn/yvIghiFeLgaRzENKR8ozJlKL00mnVf0oOBZTO/cCCTX4A+TDBmmcIXkyngjt
oHyChLtgyecDjaoqj2N8y2AAmGoxVV9FMFOBkLVgcyz6fMpCr1kuMwWrmYYhwl/UlKSgGbzySiAC
3Row5fdOouLEX4AplpZIL+KGnnMuUKaU8MA/BoBVbSJl/bAhw5mmBXEuLoO2t9cwouCIjzRF9icG
lzMg574yR059+rVHPuXrbJZgOMNro37w88tENMKnQM0jz03olI0zzoJvC6KsuC/z0NEPjGpvDaKS
fsWmtCRB9Fx2fUpaEtfknY1yhi0wcWTL2XEk6xoOGVNI17aH+Mg3cdA4ZeQBF7IA/MBNYMsQG5BO
Fid6O29/BstZeypV8FH8APffsdfQWQVXwnrRb46P8nc//41XTXF764R2faqqfdzEOBFiun9sG2eo
k5ZAt/HEjYOlXpc2uFmHKNFfi8lRLCHGAp+i7rBW9Jue1YhnsNHm1ysx4qmURauWAFC2VMntnQXO
ZlaypClLAgF8sWXmp17cDB2SyuKzA0dqlNqfmUqsZGW/Lup5BC5bbwNPfpkkocn1u0KNoBNqAbXa
YdX9ek1ArlHzJda9mGBvYsqOL6kwJZw8G4Du668DUqVEB3AKjZXT4ardPSrx/8EyUkUH42q2GjIm
l2oMI6iOM/L1yiuta01kPaGT56T3XMgTR5ODVN0tTe7hkzNFu4psi/fVBX3fU2H3fRQ+4HT8rRtx
Jtk52/2Lcv+iE6Of++7MAgz8kXIWdC6n63k/QbmqUBoGKMimVvm8tABEWv55+vsphbkpltc+PkUR
MBwaNID8dKTrnMVoEcVE3MOnEo0I/BbagVIh2vnQO6EVEi3XII68Fokn2hPsXL3U+TAqNWW+dFQG
XLWzn45+howYLWAzT2xrUMKiRyRgUsH14Mnw7aacIUeR9BBIxpyyPKjh0vtd0gDnnqLgzpSUfgk6
cnm3uq1nXXyyhhpaW+j4UU/Ch7g80EiqtA+qJHnP5vCcQkIV90PU9lFq9M+kmPLBeEQHGzqTWiTj
ycF4S3tDQ37tgX1cq8c3dk1to01zyxRmOMDRByu0mOu29S1bGZGi9SCTwKKXPVRRSMd+z45QerGf
CWJWCZj4h7nQeWn+BT0DxkpJl7zOHXslO1z0KryYgF0DzQjNHsH6NPLFHXLhP5ibPjYPhGPqJToo
d2jCk8/SyGALaWnAoWXO1ovqHBIZ8qiDBlzJTC/RlrdJk96ObbHGCS1cH+O06/Ah4jtca9FSg1fq
yNsydFCS0wGhcWbRPqmIfwkdqs8p0UbK0GJWpBEUOZii52PjUY2+cHVqHuJiwBg6XP+GRhqvbNvd
/LouhcamlAVrF7rAUrz44aOUJLvkUcqdkrdeVtyJ+Id8sJWVd/nO5BWdjAEAUe7ShOf9gcqvPS5a
bKVHCTZkphZ2n1EPX0R73Gnsh7jvINczDUWUnmyo8D3ZLHWVtmmQGoM7dSH2feWih+IqGPQJ+swI
Phj2eDP1W1Kql0xd5hcJq1rKyEFWCqhgnrcOZztCpoiszEokAvPAUsooie7Ac35k43wQ9hSvIseW
3zK9k0+OJwX+gGY2zIJTJpLAZpY88zr7EULC1WpO12YiAKptz974hoA/YnimEr2X6GFZrHGlpD+u
BdMM7jUUHlt5kCuj2vN+JXbLc3EokwVt2MgZBaix4NARYwQ7jxbi6Tu2TGPfSX09lssqXklm/x5p
TscpXjMqPD5C4hjo+B2ZqiwiLTCoUwNGEDzcz0Y99G4K6ENPO+2WCz2FYlP7phZBYnGLRKj8yV/Y
WS2+MsAqUU1rnRRB/EJvgaIVdn5OoeMfpOCw4IzXfuAUYL51pQS7jhpSsawADfr0TKL51vpB/YAU
X19GKUfqzqNtIqZ8R0J1jQ2mEw9A4G/rEahLOzNOEZJX4TeEHtnjDrsXZd5JLmcX12Oo/hsekEJ3
R1kYFJygIObETVWIPw2EtWhtFpLQCpuB7VIvWRJnfCWVK5WN7/yi09OkBExkEH2YRC1fdaToUnx8
R+xkf32zgVlSyHsDHdnybsXnOSEN7AqpJiUPlaW+ncBZ6GeR1b0UBCEokvH/vD9sQfFC5aehus0d
XrT/Zd/iMQSHWAfro4E3G3cIBCCRHF90VrXU7XHYepgN7vDJAqNoCVh9tceiyQYZMbCfLZAAynuN
SmPfqkX+YWdOyQzhC6uKuTMlDb1Ov75iCWVmDEG4b1kikaiYk89aiBXu2zhznWJMPng63mjsIy6P
XqXiyzFugByuRbNBczcY7F2gyrFSO7X/NgXQIbUA/vZSRqrXf9I3ok6xSZu1NijmCXjOBMQrLMza
QJmxwogBQidWlcJpizgqKsuziQm/hb1MTWtYRJZgZMKGejuMfJpOwr9GVO6kMcGs+rL9EFFWPvs9
5cTd3Kqtn2ammv9w5zJhHT8gyN0qJACF8iW9aeNpkH8TdvDnxRa1bgI3r4vNTOdSrlVDxX3SyZSP
CMz8UpSEcR7/6ulnojRAdfz5cPAn5TtXFFbIdwhegy6itdvf1PxZd1wKkNsx52ldmeor1n5SalbO
eT++LV8eaNGgMYWRiNpWYESuZpzDXQNk65b4KeCDOoqM+BoUHLv+jP3t/cTrYo5InvuvpUM5eGhL
MlH1AdG8fcT6kd9cuJSnT2gUwLMxgYpS7sjg2i/Bkn/FIliR24pcPP4rCM9cNVR27oBMGrs10qNW
LA3OopqcJEFmGzvkLAiLIxI2Ng4Qwi+ib4RE0wOjHN816ZaEcBkn0/ODLBAP+OhJ2ywbVvIBM95e
ioL7o8xIBDp6lIpJn62/WPPFs08ZYb/2jHqVqFS6zs99iVaF+ksvlpLSDXDa1kwE3HoqLJwfFTCB
q9X/M+1dmu0HRbmDvTpIaUyPsoj8jAaad+NwxmNqJt1ESopexLMVTT32gHyUxDeSlg8HZ5qx1zPs
o+t8khcZU6V8c5cxFk3WZn/V2ZZCNzw7TmX8iss3utFeeGm7rppVgOCDJ99/o1/+97C5xQNrwRww
U29pwT0gJUY/bBiwLyH2nvGkVoUA2zYzCk7fXKh3mEaSs/aJIVimqhXONxY2m/1L9aCjVCa4vRKp
/nGi4NoZzdyXlbqIiMi2HTEg1pyoBrf0jFaL1Bdp7PhVWtMH9Lahs7LhP2TPmkqH0xWfy7grAGC6
EtrlVpd4BjcIcAxhzBC8N9rstLuV9tUKffu6DRTJaN5/1tns8zkgEWTe3s/+NzSsPVTP/jih9/pd
TRHrZZ6jrlpyOflKbv+OwJ3AFOK3R63tLd0nOXcSSxYrf6d94Orb4UxcpaCLbZhL6R0IFT4rq0YS
0d/qxGwTiMrbaIhhASrw1tawZvTPWOxUf55ayZxokQvRV5Io2ITqbSGpS8fsx3vWnX8duygTEBst
E0SQqSh1ilEpY7n53tqdVISOZ8fl86gYJXJsrLwSHZiAkBcukl1EZvy16liYJeZJkPJsEroXD2FW
keJI4J/pvZj0FPHKKYK70xvLgSaVo7NeQ2wtGRWH5nvN6hzvzl2h0jO1fINb7tU5lhceWcde0vJV
BHAvfWxFX76ELOs05kYOKW0yql0/tS7v4xtj3NBG5TJX9YmVfmKqyLahzC8z9D7gGY5laPcSixM9
tQ8V8o71FitKeETrhhkLf3ubjna+4707CxWyrpySkH4gd1Hthb4gNMAju4ace0arxCDEwbZ86mIS
3RjGO16QLUnEnWLgB/+7iuWeP8E/u137jm5LXlR11JFa9mKf8qtjZz6WnafJGjN6BGdSbUTqhruz
2rGzGjUt8R5AkFN8d90LO/fGmXR4Hq5A+s9g+2Ac3nyy582NuwQkkDB5J7zP6pUbTGnm6xtd2ZEG
AYyyyTwQVaaGI86iCggTx5vD+ghM6+7+DEi4RN0f2kFmmHt2o076gIChbMBDwVr1Vg5kmMDFQfhA
64JNB2gRRC+1Div4kxIZS4rKIcZIAaChuOxWS+4tnCVyLeQwgKytDEDTyOmYbG65q6bVA+edLdN3
mGwycP+MKKBe4xwmERuIpnRi4uwJdolDFvqNrih2ac/rSXkzAe9yH/CgDZfttpM6MMZjq9ixoYVR
r++YyLsP4fJbEv0Zu3PKRb4wjYJnLdg58nlBkvXXf4KNJVcvKpj2TAaHcPhrhL8b3hEgkq3gTGND
+0cYfgeW8s8ZD9VcKHq3gqt0grTttnSDydhtHBGANZy87XM2t/kgXYI3DZdQdhyL9zkPHzGOMsP+
DZo/A6ms+abtx9cipdWEE90FcXqWkyGrmMy9krHsCcxxvOOde/ixjSZsjYYa2cGRcQCvcnfcjjYN
KmmKItGtOAwadmXF5KyYAqDwTTmvgcUt8xA2Vy0UNwqxSN2PlWzQdKQdy5P0Ny38M96K7btnmJ7u
oi3puLDkyj0tXIYFb+V1ioCIlBCxSoAWTANNvsQYe3w5ibzdIQCdJCjBkXIQc3v1enmJS4GbxW+5
N9JnrKOYewvP6e/J2cThDWRXWoCUxDjO5esGPaxB6HwdAZ1Src/IpmDPOSQiJsFZ/CHjG9F4Gocv
UEn5E4gtx3RKAMXfDFZeJ8i9TLqrFa+askORQg9bKAubMmLWSfBfUzhwFLOWPkckfEd1sbt8PHSl
Cv9i6Xs3vykhNc5ynLeL0wgPdn2DRz6mzUU7qkMw5j4AA1nHtg0I/8dAl2Qt0SUBcsw+/RZcNsot
mzxyXEQWLoUxZDByeRXFX/6zWLOhNVY30iwwtumjl5Pe+jkaJg4ObJOEsrgpIuXKVuywQ+CmmudC
dCjhWbPvvR9HYr3njLYdYnYpKYAsYqZ+tG9H1BeUfEhswkcH0WHtSodO7W7rNWQuETT0Bsc63mOv
QaFCf7ZHinf5x5YU4uWpxs3PX802rbH/SocAee95KSGaC9XvzmaAGgo6HJTyN3tztZWskq1bNild
wFAiZTyxnkAPbrCme7KD/K/Nz2A5P8IEsTQQkn00AkOvgRb25H6jxEe2ex/xjI4qxhzeKwt8wlCR
3rRdPxPW/0d5VD8+QO6LXV1hjuh6nXuPoorrl+3e7r9TIAbC0IBd8ppRdPHpwMI2oJcIqnGQYSmC
ksWOMwZU0KJh/D0qVcaElFbn7mFuEBChM0gSnlRNdEWrmrPIQazJY7dA+enFvVSmPTl7Ky32DyFD
4iMFc3/Tf99W2eokrR91S8FORm6ZSu0LROxmAsdGRq738AQl8sRfuSm0Q2jE2m7dogN9iwlQPWZp
7txJZ9kMaH0KFBvz8Cke5N7LuCgRKClTKMUarfuaDNThi3ieMi/zhDBTvQA8mx1U8qzRzc1P48Zs
3dbQlho5UuIX5jF3+uLDrFA/N7FH69Q9MIWh0oCR+ExWfRu8mmX9NTuPtXpz4MypN3Gn/nV5o2vR
8fI8ZH1+ewbtTbhefHxMGMcg3tN7A9KmKUk/sBGpo0khXGkzxvzwfd0/nkrGJiRFtyzaryHRtEIo
U/2nVVq7ykN8JVKp7kC+m+lfyxXUYED2m8kWonlc/GFUOCex1SDXhRgQ+EUis0W8ErvQvczz35Gq
4GMOUGsCoIov5uA1wCJlsWE1v4cIBQ6fzx1WSYE4l3wQeEGB81kBlBMmZhIgFsQNqZEr9ssfS5Fh
BjvtMzsTPs/FZOjt5h+m0y0BB7JPrQTEt/2Sgw8e2qglEZxcOHe1z5B3VmExNoV8dTlTh3h1MRcv
9Kv+RJ1UqD8z2+DfAZVhYCY+0EX6s4Tjqn46x0veuq1LuEZ7pcBwkDeLicdurhleVdhJ1V8ozyD2
IlEkr7A2+f8cdMwRGXHOmig2Rmp+nVBIWUD2zbTNXEGxmEerFxV5Dstf1iNEafGlmTo3BSByQtTR
pXiWvtHE2AiKdNQ4q5DuzWH9bR6JH0JhOjM2fmx8/Bo2u292i3M/jzyyV9TDMKCf9wNrQXwp1UnK
reXcSv2LQBtM+YjT3w94H2W0ojIeWlJvznUR5gZlsu40x7I+jUbqFkum1WnIcDS+C72U5DgG6bFG
U4Kr/1HttX0titbDaCTBeAJ9CttIP63WHc4BBHCuiImXQgwpytXSsBrLrkyLqT8dI8xTLS98+aV5
0UJiEZervL+UE4uyoez73PAGzP4e5E5VXnpLXBPXC2vbRuMPg5qs8Ko8ZOCAwoRwCdXP6HKl+39K
kIJmoRvXIoz04DZJoXIHRzyP+iYU17DZ5go5mYgK9qxe93P/6/x7Lt82+oHSNw8eWgL6MePL918I
hsWPzjz8GRh0kYZecbLb54GWeK8Q6sTOXRpmCjsFFhLTFMAOkopSlLE5JR2340GEbYoC7Y5t25rh
lGxf3/kMigU2H1iumfcM/54c1lxLNSzHPRV4pIbacW79UkouxF7qMwyuWfjJlV8QX2B70O/bpxD/
MMYuksFg3h2vTabZEwNrnQkr2KfAjKTl49QnwFLB220CcQnaPKt/JEbIVFu2Ok4EnvjzuqDteBfB
JqmlZws0XUc1X3X/HGRfxEkrFeD8Tt35ifp0e38bPFwtuUgCg9gCAm8/OBdUkIvQqgmjjMEY+LVV
HVGJP/4GJNg1KnJ8XxAlJZrvQ05JowxE1DuVSRH94J19l7BgMeFcUhTe/Bgxtxe8h9cVqGPayKQ4
tpS+LLqZp4yQaOcemkXoWIi4LRbsrY1e6TtCjVEkR770jg5ojb3pqqYYRIiyQbLEHAWVglvpIU0C
ovpvdH21lUDU5Cc3iKmrYye12OkJbv5V82YQ6puNmJBVIg/uOVRPKXF6blYVmSUXZDeM9j7O8MPu
xbVpwHSClHUyj2uzd3RmfRUB9dyLMb9G++ZZX2y2aAWBW9PZGZLDN54i25xEa/td+NB0xIeqRWCP
s/YvgEcTFbkilW2JWrJ/YBFxGg1yEjb9rIFQxDcYcGe56I4QPMKs9aRR4sY2EE+LdSuLQqlNG9zl
kEZTxyobS8Vyac7vkh6xZeoLSISTi2dTlg1tRPXjrEjcfbu+d3xO6JPjLDOH8ETXANPlqSnAXV8W
bWLHxwwnUmbF6mmCIp6gOFuUIrghvn/yRZKR09UL/klNhxLeMjwdoqwjClq5F0xD2MqTmdloCCbt
ZleVTQFdQFHlN6k8B64qsJI9Lr3bukOdump29PTE76Fu4wMSA0fb3JnnzW8zJWgCeiMFX+17/YXF
pzscoaQUnZTq2o35GbjBxK9sNQui+BynPop9xG/9i+Mo8ZiNboer6Wb+CLHhFLJ+wMIZlqfdhOnN
kjPBXFeN9ps9fMaym1M/QnrEVfXTm2Rq960cs5tgK+c+sT68kg7uEmo1BOWnyp9SX/sr14vozZEo
Zp2uIruoDzyZGq6w85Iyqx5OBs2jH3YSXoKokDI5rhITZ7LBpD8Lz5TZC+OPua8Ur0s8zeF4srim
QwzFLvLTtc1dRj7n3BIdNdcd8ZE6QCPJ0bH1dIuWDT46/RZjJ0Aqy0Pm+tiFTG8pSIwQ9f3+jk8r
nzoBGVZVmsNJ4mbM4Gs5RFT69YJz7xHea9oC8G9mKAAdV0+1nXme710HsEJmAvp2JUIk/wcYPq0D
XZRH4FS3TLkOKawUXp1zmfF8+bqhb/gChcgrU34sdaoQDrbUaaREfRfQo6HgicXbqNHEdj1truSK
yhB88OjQfH6L5c1iBzckluFGBfRFmsZIdXF+PJN3u9dkk/xsJ3XSMxrzutObax7lBigUiQDco0s4
lGjilyadIe5P5B7PsKWNYN3tJqBrydj3XVti1kgWY9gCXjSiNNpnCkySxOtUdJRE07B5Cm6f9yc9
e48ePqSPJUp2zRcZpDIJheNzV+BrpKWAYy1ZpZ2NNX2bBtrTiIg//5ZhdmReAg1MrNGr5Zu69ZJx
RF5dGaD8w3XkUnWVok1hHnT9hrYh/vP60/HlHP7Csxq1AM9tewq3pyaSEk6UM9TbDy2FJCvoxNm+
bt2qQruAu9KzSoUFncx/ceFJas6yTo3jIy4lz8fkoOj96tZMbVZhPdbUjr21YPdL6Bt7J8Ox4Acn
wIG6XSbPTAvoKnpABCXH5DbkgXNKw2dxY/n/MYtLwTzOy2FA+NwxfYqDcb+ez+aSJCsRP8U/a6KO
+65dqaEuPpWtKnn2npaoRFWmBRxcTSeYvP5yeZONg8MIqux8wRBNRYDWdjK9ornHBRyQAdimcisx
WitFxBNGe7P8T3JzRjxQYJAcTUKziORsvou2MVdCDEeAj3BZ/zSzDezNJq0Aowk7XtTbl53gzOp6
jFPP/y82nf0OS3ssgPSaNi3CsAX6qTmxlChANuUXystqBHoYjYiw5zv6Og03MzvPfO1/WQQR7XO9
bSMkDh7NBa8Xiy+WnWXOkJS7AvOAYhbycPBitVE1sTfOoFX3ZUkgXZAr1XmMu59n2mDoXJ0xKHgQ
X6FuuKoUcN/soILhmlmrY5gLa4X9tphNhJmrwVvg2tNLJ9XzIYqEqU7of1WMyz7COh1E5iAPo0BU
lXkBUXTnvaf1UAkqmDNVZENpwPUPw/UAQhI5GzCGv0tyP8fl1PA80+i+NEiWchFauOTnhjlRkI07
0H6EiFne9gOYJ1TcQLpurCJjUcNP/Z9EZD5131PKanOOQ8k0u/9QP14kV7WVTqz/Lf0/CxIKTpKh
4BHM1qRA7eeAk2v9rAP1+jbOrTw2fVkWRX8BJhOAgHWBpn/0GkEoVYDjUeTz5vkEx3mFORajjN9W
bDjd8/Y+kexRfHwdw79AAhyTIOgPuPPfY2hSVrYRFQmvz1V5lvo4Ju/gVPlhL2wqYfww2mgluya3
oCEq6pCe6IB0iT76TaiZ0stgj8tj4PHyDH2aWjQicOBIYLUwW4Jtq57KpwBjkRCqvURbPgFB37VQ
Jlq6oo6g3DJBLhYFrVazPiLriAvcl4HU+JNjihw8tMRQGhOiz9/PSTAd0Xy0CbTh/TEkvGaZa2Eg
PndiTXfp/seWYf32TYCRE4d2LUHXSLthQMNiKhpZHIpgLqoYA7zpVfdeGUDj3wUTSP7rylTH5sor
2I6/IFw+ymT6wsOcToL8PJHjHuxmpjuboRU2iVi/0PfvZCKWts07HW4DpoA5U8g5u6hgXD96qtCs
L1MLUGfnq0lf6eaSY35jFZiH5cgt89ChFWTpxoCB0rgEdbkqyZIeeG/OlZQcnr5d6Q93VJol/cpg
TI1T3LvrwBwjckIS71sYvpf17tGq4cud7WWDqX3MqrOW57mdqOFVSwidkZ4KofE57c7aMDi4vhTK
5GePiHEAeiWFFGRRfVlvoNyrdHXHCge2pxtoXAVsartjJyoJpfLn5uY/gqbny/vuW36ZbDNIxu2v
Cax88pEAkMix4BO3VGgLn//dAuH7mYy4OfKg/aa19k0S/a1g2SvhiX/HujGae6vf5rnawygNbakD
V6Uqwf87C+2VddwF5da1P2Ki5KoFhfME+CoP65MyU43THifCGZZ43/tNC8CuI0vyA2UfX5i7U4K+
2429cJ/7hd8W+k4ep2/8Rg9ohz0wdE5qx4oemxhdjCps8Ud8g+H97QmnRxHk24sbicD44D45FCRG
AJIqnrMvYK1JcLcLDuNYGbrFatppPb0k+GmGC0Q/1518faPU2oHebxciM1k5uvzPSa3tKTtEmUfN
BrSn3DJGvvLWm9F6FsO8ZgE5ZcushPc/DQeuYUy8OXoNQw8ShT/3sdUfKNR9jn8904LAM4F9PZ1s
4jzfOk6LX9NRDLTilQLjhA6fKW2HdOPBxH2OjXu5ChzSSnX9wRbl/bzE/kMpOFXbNX9Yfrvz3C+/
LEhqBu9HJ4IZ9oLW0UtljoXqLGVeTdXOHyAExo290bzsGOT9yo4WPluyQJPid54tQDjQJRt+/ySe
+R32M864a9D+X11IPTclo8be7omWkRc0qpkI2rDJRGGTZOamsNJTbfMcDPwVxWvWzK0gnkY21FJ0
JujULvO8fJvyetmzQ/3rC8w8HB2lQFmr0F0dGo9ONjUXWSmpTSO5S/AcU8Cz+pJ81SJ78yBZpIGe
EZlGi6r3GlRfwQqpavGKLi4S5/grTX7cEL/RtS3pTHfI8J/uXM/rdfo59rpTwRZjuFcB4hUgwGpT
fEBBZfg0WCZ4EP4GGhwoX1SdNyu6ZUdUFBEu25dbTMZmywsasIBjGSo/6ia77tI2fpNamjPw1btD
qdwHV7BGyhHi+SfvEwBRAt4yBqgJ/vQ3eMN0HnEoG//c8HB0gVu1hQTLhnRuXkh3jj00/J8I2eTL
gNBXQL2Wfh2n7IP9VqZULa1WiXzgSXOswyWJ+EULTuZ7FE5OalQ7sZMqd5MSeotYOot55m9lbXp7
yUOSMv/5/wb9mGh60NFx4f0pic6L4q+MSyGu/40OwxvBdLCAOzkaxxZ7xWOr/0+1gTNLIXDhk68v
aTnmOlWy8t6ZNTswqZWPEwF9pgBVtxElh/u/1ZhlLE8ZGtuikBeZuOiEE3eJglu5dDKFs8Uq/BUY
NhptAzYPmTWQ8y5hdHLCKdkL8T6muoelEWhdUG9Ib0IS94e333J0g07vP1NZXapdupzApbrInMRt
Wgh0v6gUYSheO0/LnMpI5ZKQiH0bWEkSigBLaHtNWj9Lc2a8XNwLnNLvqO1sOouCv7x8BzupZJ42
dWUMprh8i1fujgdKmPJoJsRO3VGMdV+C6E4M6/a9Vw8Qsor8M6QQxvEn4yx8aZ0zTk48nMNT0XIT
AB0y9QX/DKXBlQTZI/K4/IDWy6hwoROpZNe/RHf0wjKbKpppsAaulJCWi11h/g/67Vb/d9gKTRsE
JGuGyqRVHFqOpS1bTqu2p0PoJ1cr/48WlBBGFj1JdVhdkZel0e5nsImVipgpbY4yDL5hUHoHBq/W
EhwfyEgX5Uqz87cUd2kfNIP2XGl3lw6S6u7xQQprD+SS4NkspQxUOjcd7DdorsrPKfp0OU8K45G4
FAKizl798qIP/NaLARdk78u0zWPXsiwTq6zOcTGVsg9aS87ghGUYbZHwuzV8/voczHJgXOZ2dDch
02PzuzGPeRovMGfXX4FZJXRg5zEMqhUgMz8KA/PfoJPOB+FzA+H+99Pp2ekf0AcY2QdEd1KN9kFT
zvTX0MxFdVbxb8JUatCAL93YKESQYxaTEj2h0PVLB2KajtCK4ehs1615Nhb42t/rUh1J+xZqPQWZ
lWxfi0ZW7B5Tny5LpCY+YRP2AZJqrG3BJ0Yhp3E8AAAHFEzMu69cBVZ0p0eh7InSYJCNfLhJGhIe
kTnwxL2H5oCt4H+7XxhWqGDJR3KIAJ+cPQHcZ5IjvSeQSuoO1o14J6Vk05S+AhnTefDshgGCKSiW
983sRKrnIeUoKTyIfBeox6tHBx71OXvRKn+1hIjyA7lMa7X+97NKaLqxAzAnAbXSVWGpN7g1a+O/
owA7pr2rFwL8ICL+bDlTiyLuWBgnE/VFGgnOY7XtPoxITwF+qJAGVI/7l2kt4eBhie9VNVQM6+ps
KqKxV9DoGa4NTr3rlT47i1vRbEnaYV2T1HXiFgJ7SIvYg01KkjCiiVYsRGqVlKMeodRfnFSAsO64
FnHDtESwwt6sLZfUXWxo/NTM9T190TajePohHnCasiyzVHdZPoqgMtRs3q3SbMTNLMpz+3iBlGMI
tpPTIFPzA5/5R3xNCaxtGY1aC4axvp/AKXiGr4GzYgtsJ1ya18r8UPB6iFXTbTL/Pbes/S5siFcu
aGFps2yqeJN+nlKD7jkklgUDlfvVwt8C+CTJeE4FOomHVhEsNaroTnX2Q4Mqn9XnKnPJBNO0EIOW
HNGOh8ww/uK0fXHAIk34U4uaMcYwfnk03sa54AwfCF/24mSZQ6SsrVkH79xu9t7+l33e2aFaxKry
XyQUDGeUkyR+rjqbJW8BnPWjZvSFyQgvZyhVLh4VjIcnTi62k0kJmf5Wq3hZmE5qSyy4pamr/eA9
BFcxYhv51plWvY0L1be40VYqZWMs9Rs2c/d6JyDGSTM0+1Vab5BAf6JomCXkCEd35Qfixx10Mc+N
ICA+SL2VQ4KTnJzlbRC9b9wwKpkb+dgcYG7Lg5+4Od1ioCvsRHdPzg8m8Vtyo+vINKEPLQ9rrl8G
ITcIOlkwfcy3U1N5BXuPESDW1VpxxzQqWUEiMfYpFOCtd35X2crdtpZtWO3ECEu9VbsDnQiyo9lh
MCw41fXbDXwWr0pYsgbJ5FYM42xaVMzW/48lK63T6y7vMF74HVjqLr7OuZ6Y/jC4edH8qHLhzrsy
3q9R4QnLfy2xIsImbRtk8yj9o3UnutiamEFLoiqASmBiPjvTYQ5bpum2yFaiH/KdD6A4rtLrYSfk
PTJhWQ0nkImK/MZeOZBY572UlX+us2aD6GsyPiAkvo9TXcieKWDghxELITCo44SQR2m5NRY56Exu
T6PYZYc9tYmyNEzi6TsD0SSv1vpIId6O/Lt9p+M1QQMRAVfOf+9UC15DuA2FRuwtzUQi9e0IfGgm
H3p0uUBTo2OC9TJ5KN2R25BhMfC9ZcLBnEIdjHGBKi6FJrZdIlOWwJo5aQe+NfSx44d1whhZccOE
NpFI3RBZCEcGU7MEaaTjzo849YQYPWvGyj0f0PxqCrh1epS89H2ULOQN/ee/dOfVO54qj3wwzvRm
M9N3fYk+nv/hqJyNozfreo4kjQO2uzoK0Rqs0v2+0XWYIzgUxbFj0hgX1JTtiRkbXN0stBstKxX/
ejatZnIQVZiOlNoIlnl1dYF2x2328HygVcJapxGPQsLk5AaCv5q9kEtN2vA5EtlR6O4/ePkWE3Yo
lg0jgCdlKYjbwx5an5ML/Q/C870xH3idsexZXZUpSTG3P//uxt50li2pSdFI3tUA4XzCIUWmAnPp
vpDBch66G9MB4siwV5fkR8iihwDw2ZSBp4/VoGTT6KPNJEBmmuHLp6MJL44xd3TrNTala+P4TETx
8gP5gZiHPlKht5jhsbp+j2WsMvNgZjVuQN1Nx7veGC19efaAOIMZc7PzUfBGhkINHMpFN2LynGNV
tN3GABi+MJPem2DDC+P/mnd4N9eJbc0BHmzCeVPjYQJiEGnC7CyF5AN2jbW25skPuqjyfh8afF/o
XmeD24D/NBdnZHDzMnYaEHg6YqBGRvLIZMxy83CencWPMWScqF4oiKjudGCFWCG34p+SP661zNGb
VT/XOcqOA9eWVfFA8nPfnI7I4M6OY/GRxZO615QttPXHoSLIWtnLFyXaRE7WTwW/UQnOT/7CvU2k
QbmS2omF8Jj4E6E1XExOkAxS6ytjzGA7XvhOnfFc4WHpkQZyJNaLHuF7wQ7qgnt8z0UsntqQqiPC
AP9B3yOxdoUpLiXjdkAPUINcfyVo6HsrFphDIl6Jpbdx4mjR36RvQl/49eoMhXbOl/AzalxtzFXa
ib5cTK/sts9T+bJa8p9AcRE4s6ZmM1rYLO4u2BDufgn/jsIhLAOwh6qHciXvcolZXsIf0sG+qtvY
FvXVMyDRzE3bwmn6OA0dAdwvTJMZ2eqU0/z7d4XlvC0UpKVTQFZE3+sy7xUXXyKrGoZraWR8EGAT
ECYrzlBB2rxlEKYrWazX2RgrZC2ZKRyAL+9YWkcNONUqVLThNb5N3Tx8DURxOh+hpCDnJ5PektyY
WWCD5mtXQdG/Yml/Zf41lUGPljcN6UAxUoexPusMq0KqElf7Sn6TRG4SC2Lm9866OeEqqz5TXolY
X51qqfjP/Nz2RP2E2jrbtl6gMpDEgYZrdih5RwklkXSgNu8ZxJpVSyQHocqpkAI8njtMhp/ACLC3
jsHDNU0Hrl9qZkAxcnhnzA5tsvECfOUcPPxPKmx7bPAUORRba6hpYwqz5CxqwL3j4t/AUd/CDYNk
6N3GDvsPRYAW0736hpER0G/Bl/bXnoVR5fWM3PSVyIfrYGwc5ikkqIO+3KNfEjFYk1ljekO2Tmgx
fseazxV6tzRz1kX33UGIgRUyoBJvh/hn31NR+oBq8V7oE58Qk00MKYNWWg6W7HU2yTsKzP4yPQ3S
ToiQDXrezo6o3SjcLqqYVilmpWYdNJ+wzsUQyP8632ZiusA/Y58cmq+pLzpyG9C4mAN/nN8khoE2
FX7lHOsNPuJEk4NMqpOlKU/RAV/0dnYwhzAOdEyl7+AjsnV7YIdJUWkntyha3AkeeuzXRKS1QhX+
N+eYoIZLaV3O+F1Cl8a0C0kPdeii3DyJAUWurxQfg3Ak8W8N3M2l8FEoMEeAHr+foSGTcXiieWRW
SMIHu+HvKaFcUnbWjznwdyGE55IcwE7A80zfB/ZH5gR1q3WFPhpp8+qa+RIFewgEptquTyg+vyXq
AkgaRuA1DJWmzRQOsjXtlm1+N05BG/3jA8OiTHY3igBXZQs/HhkCbos0DI7PwmMTbOhe1MsESVjz
UtMS1ur6X/gJL9Hbsp3AAW4Fg0bgpHJQoF7dcQIdghCXY5VxWf2ABEqsknHtBqI40UMi1D3oCW9J
bYpEO+UjAqiyEmTgyyEQGp/NBHymVtQXY1/p/w3nogvALhkUvVAI3WYgZaA1WLxTZPfBcR0sl9Ng
yKNYAAgoqEcrcKDmvG71WP8L6EwTIW4Svk2izN7dbpifQemjc4rW0kHVyZp5gGE+WnFrhcU1h0OW
4V286TTMk5w2TuXYu3Ci4NrKpYike0tX0AMt/waAhZlWuNCt6Dn6b15mPAER5Tk1psVxMTaiDLQn
FCFdf1GCglMVzqLdk4Fuqa8TYsOOdW81uuamH9565Ew53vNQvaxFyLziakGRU0pC0aBZrcQa8Ksh
bRfeDNHC/KqCR8Y00CWO9ek9Tb7DUq4/kJRtNttwUv11GoaGOmFUw5ws8xpir9HIgjd2vdU83XLd
V7b++k/iBHIYwDQIJZyWuYx5hI4sz4lbxENn+qqIrHRj4xfQLqz2lzv1Jyu2kdCCg1l424BzRV/z
gWL/Ai6B/kry3R9hTm76yCRp6ccY+RM+JmSo9Xyk6532Sf/PGgL35cP5KxhYTjy/aN/jm+Ew2vka
O5F/6gSMNAhM6vW1CLukeF2Cr8Tvjr85x8j3A45vk/aBFtmTsU4Bh1xS0qXz4GiyscdBJqwSooOo
Rv8RbO9xCNbs1qBSt72PASZJo7qisEnepQNAow/gUi5X/mcabccB9X7B3Pw+bBd7xyUu5wEDVFZl
Fcq+ysy4l/Z870jdi3XfRDFiT+rn0PDXhxPRdAQqBrVu9dGXGJY4J+LecuW0yKHS1s23Twb2bBtQ
URn+H10UC/zkE2aCiTZRt+7T/3RI1DlJcoeCL8yTHHb6W2uFpI4WTLO0n+8JZ1Zjk2xT1U5XSggW
HLzPC5uVSZSiZg7II6PRkAuvk6lKRwUl1Vi+PooPyIy2JWYHnblQHJbu8wDMJJMUOYUkiZ4EiEmQ
p8gN6yTTlKFPOT47shZm76Uy4v5tV7SO0Eq9EXZCi4bHor8uiBZZ3RNfpfxVCiRFnYJQBDhCCami
iR4Zewt8CQHe3ynfQLzMRIcwKJ+mSOgpYMTjygAgRG3Hur/YffPRorD/FR1VIgJcP0VZ6vD2Te5T
COFeSnEIXK68ya//lJq74djWf88EFO3obsclLlELLlphOVGyDWoXw1DSqSBuX1K8k0ot7hU66M/D
cB1MTbkNuE+i3kM/QG7BBzZ7B4WkphoAbOeAam5hyc9149hSS0+4lBpaTwcoFt9o7kG6JkOPQ07R
giVt3B/7ZtN0NPz2CpmuFj1AtnXbSJ2WyJ21FAPr6wqN/SgsEecedRDun6K1h7w04gk/39RSaYEw
3hBeaQGq53KuP/6J61qEpZcXE79vRRMEKHfjCwipP3qKgRjaTlpBtYzOs1iu8gaMxbFL6tqJaYpN
LfHdtoZ5nEw08VGchGqhTFP3aM7D55UnopAj8YchNfCXzcBKtRb3YdMLGK5/0iaKlZqu0b3Z2/iV
43yPWNZgbNqsUtYYCvbvsFU8q035ot4O+nkFJ+gnHQ9xHxBfTH1600XtWDkgFLA86IojpZLo+3IY
B9meuee7LMTE2+JikzBAcTAjORUQHEyZDwKHDEYYi5rRlL6cXXD/jMIeY9nbMCY1ky0qrwJ7SZcg
6W62hfTVVquThvFzkBoTOUUe6aZZ/Qyn2vS0DFuvS/WjS6EB4HQOTGEqxewYqQ5VCFlmmHck3oHG
9zPwuDYwrlBgApEpI4balfG9bu0Im92Cg7GBd53SzTWcyX2nT3sQO2eS6KdcuoNrXgiSZK454NAd
MLLxU7i5br7vkVpz0c3Fisl5xGND5lBpCJK4T4ipmmJb3Q+ziAAQ0shyACA83RHjLd5LTlQPnNbG
z7Nn39BcXnUFbPU2g/ylotxqCEVMy9H4BK0WBSJu1Ke92DLlzx/WzPclsfyuMoU7qie/ls3T8yIB
osJVDCt4mZyBVk/nR2Rd0WKz9XyuQN9kG+ZVHEpqgOWONgWQ8myN2eq91KnRtPdpmIeOfeoruJWb
QGJ87h/N6E4UyZmzfe8vS1lY9GSiDRubNAp6Rlx6wppgzm34GAfT4b3qV9ttEqas/UDSh1yps9Gq
gxlXR7LfNwExubC2nIOZReAxN6ru78N1NiH5QfbbPX4z1h6h1oFiL3GzYB1xhLh+Neivg5eOq+a8
pUeU5cE9mVY7gTieCsu5xlR26HHfOrpTfmgaR+Si9atv+ddEaB+DAw+5M+UnhNvhc5BssuykAMHv
Gfy0SPbm58bojCmYW/CfxMMHzl80GpJRn0Q5i21TyhDIbVY6USKpBeOqeGpGYzTDymNe0kr91EwJ
lj1mkljf4XND+MegdCz3p/9O+ikJkBfcS1+Y03j5HsD7VcTTBWXoKt2FprLxVeRWqUJNpQ3KtfJS
fFQa0KkYenEhy03+9LnYE90K/IZdwmTuQRwJKTndFuzhprYs5m7ycNSso/kuwFtF2bMlS20FjLkV
dP8mmNIixt68Cta1NogQYDbjGs/riQVmnY7lGdpNtZ5astMQDjhKMAC/71KL7+C6GJ5xcyyAm97A
xPhMvFwNXNS5PXDD21IqMeLvEdL1C4hgnhl7JFaYybaM+KWG3LA0hjp21kpUP4h38ld0gkfI4Q8/
m3JNDrWXMwzGKTsqXMhITQdsEPm4qlQkzNvIBV5Cl7ZhW73LbfK4CsL8QtJxX3ISZKswcTR5D/IY
Vxf3uC6nrrmsST1wcSapQDXfqBL5GV+f1IlWqq7Nj3MjNUX+tPgzwhEHVySFZH6WVBfCm7RqwXPx
xvMazclri7ye04ZKS6/zwqeNn2ZpwVRf1rhp1gFPnbqatJLfQiZxv9+ce7RuHSE6vgi9mBhiXJbC
A1SS0Bx/0JbhaIiGmIOGYwc1XlCUTw6j2Ap6jn337ggh2x9UEDxiX3ejR7vtHlaw4in/eJHTpJBy
qk/sgr0ssEIgFqev5XwylgWY16Llfhg9jlUqvrQilMsY+M+22YLyyRnVHPC71v/MfR4Oa1aKgfsh
9zE6Dz9irnklWKH416cxE+vRb5nYrXd7mig4/kyit/BEJcRHC+tNDO/y58WcCyZtom+bY5UalqKo
QYPAgd2/l3cGc8MQLY5uyavzrvy7KCQyMUR1w71WW9LUqtq4rU/JP3cTLviCl66opJYHIoWloifQ
dmLXE/l8V8DIFObGoK31d+VWvilMosBZ3NQsCJvL1j9ipL+Pj1IGox+0sADWXXSWnJwzGSS2kifd
r1+y8RJO2A3MPgn+ifD2L5cLZaN/GrW53w+GEd7bFQMydo1oQH+d1AV1SrQsAy1/8/OGoDi9kLPK
5GoxJOG1CbB7MmqfsZRWW8CL3nI6MevWGOpbbVm+UA/4Hppc9fv5PwgpAWeYy22qZoGne4+f+P7a
pGpdeXNQxVIo9yr5unIOrLXVkiF8wRuDVBGWc4LeXFtSi0h+V3QYGSTjpZNwzu5uUU5mMmk06UY5
nEdN68BVSBSaYWEOMR4hKcUZ1olLDpBlubKvfVGBjIWwEgyUVxFM0HGyXpf6JmRXNnbYsl89Igm2
pusJ1I63kYGNqLGdUq1PcMb/PAVWMQXnsCnANIMp91SP6S7YxiEuuChiYDCkMxmx5IudaPWpXyjC
nndRS1nZhkKkvc9dt5F5nUzcJgySw4s7eCqTAL8aOxgDoUGBn1kNP1Bta4DVDLMhf4OECf9ClBZp
I5rRD1u+KF0C+1Ycb0vg2DFMmEDGcAXF3kSjIuxcehA4N+Mwu1Dub4W0/8MAeMgA7Xw1DOw4JvJk
K/jSvNLPgstCq4CQebGCL1JQMEECzvm/9K9jS9TPEpFz683Uef+2mmnQzkIYxdxLj5nyWC7/+icn
8KJFZxSLYdi22VZmMU+MtsCddy6uK0sr8Q73ACRWNuQBd93k4KZnhrrGNUGoo+4lQ9iD/EgzmWA3
CPELPRP8klFA/CdISqcXe+cth+tH/Df47n++T7Why7yLNa1YrUUc+3FF2wUbMBxqu62XfMrbgqyU
H3IOFnz5YVcE6GoQOWxz+bFZFm7pigm0VT9FCkqup4L8Tmrx/hXSQCkkdL0C0eLTB/QrNPqpCisK
6ea0LVJzm7AAkNZXgdz0IvEu4ZsXX4a6Hcb1UToPHhFo6+25njXeNQrOEwvvK1pgqWGSL+U7cPCN
kmubuWutN+isH1E1ks2h0bY46MnOHPjaooHXktoWka9NRCdmJCgMpgy9FbcNqsq1MfcOsNpET+Gl
/vETkEU/kUQ1giuehWq+8JcHNfyYvxqZ50EioG7tPEJaFf5Bxb7S+V2aWW5TPsfeOVQ/zeoFPdCK
5ymCDD6r2AddQYX/wWmMWbMNObdxsoUmz1YoYHZHzNbw+zFlqGDc0BoEzaI+dMftOLV/KKW5BGt+
tm9xDr75lGyr28foOGQoWweHQYN4jnXERsn3S1RhPMQX+S+uKmTpIizWeXZ+rTCIn6m+ra6YDCqB
GZCokLT0aexAxXHqPwFu4tLH3yK4D7pKbHEDct0/SXYmc25IV/P4QXhEeRRAN1dy3ll9uFEXKqrD
hj8xXZ30wxTVDe+fBarA81itCHKfqW0pghZ+xiphj5CnK+vzFp3+TqS8K/WxhMuGGb0EoUH2QGdx
MXS+hmXAmKby48v/Li4El/LPgrCR/wreiAbYRk3MBq8s3DlydWenYUPZzokwlacIq8ZLYE7Phzxq
oFxOBv8GrMlgV2sC85wcx4qrj+ltuqpKGecd724VCycOXA3bIQrLUMPeSlsbRdOHbhHk/K2OsDga
UtJ5bFsLu6EkUsnqPXFF6Vmg34L9TXkfIGMMuRboKhgD1V8Lx35OLstc5IexKpmsr31yjsufg0YI
jE8DQnKVA85msN8M70d5mmW/rkeb5Wm7XDemO+kqZZmhBqWTfB5wItEcneJU1iZiP49PzP9ARXoK
BFnCouvb3z/VoYDm+TItehFzAbW8WnhNDVvFmLIIV2SmSOjS+pDHinHE9pKup9znmElvewwx8bOI
Yk/9M2tY8ELyc6eieXLEqqJjdnWB/pEMbS3ejxGTYeIMth/cK5CtW9WBHOgwH9Qr57wEdYi8RpUK
4AmeQZCjxYTlWd0fF5ZBO77ZOePx1+56a+RoEwY06K1BdCskAm+uF68p3VOa5dYFmyJQF0eX86Uk
4dwZnUYekxmJtrM3+RLhKDZJ81nG2zVKgVs5UWc92BMieAPsCiJy/HSNrGxWgmOgFkOtIUa24CDJ
Jz20mevqCzfDtjnDOXO/Y5gxiPxNLGouzTB9+iIU2ysb6hsBzBq35PAP61L2ofxbwtFtCQSYF16v
6WgvXjgCc6/4tdpEodmuXktyMW+5QnbxhVe3y4Yr8dvreeQiZheE7bXiScIKCAR1FdSG3LfyutQ5
2O8d3nb57Te8k+xBNNlffaavvhk0RAqlpTKYzouRezTcKh6wcureVddKuxcZ+RS9kNdZtHCUnlpp
SoFiKOBQsIrk23jqcP7VCHalr5l9LuTHMlykKBmbypzSJ18cXuVc+6L3L7RVv5J+Ux6xNvqwDsjW
+635B5FiiwDMwm9kUmXLy5fB3S2xBtLM9gTmPqYU35LNLHYtmvqCdc5TMaBcJFMl29DguCSzTokJ
YtPb6D8paA70IH9xnPbgcYhCxWmEraV1UgMEnxhIJHtVJ9I7fO+iMpKzJO6an3Hi7JIvCBHe0+Qf
HP0q5MTx17wwcV0CRnTzDqzfuwAzbLqgIY6Y4872JhouM1UeVRpr6rjfp/MkaLgpdIZUphPcObmH
3KW2j9vC9dQGXKHMb9vEbgY3SKJdK8xn/T5NtoTzY63WyXi4/WcCa+Ih1G3wcSStYWQdcbwukO/E
OFnb0GwU+6pvK6kN3lB+1Ae7uzwWoM70RVLqPqKRvs85e9W+MLjQWcCmxb+z7zMzfFMLfE360AYF
qvYFpSk0BbXXkHgujzw+irhr6kcqaNK/8exd1CZodNfqm5j7AXXvPNFWC6/6APudUHootIIK0jUw
DF9L3bxsABLwtJ5mopk7cRpwVxEm4B4n2FrhH10tq0Mxgpjbzc4VNZGtZ6QqNFVRhgpp78rB5/YR
3A41EC9Jm5hIdPt6LoANC7I7C6ttuEVWqW4r9pksP53klevfV+8XgDKlhN+43AAdyZqZ4E8u23b8
ngCOFllL/QwH7wETXO3wzrf6smvrQcyuWLzY5n+ct6VLVcN/hdnmZ/q58d+KSUN7Tq4nYAOh38By
zYtXe1Ews+2OZfT7O7E2uzTU+eKy2H4KH93ZgFDVTFI4J3hMzlQn8hbW4RNRFpLTm+DEGCDiauha
8W/Ihn2FEcoLhS+CPd9YSQXzZGKq6FniQIImxJDXyQmp4siTlMdsFvdlFXu00OxQXgKoF10OXdq+
N634aTrBpBFn7tcwnpijBe4yJkDZolJs0vPB79OvoJu3k3PZpOvEPNeOvnqGxU7PqzTKXmDJ0Wio
O+IOlEwYH08Wt5mnPYBgvjZeun4nMewrC1HlhgxHvTmZgLFzLZHQ5Xbq/MS+TWtOr103ZNso4983
Uf/O6DBxWzK3ZC1FGUAwGmzotr8jwpd58/koTt1WYl1qIRel6+kmUhlDgG4+qmh0NheNlGFTrzDp
CLFzDoAZnj1w69/tYIdw3k4t0a+Mmb5TgTjRTCIQC10Wavj4SXKBNxHSBBDHX+gXQV2oHnim4aGZ
USVcGvUA7CRDaPR5BHp5qcCQQQrHU0+XGZEdjqJg2M//Jz2vwGaioQFBP7ydU85s9Kejl+nkHKpQ
JCkbqpdrFfu+i1m3eFKKTCSjRTeWwuAqgcBVxxH4KbIQxryBBN4zteGmAC5aR1jVqOzsVbY7SRxg
RSlHj/3eC1YAnztJehuiMtvtwYM7/tFmw6ZcyCHcJORWsHQexvFD2V7JnQl68WZ8sG50+8VM3QYu
sIKn2KncjXGQzlKpRIHwIGxiDriFUlIXDr9I8YyHnYd/BXMPE7utHkOQClEGVK88olOa7UlAg2/e
3Fbl4IceT+kXhyPP7A4MdZS53Sllexk+yKaE2K+J0Dpm4OsKLtWZwlU6ri1JQFwBSPA0kvMAf7K2
0FSTKXmDgIbu2XQ6NTu/cX9OsAgsuUfUEXPO9pm3V77eDX6ctfsT7ihXmluqsG2KwneT9Q+6KuwF
MhqrnHxAJMVXjlGSxyJQV8s7VTV4D50cWSrbNc/UI1Va8YneQe5jw/Un9iSXaSCYUWA6NwcQcPQu
Jus+eUt6mMsPAmvBiwdGFkJFwhbqsRksW0WkrvwEF9Ir9qbORcPJCobN3kZ77EaYj2XQfA4CeKoi
bDKfbw2M2YqbsievpsRpw6RRZIFSNLFVZGX8AsHHHJatQdyGmlzBX8Sh8RWckXkJfPr/xLqcaNaf
L1im41MHKY+oyul/CgamD5/maipsHBOl9egiZVDe8Jl9xNbzuKjmvInEms/3nQILkc1o2yuK+ZFe
PmgLW3Y2/i/Fgz6F7vXApibCM2i3gIcLknQZKUQYTQAvbBnFJZZcq4KG63vPJ1n1Tjakl3tQCJNC
mei6b4G30UIQif2XtEuN/F4ytfApP2h7L3oEyLR8wpkiPn49FiJOhpBiKU82id8caE2IbslmJdSi
eRfqiZ+RzTXVrT/DKEAgXKumvwebwq7SdpYuMyxbmzfEXmYQSGOMglcMXjdAvrfM08eXM1/VsQdJ
DCrgEOSBGhLbsVOG6k4rIb5DW5KWxd1J2ppz0PdAWsMqEzzlg7KetACivd/ZarC18UHQYW2SYVCo
yMX70X7lkA+F7kjf8sojCqI5LBTMMuwWVlmJtYUeHjBy1lafSAp8ZmpOGQ+RtpvTHY0Jg47ued39
0Gd1SIkonbhNAxRed/O7MN6r9wUXPLMGDtNexCNrkyAt1wGykRdYqOgS3BpQ0K7MkGFIn5Le0XOQ
Gup59L95YpaW6kParz1s7w2lehQRnwsFZH+cXIind45U9zrXB/qfeY1C2j9aOPSWUVBH60BBLs5N
6d9jWX4s0jvJ6z6faa5dpX3p3ERcCO3Y8Ar7HMVoxhR0jbLBq9HoJm1xXxrdlNb7KMiSVkE4wSv5
Us2Nei268ldISNsERcX1fpK6cCjsYlW1zyvvmwTvgLtNQn1GvHrMm0iYmPSzIlWwIrDUCJ4hGYDN
JBpe09OJQ5uQjOGJI+Ehn7WL/N2jq/+Z+aiKcwYycLx/qmIyIyQl7ktBHuCdK/dImC69ooT8UDcV
6NmK/wPoXRwLWbxc3Dn3QcDqD2nPa9yB79iIldusYbudZy5bwR1HhrH/AiRwYYsC4sFmdbhriJ0w
VHvcge60ljk6PIY/Ar4Iog0q0BOdX9S7/W6s59tolvirjWtma66nsNDAVfTF8j9Z0RzJMkWxHvqg
guCtScwp9mfB1HWm5D/JYuqM/EKGh15wdBVsCkdhqEQj9AFy2Hac66vfRMPPqOP3f1e5cE3C7zvt
GbAGf0CmSaZd91/wpy2aeweXywor2sQwgKDeIPq41WDhyp7QaxiDq4ipszbY8ApD4emIYnol7aXG
yJ2ZGbnbP7XRaYglMHpWFNkHjxDJZT/yR1HtABzYjfrifOo45WM7/F5NvNafaAwdxBXGDPCOIOU4
kb2AMZ4VTl1ZVduNOGLHbKGc3dd/vvsXO8P2YWB/9SR1+GgelU4SFG1ifj/Pt+fwczCwDLyycLvq
XMQ5yCw4d2zLG1DhGFmnF0EMIoAfUpIPOOM9TjhCoSkFYotrcDvPHNgxjS7pREPY8sIsf8DebSMe
mKp72qUPWZYex8Lp0Hi+m7o6ieckbXUTIpNqw0isqEw/UZ6Sv0/BXninpD38wpdLemZw/803PiHi
KGYqewiomKZ9zKmoAjnf8l7uQ+iZBq2pTBYdf8Ck51zLheQGN+P9YOJJ974Bs7MKz9RlG6dozjIT
wSDVGvN8n6WMuuBqUqf2jqXymyiXnCVquqGcca7y/nkzh9ZSE9H838aLRc8iDQgcNsEFDoTrR0c9
m8+lfTzJJot/r9qm/0cYZIOBs6k1iwVgLe2oYJggFodRSIAMCaAafoEoD5alB0l5VHu0QElcvXE9
EMcnlUTnLSOLmvace3ozXAXEm3sGVxZ0KD2FpCcSW/q5kSsLMtJeQBczOGiGh8f+Bq3XUClQ7xMy
Ws/VZITIRljomK5hpdIZ6tQPnUix5ECLfWfqtVxkCnc7DUWeFEsQdo7zMYLj2SzwFlp/LxuB12Gw
VptP8JStChdH/OAPqO4Q1ZOduvszrajlDWogHLfTwMO8Tb3jf2oqR8NTO8/JEuKYMxetxwuciPVk
IkOj4RcvCcLEkd9o3/Ua0vX14t4YctSfLX0gQa253QPP/2DX+44z7+nzoPud6hvv56mDyBRD+rTr
Hdmd3lpn9+RxCGbFpX6CryQZxMp+yvV/te9Oq3uzrBnek0Mol7W8M8jm3Z+/Mc5+lhKySVhAZivN
EeRoE6HxFGv47RZ94Cn3j8w1Nr49x6ssp4nKUm9t6gFGV9HhAtXHn46SwxOxVud/USzwA8wdcOtq
Z/6775hmsViDlLIv834wysQCd+NurtNIEwT5Qs+1BuOND0pz+CuyUoHrjUqB6koIQ3V+zZITU5VL
feHdkY8nDc/m+/GqUarMvWjLZ7vtNujS5haUPmq71S5hajWyI6x2NmXVzCKjf1nxC49/8s+nGG4/
hfAj7ZQ830VdPblTR1d/Jytv5UwBvaFxpMqYJZD/cY1LzybViadZYZxw9tiL5g/nHzaFZDZkR6Zu
OUbgT+iy1wrzZq8M1EeVdCXmVXYlRAncGtY2f9U7GBE2mlGAEcQAu83y1nUz9apRKMt3cK58HJl3
oEulsbOLVNu4orkvVkH9+wl8hebhyifGYJ7NnFzizw76NZpUeP04jEKoqJD9+5qptp9WCIbTBWR5
XifSinL5PDlOIE6tpOXk30xw0wR/rALXedxocbiORVncbvazEM49zQJ6knPjp61FFXXZDuUyBWqA
utQiQ4VRmfbt/PR4EkrnnoeXN7Vbsji4guYvEQlD3wI0/8BFJDD8JD0dee6MICr8iza6+y3lzZTg
IRAzKDzBWhGq43DHpuISzp6XXAGiR7g5l6/4JiSr1DlW+fwiwnx0B/z2fWuGLwDXOmBwrvQHNXD2
P+QyRrNvg2N1RyeuxU4sMN1AW0I1GimoPjJM9lZim7MOqUurbzQCgyjWJ3YBiOWeJhhbugufSdr6
Zw2daFTmeqWZoMuGPqR6A/1pjGOcZkoGBxFm3MooWPN0rznJ7Jop3n/3YcwPQbPosI9lyc13JfQk
/dHeYmzr40TCbwBxAmTMiKiBqonuTka8Zs2Rmoa38mOmA4k8dyiXpLQ29/jRUIQUQ06e5pkWF4bX
H9IP+jJ6y8hlFtycTV9vEC6XtabuIQqlZJz/M0loaccD3Fus6OzOkSKLp+9oRcUp7rzuc5monma+
c+jl4xbudC/sjFN8Vibcs0Zkn3Yc0mLyeP21Uv+l/Ae3hBtmWuzKGw6dSHP04k7n+C+3YtSxf3Yf
fTVJLDqCJxEaI3qrwDQpPPLkSfE2rR89ivx95hDNSsLoZz6HZQ7IaSrMclUZgsmJDq4V5EV6isBN
QDYqoWfPvDTirx81+8gr1gXR9aJtYRXQ5AaKqACwLI3A653VSuBC1uiOQKj6fkp3lU4wAjJBx/oJ
OgBs21e+QVvCpGa7RnBpEwG9d2fkTaMtm6khzjLJ+Ym45pj9ID4NHdzXJ3Zc38DkvqRuCcCDm6As
TVftMkwoD8TPCJPkbud0ZUHHYE9eK4l/YOMKxnoD7ynu8iMjLs1PODkqMbXcJ+gBDI84HhFOPQ+U
2tBohR4ZojRotTVvP3SfK6aH1tfg4YesrckvA2nPFY+tOu3Q+8CWBT0J40MsJO2opU+FB+8TpOBP
dCL3z5M5PPmuzQnNDyL6QwF/Pu3FOPhESMVQpo77Zurcijg2XA+nkH9nAWG3H0HxjnynCOu26Qqs
eRitosluj6++nbW4uikFORVbnJPfykl+jvNgSUcIyfJzOjvefo3Fxhtag5H/gdskNRFRcs8Qruz9
KW2pMcSeu5+Vdh0zBOrZs+H9WzUZ9WhhACGjIunHxHWvwGaXpwNPfCFYb4nMLE3H+nLEoPiJ+Tcu
ViWl3Yj5HrH3/XQqR5Fon8+zB9BGUudGOWiZYvh7WFqy67MYXb1ozoBbZFMfBqYa2Ig3TUpVVItU
4cUtKbEASz29os8QvVq3JMUpbz851CesHUHgDuX/kcYIfb+l8lPNkVzujD0ur/G9mQ1yL1FWplDe
/Kdr616aVIi7wTqlL+GOM4eFL3qaqqNmZG8pmXT0eSHBnPDpMy3uerKi5cerga4hi3tj/u/DdC05
EBZmsbWylr+8xchnxc4Wj4cROxGVEP4wJFR7QBu9QJoB8smb1Irt4BVTGEbik/9zuYwcQ10YdE/i
ME+G3i935fuuuKiALyVN621J/FhSKYD5kUUmLJaNXgKdW5MVZd7dvyfIfkZt7RlgsDpVZtgh6q3T
th7HsMNH0xBPKSYZOPdoo2FRo6xMEvJljifgxivVUCe4G0G6sPzEnpWNsILYtOS6mOwNH8CuAFWS
uFUURoGtzzHz7PkeO/S8JTRrkF5q4D0qOASa7lrXPdXmnJYQREpDPH0Oi5J7+K90cdiaiFGTA+3f
3DbJKGSuo65DA1krluKUbkUcADAW/XV5F/EQ1SrWTxnsb83aBbzFU5RTLz7bW/0PLyc2lXN92B34
CQBVLzB6WI+XpwhHKVtFeoeAYGdPbq46ClxdU5Ml+L85u6NyjeCW5bKypRH9epSpBycwZmkH8LXJ
YtyL1oi3GwNY5wyYINTOPlq96TC+VzNIAio0OpTfgWXCFwKIieqB49rahOSP9sM5mh+LHVxU0F/c
984NstZEig4vm7AbYzNL5XbCoMcc18KH1VlKoLVJm4IKhqmwn4q5F7hHvF/L+qDmPWVEQbeeW3cp
yop+jE6NKU4GYxZzFgiSmoGrrBhD9I+yua7QzG2ZFoORXRLiuaEWFgB+ggbGxFbSVfV0+e4h0ZjN
ZIlGh4uYaCyrV+2BPRsdzFMvkoxC+gbEwfOu/QmOJdCJ14uDijrVbVpV2dFQiv9ZzoZ+LYrIiX5I
ucCeBkzbMgfSdbdCqKmuT0OXYWLh3rWNXawp8w/7aMFW+MXZZS+lcpMey71PSu3imaJv/DNQB1xA
6bJfCpeSfeEPt0QFtZhRRxhwnVhUm5as99ejCeSMwpKW8LnoubZsn22j7uPiphU1yfVR6cRUr3oB
LgTkJzXPMs5/yN4javW4nUmntdGk3L5mEEkYIrvIdttoEAYVPMujRm284zP91y6EkZZWoNHqXZE+
VQ1VOY6cVjcQ2HWR0z4bPvwBtr9pKKjDPZojsAehqHNvRXlHdWHaEM8sE2qf67nRVwzyeoff4XGN
LH3FgaVLvWmsd0GWH6c7G4HsdlQexF8QKTJBu4+7to5Sh780enJF6tJ2DZ2FP/idC57FiAgd0oyj
X/u/eZOZ+pUS1mIrDNvsiYeVsIgBtCQ0nVVrzVaTcz3sykmtF+d6piIpOpvVUSOBIc1/aLHVm9Uc
LMhzkl5/9TFd1XrH0bNizBuGd1vm4vYk6nZdIU6B/9rFHRlCZoTayyuxhxGSDB1EV+h9efbRYVO5
YLsgukQwS94eBluG2jTjEf3OC9pfmvC9ELTRKiF/5E8t4+HObbF2KeSc25h8iYkm4dNuJxnzNi2V
9xWCGfKIV4KN+dy15/G58kB1gbY+d229HX1pkgp3xfml6LFtw1mxcaB9BS7+VXu3v5lFNIZMWuFM
iO+cHEkUao1KC1LLQB8tcEyI6Tb2lo1rCMAXGnYJKHpk9JF2fQDPJoF0W7IcmYMsvMnEMtK8mY9/
55Y77JgySf5fNvceLm6vmpUzS1eSzH7tcuAN1BUOe8HMs0JpQnuWCuYzTku9+AlMFULbqHTw7VMk
+MRjU51ULUDYVqz6Mo1DF6G4RhXAL5rf7hOym82MBOi/AuVnCefy21lp7+pft3F+g6Vwkmd4sv2d
ESeArYrSuAM9SIaYmS7+4JEqekL+cr09GRjl6hNSJ/JUaWOUQ62fs7nF7wwn03z1+LQJlcJMcdg5
JTbo+7OGLley6AMFz+MOtQ3JAIHIL/VWFSpRrBD9ZlyF2NjNZkkYJtxLWIR2fiN2hLx858Dij3V6
wirhZk8f2jnQ4FlvPgxX1qqUJa4X0jmF/q1lE5p1FRwbY5TW6I4DB+6FyfItYZMNUKTtlQyX1zYm
Ienev9Exkrzx5AU2o/zwAkbm+za87NDE24ieqsXczqY0bLJu1X8PD8w4Zer/5SyvJC+VvZ2/UyY/
88IQLtdRknWwAmQV82Ukkw3LRFloFScyPXhgEV2sAtH2zgSx3aiwqiR4XidzGUINZSS5Aee0bSqU
FccARd2AQAfG/6gX28/rZ1TBNOuyTqhgyLukzY4vWBMyujeqU8fpCFDdWl5kmvNojxYBdkXHaDB7
Yuhq9RoxUhqkO9Tne7wUvIDpE4Eh2YG3qcGaePKBaxGMBYcr7ZWKBW0Fu4WcsfGaMahEyj9pcILQ
BaSbWRDy9LCAUHcRwoI3ne1OzCLp96ddufQYaAb7l6dbWI0iwsncGIZWCZfIM49BKAhtfNVBmZcv
li/18Bf/saz51SPSnWaQD/yE8Mhh35DeKpTohtmOvWmySfbxVCToABz/Ewu4AyeFADldE8Zc0YDJ
3SqJf3MkPdnOPxVMfz6H2XN2MhQymJ5vZ7egFGdwJ+QAfEK9tOw2TkbF6qKJltWyYGryoeyGjNVE
ulNXkbwK6xZ40eBg1WEH1eTbnHNjz3gvquWbg8sPf45JjFcbaGazrKnFlzc9tf7OWs+Aa9C9lRiN
aNxHkzlmvFBVgNk9UfJfkUcN5VUQpHkpWRNVvgEYbEOaFew3LEypRlaEEbFfAnE7S+H3ePY7d9DF
c5GdtCrQmKIHM8jHKIOKdhFpozB/LfSOsw4Q2t0QozL1VgDPAyKOKAyGurElpsjfmdfhrXgRkV08
GleEu1dbJax2SIa+fVkre25vAUU55v+5HAQH64kvDYAIBApFqIv+RO5C3j9vgH2CUFDCK9yukJhe
ZkUYUWV2ME7LOvJVX/INc/PFVIShXn14cKYX6cUdqcJhKzjEAcgH+L5kdDrsd43Zey5Rp/EGCEht
kBL4B5bPuao1vxRnNaB7uuEs7R1FWgDt8jPiPuU4GcEojQdkltbjE9ITa3zS+GDYkAZGE+9P/J3Y
a5l4hG7h6UwiJZnmg4kEI4WzUmFf/qKYGaO6SrCpBvJDGqOQqx+c2Vfqz0OBtYj0c8+l4390R+zh
7xE4GjOEbun8BfRC64sDTkPqkSeOhWeUYIHycpci4XLnE8txG7ENf9mDVnKyG0KTBnPKs/rA3rP4
SnBRRMesmjG9992GoqHdDlc+JZ7O8B+DAC36hEfGBoGiEERPongO1BsmGXy6k00ZmeIXTwIRrbZT
IjYKGboMR0MIP4pd0NW+HAO9aWZZH9m0Dz1B0AO91MPQxgV2nR1CLx76BKs2mKXDfWcXWB6e+zIv
wUC8niSt/FO7Gd4KD24fZBwbbcLaKb/8WTdaZ5IvPWR+BO1HW6MOLOL7Y7Nk38vkjQLakgvjA3u3
MsjGR9R1amjnw8/1wYpGeKJqJrN6Qi+n214fJaYLzLyWRB2HZGA0YrCkP6Gs2/wD6h4a6SVtbCkI
dpsAQQ49+Oq0T5QXpHnIQprUVKDzWfDIYysCMHV19AGplFaJiIa8+17H/pJkCPUhyM74pSELh9BP
YOwdIHEkg6xitMox8suuBQBY+ioLUJrJ8el1cGAfXVtRws3ihdEQYIRx4KLpwzGzMvNTvkXPXxYo
hCHPLF3R3Bg3C2mp0uVcs121gS1xvlwvseRIV8UI90MIc/zI+8dxfNo3JZcoJZ8lXla+sH3q+K+H
hXXZOHz7xTYSeseTYiv/N11fxVk6MeLuhyldzOJ2S/CsZF8xINgkT2xHsZbZdbrr+Hm6I64FGXxn
8vh6PLZFYanGvLJH5KO3MnH+R7rleD9yU3cV4qGhXzmJmA/iuycOjb0A5RT7bYHgePUeYUz26vU8
04ilel9ynFax1UyLh2fbs81nVfXtI2Jpfsw2sYKF2a96VpWUDvCyEEE1oXt2i/5UmxdYM+tL7SQA
NpuOMQt4eqAnCH8QJnI02YGgBOz1A+lZByBPCWw6sZhGGahNyVmP4ov2kKOyUgSmDGhTbzNkvpkC
Q2pJw5zNkajaTWLmUDtDyBLLOKW1CzbY/pUFp8xC883CADH15IhymVmHYTmocs704RR9vipUKcFC
KCDmHA1PabC4NWECQAcTsnnlCfUiyg68mlwBtlSoiQ2PRuT/qQQgi/HEuMJAmtQYlTMFPT7Z+nLQ
aOp8hNAfkxqwirizr9UPDxgHcuJYZkkGd8ZoNrq4WWo3Lie0FA6n64YUNDQ7ozi2DmOw4NuVRGmq
7+KuPyDtZoJO8skxza6Fmfo2XpnOXWwjHCRsOGYIr+p/g5tNz4LyrKpn15d1+17cOA1HgWDXSuT8
2uADj3jFyKRdMV2p97Mss2IT2sxj4rB9OLNCof53sVcPPtb/lON6MBnbgR7btPiP1WpLPbF3n/s3
3ZjcuO6+cSKVjshsRX3ImBlG71Lo5wngYcXhMMLmwlGtlX9hpFuEdKA+sH82xBHgy6ybscjNmaIH
iP/U2vhS7f75QFZhVrAmFPLBs/3UWEkF0bgSm5OQpMo94cnrY/pCXraNhgwzu84kymwlNNgUavCl
KrXYec/N586OYqPpLF5DIiDg+KKnz6Sme2cMJgPt8XaxTfEfK4brAd/aNPTkXZJZrhKdQm2kHxZb
zIFes9ltrSEy36r76Un2cRJWOE+VQnU7Gdiz4EMPoydiYelSW9sA3EwD0odkNN1HvvjgnnIbehYC
JWHm1h2ojotn2nEUMD3LgeNcxF1rWP7Z3dorO6P8wdOXWJcemqa+pwr0cqhn9vQd6gBlF/M5YJ4c
xbXJWQgIIfGlznmK2TSlgv1W6I1R7oSFAcWK4KgaFOurEwWIJZ1igzty/aGMpffFOUpI30BC5VeK
TM/UiShKOIq41Zfxg98t13vcHYAtfI/5Go5cQERAh4rTdp6CL/jHcfkCuTslAlJHA4djUA0mrkYX
2CzTbREv5kbqfiwsN1UHGIa6EsI6U5WwIzr1im3GvB67lamQL+hswM5d8wMLFqFXIDY5whizYqT/
eIvfIYb1CbfyACnRxm3KSYkPtJ52XdLXDSPrgYP3von3kjYMbi7u56mnRAT0u218RW7I3fzQFOtw
QzpLOi/xqNrFpfg2l0ON17C11/LoWRnA5XeoVqQM6e94JX6PqP4HSo0A/7p8j2GUri43gH2Ri/DO
E61hruS5XUkvqVpLszlAHkcpDByx5t2UifLMXroZeJbs5POQPN34LBE4vpW6Wvvx3tvFrkGwKKT1
dYFpOcWGcbHj5wUJqyZ0reKa6S3xI9bNTXeISY/KhaLGLrwMJzcA1ZZk1JCegj1LZocVvTtAC9Ov
r5cBfhLeBuf5W1l+9nKHwJ78egls+YrEOKlnfGn+fEqBKCJBU3rDIGsIV0tAZVVIe7pFg5Ehqbpd
S77rbqgaVuqAPLjXFJ4wjI3d+QkCm+28DYoKq0BhntRtWuyUcglfo/4O3cmfAqxLcZg58DlszczL
PGgr0OAgsFddw4OX85RjHDFtsrzeYknF7CLzDITYj3oHtajQ0YV8tF52DQZMCWTiHVCBq4F1mZ7p
ow9t/mpiDHjOSgAkc1MbuncPRa0e8NFJZRDHJlgxBUwQyrxh1yOoIdTzg6eS1rFUI+ltw3Dl2JlM
tQ9T9K59mbGXmP2ZbQWG4e33m5s4u9ii6MGEx8eanq6x1iyOAiQ8hqh9E4xtuf3LnWewIraXqG/J
yyLChSLwqQzFrO0Vhrq5bJGwTLA/g3buuyjcAGvVbwHeN/j/4fivEXeB3uTCM0Il+DygYhZ7BaJH
YK6gP/T/TXm7zQ78yF+vtwpgyU52vW/dMUIm5nw26kak6TNEd2HrB7aw9G4JqCKAWXY2B1/KMaj+
LKW9DtAHVTKq29MTlFpkulXmbe0ZNIu5lNVT4nFLPXzVzJWIdY3tgMwbUjblUhVvrhkcFpGBv4NA
KlbbdX1P8cDj9IjGKaCU7fHzYChxTt7NhOyvl1+hi+x/q4fyOFDEt9bjiVtIsVFmJVc1NibWHeSk
BJ9SMZsszK+FVbus0Od3U5aD9sTKsw3SH7IdUHMmljgoeF+6SO+IG7u9P/fCkFnmQWBti5qbkQPU
eIib8sCfM38FkJecClJQb2GbmOAhwUzY+RtNt84RGX4WypprLnomSvVBTTwf5eeo/m/NS5F89ogZ
XSkTroDfmHbHASxzSeXc8IXARdtBaMJt55dyUuJ3ua0KcZPuHDt+zirNTD+2KXwtyTnVbYU6mfUH
Rp9kpjO39cIuipOyyLvf8KqvwZlXAkg+ohdb2x1+YXvolG7ZWjvzqp0g83ChLAZp1idumE0qfUtV
AjbkIp610ar4hGK4iCrO2PAce6AUtU/I4V7rQWRS/Qnmj8ZtNF27MzHYm86Cf/NIOYoR8cxJI323
bo2E7/LuZROaYixs5h3FXH18jCNY9R1UdWycJaRxG0T6KEuYjlt6WpF6BEaXnpdYcyXl/5vFr26G
RWtnl6guP0YeqaOE6rTd7f32yIc2hTTB9nc6vUEz54n5TeyqMSDT7M1ib1XYkCKGcSEgIKZOk/6p
h9A9DRoMHxXvB3qSJ1cXDsb7ITyzZkIiS5wx6jAh0/YQNg8sB+WD0HpRasrF0GFLRYApwWwWfPq1
5fHCySuasnoNC6L2XbdQX7hLd8Q0VIgPaQqXsmSAK/IbXo0Icve4vlffnjwhJV16adShUzhQat/T
smCx1P5MFLwRrovV8M24B+3/vYlhQqDmpaegn1XiXf87HHCMrjjzt4DNJoGGaDOeExpxuOQh9T9Q
y2RoLOhYHasWOTOsz2jM0n0AZPQwiavjA1ObJc5lm/QFtsthKBwnWSpWiF8jqGUZgvPcHmFHz04U
jiMxiUQHsb5P5pjukA9AMMbDqElKSaxTLbCMMGDVOkqv+y2ND3UkJ+vN8wwZxjkhIJCbmUQn2qVb
DCAA1yGUDfjtghu2HtiTR8i6OsDXePjfvhRHihC7+yHYmcEuzMoU3FTk3t9w5QEqsNvuX54REjnD
PLHVaNGUXEGRc9lb/Z0GHW5ZT3owhtXMxsQaPSbC2L2qyNkUBIlCkkkDll4zzl8s3IuwLixaqdBP
rWSkyy9gjdHioWDPq3vvMEFHiHSA9gb9hNkrHzFqHIU+POvYWXaq5sQ1KLWwyrm8VFjVRi1XwBN1
Hq2HvXvv1YFjJCBIrKGI1woWdZHbeQTq0r4dlNMKsSzo+cH+F9DOdKyW04c4XxQ0WCAqTIDrdy1n
3fTax9lUwcWSl+BCuOMvTaOgSTpgqmmesHjf7ErVzBl1+ud6UxBQVnFTHbWKGtRxG7pLDNu3j/Bk
KgrKObmZLAdkT+YvmigZGT5mZQJ9sQocrGi67BHoduHFDaqoEhUk5IS1F4ZDENH7SAN9qprUEnzJ
/WwKyfgG4Us5yYB2k56PhiOstAbOc+3SPTyIkXuqyONYt+07qFS7zF8IyVizUpAdsKQvAvT27vDn
I/++NytUNvWPWaCq93KiCrTVXOaYLfiiVaxuyeaYFyr26kDvMSj3Nngm5/D16zHMvKmFlhxa1Z4k
Nz9OFtsCkIxcliQOb9xUuXEqceYTMP7Sw8faxSt1VSjcj6N2KBdtIz75MRnmqxwdbH3l8q6ke/T9
BKsCf/4gkOA5L2rvaG0pM2IMstPw9/+D8Waht9aI/wtVA6FZ9SBi2rITVibsONJY3y+n/AiSB0Lq
IdZQvtFeGbN/+X/PXD49h01xdD8l061PLIkrJ7P0CtVEtELeelnnk+OkrnKIozfqKbxXjM6+D7sq
bVFI8wXC0M+sv/lQh9mNiQdBGfj9oOsmJ34J0b6+dSYgzPshOepLeXwNcVPX7fYQFFw0BU7nnTr/
iBO25DuLDvf2R8L3VnMGQGVy4SxBGE6CCDY3CtH6MPEDYC1/+5zcIIHHXOUTC5mvr0UCFawOZG6r
1vKFqBo1m+ZqZPMqn8amgoQmBpH5fTos3rlk4wTotKVvCjEnVXhaluA5Suv+ephhhI+d48EsTiSK
4Fhj8f04Vi4nPgpoZZxYQLvdJB5DrNYBjcY7uX0Jtxiiz+HV7t89q11Jv1U3PBgqX4/A5Fn7utTK
gF8KcJHnKh9R26iIAbdyaApqtQWmGOtkGdulaUWFkj78X5k2iDwqpOmeVEHrXwnrCLMX4NzMUQlt
CGFYJaiJg5axf+oiy8LPITdB7GaDlH/NIoQ0+b5/rDHZglcSYzQPjHkDbBRwUrQcNFYpvO4GCLig
DRBR0wRsAxHX1ty30wfG9VCQBB5buQV6cJUmD5gkWIyz/d2tOKuOvTLbkDXlHmwy8Flby20F+mnb
v5xquAGq/bGg+aZ6Shmjtt3fB8dutIqfSvFeIlCg7SGcm5U1fi2JGq0NLKUrBls9id/Dl04N22PK
UyGyZvEa1caY0b9nUdFwT+sFaYwG8yUpmr3uZHYWjtHBtDRJyncm6nG1fuj6iL2Sy1kcHyfKooQN
k2ycfZLu59jtkQ59aBrkOzGMdxrvJ6/+OPl30ERPFePyQUduMtMH0NP+3J+9DZ+csZU1siH5Y49Q
+OgcYDYz7xWjSxxmoTUcdz8H2vFNgHmjzcyPg2FU9mh89TU0TPYiLOlXBxu0SxMBLdDeur3r5cDb
moNWSeT22LbER8mRp3qyx2S0qDkhoVm0eUdFoqMSXktppBe3/VVos2N1j61KZ4Tm2ErWMOIRpId0
RhMJvWoL01I4mw9d2cQyi8yLA/fRN3YtZqHFjs0tEC8TjKqdjRfDFy+oqVKufn1oGYYhukMWYkaL
4HLCc0dlZpXOABy2MhtJLp5AYFVU8+1Va145KvBgjr97gzUT6satNIzKYfGedEOrGpTVFUnbpG4c
sfxy3AYxbgvKmemlTdO5WPB5EEmqvsov0vMXiWDXnQVXJwscwEIO5oK5U7JkjcC1TeNmGSo4WuZ3
mF6IThCk6XDAv0SHd8bA1NuTApAJrq5F8lg2AlP4rw01qK77nDJFVbqF0rS9nCP92aZv8SNUXl8g
F7xgp4gnmg+QcFlCMIBUDuNtkSlUp62zKtEpzJJScP3zGz6VZ0Feibtje69T+wZ/la40HgU8idt0
z2CsIQSqP35oG6ih3/fJEzG+8uLrO9ztidiYHseRi8kkflgUiWkkX1YP7hR/gENmkr/5gZf+mUy9
MdyiiFr4KtvCZ2TgbMhhU6KzJIGFiYHIU/shjL//20eEF0h4uew/L1cMvo1PkU1P6bauj4ZRpPFv
lol59UG22Dr7fq/nP4u8eGwFz7mseNk2ngrmDamehOxiSEQDwA6C36/YT/8t27tw9QCprr2Ujv6/
qZ2WUIyOpo9U+fI2DSkD0zZyPwmbR8t3MVBz/jqkXDeUFK5HRfw11HVJJ3enXMPWDM5LAJwfhDF+
UZH0trwyIUEHvOFsENZJe9NNEuczWskdOt8VP9JSWDaFooekgxO0EJJzoUJiqsN2LvtE6tlwsWW4
rmFYfDkh3zVS1OqRI5xUf9shHUgtkM7Y2GfFqZN2TOq0xFnszVLrP7dMnsGBnZiKfLXmpP7zdcLk
UCVn0j47iXmLLYDO9rzO8rcEjmmsVY+lBQVd2/wtzQZ5lMwlQMECfWY5YPa9nxFq3Wzgt7RP5CW2
QNIiEmHQ4KFJVQ5q31wVN7P1cJsBVgipc33Pk+CV7y7A4Ac5dfNVPU4vrol0CGJbYRNz1VQ9UOGa
lMD1WdN1QH7Q6P5aO7bA75DKm5FIHofOD/B4W/jsobX/uU+asbiOkRxWuv2SXaiWaKjaKNxH/c13
ICPNIJrtOdrD8CpTaL7y1/VXZHf1XT6m03IGopztzTVdMTgamIaYjwJVHsmxs9l0nNGXznyMwhXd
42E5vbChoohcaJledYNuu1Moc/vhHYaI0OIU4nGERk5v7iG5tOTzP1S24ybUNufISM4lbZ0Jhdkk
4/XJggmmHNvfwrIj0oifqlULeWeoXKIE0bOXaD0zV0BHw2dMl3Jd6WaalJFB7sYfmQ91x/3gQImo
LwUuo4GiG2rngapiKnP84aIRRJRoJiVogmX28GO4YBcy7wF4fW5tZRwRPYNjauOsX5S2fMUKZQ0U
5RXI6lJ1mzj5hgwm05M3u71oJVn+mq4ux/smvM/T82vwODCcbBhAq8xT0PWaRYaMvQQSVYVkFhTD
rQoS/r4TYNk/CMzveNgamCzK78Dr2Hr8wsXXRrSKKAJVlsPGG9JT577wVZMiK76PAIvj5E8honUt
aAGUdIQFERtytv6K376Nlbkg9hLDCDUKQQCVEZEAKdjybK1bNiRKuitP3hcIokEDAs5z7W7O6s5N
hZEiN6Z4D81Usgvhv+rKq1KH5yTnIw0gtVNTdV1UfzKj8HKyKJj/ppxLmMUbIMVzJwR7zxdt5wOw
Wb1dDJ/GXnumEbldzmdEHXbDqL7Yy5aZo/TU403Rzx6otNnEeSaCHgK0X6TP9uslhHC3Bs7RpOVk
QUYqFee/iMWZ7WHiIhCQNWN7bP8na21a++P19q3l80xXbW/hEFhBMM410QTR1DzYEEsJpT7AtQmH
+ZGoTvcg4IbtvgcxonpgquZWwc0rtk3HMgpFOQtjYw7B2C35ElSF67BAoPx07+26UMF/E2/7n8J2
6siwSpnaFo92psXPdIR1Mgj07ERCyjoqhPOP5L50duErDFonnDqVkdT66tKhpFw+qFj47dzM3/qD
1eRKh2PaZvawpOQpAbTkhdColDkwY00ihbwYYB1CjfO/qWBsickX2X+xN5EP5krEKE2NCd/06s9y
vWvGxu5vTk+A3Cz70cpND8q8xKOtvpldadqdMvvdknJd2ng38c/ePO61zzTiNrMTX9RdTseqUWGl
DGj7iG6ayT5XbNvsZuLNyKh1JchpXvV7esVEoRo4BrVxnj7BeZT+l6krxKWoNSBWcd6cLIZflUoS
veI8GOwSyeKVhSx7pmBPhtopDg/HLnbYMxUGatJnSP7wCuoYz7uUj+n4wIAOJNP/1+hE1VcAY0zq
t8waHD911flFuqZHUYtMiaWBJfaSPov4pw1XyXrJrmKHzA21zs4cJo18jMixRcWW+Squx5n10bwP
8eTGnyosU8WnY7ZB7JYiYoj4yVO72qG5DkC1HHcO5pbCACg0u2AAB2IuZB3cQuhPGY58t4dQzD60
JSE1cpYTTLR0kfvS53dZfxjJKCF9Hh2rl/sxd6l+SCApRLLzG6uNWT4uXBGhU2v77C7Ojqn1OfgJ
JmEsA9e9YyBkvBxGFOWrN99i6u/IJwlNJvaRx6tVGrv7id/vF9XDe6sfjC6tIJVDVmtxCym37004
NQQYwbMOpwI4mIa8CTsW7b9T0c3Fhuv7QK4/ERO5I0jILLOOzeRt9e8UY2x+HkPtLy0Z3cCJeqF2
ZPjlZFVgNUEsqYVlDh9CVK/a3xaXdO7hixQvWeCEJUmmUDLnax5CkQz/xTnOgVE4o1nAdvwQXwrt
OB58Svo48XXtO+/a3zdifz+eHG7awboHPHY3pCdepbLMWxrZhpgtIjrBb5G9o+pJ2wUcjrgr5T3z
e/LE+DNYbg1Q0Sh0CzN1/oac1/0t5aygjgLFw6cSK34KURjwdPz7fCT8TivPviX//sVcMfT/8evw
7NWdD6aJoLmD38vL8aHWXNtMJgBCBXyEnWwCoT/vxt5Rb2BlqR6evkZLYXz0S0yaRRlU1i+CwzHX
pQ7UuMq2NisugSl4TVpOKGOfMaNHGxOxF3d8Dw0HSNZ48m5r14PKRgBYVEeFx2PRIdvtorqTrp2B
TyQoV+eg6dzQDzeY6Vvsnl3WMemRlxnte2FZlWpLWC6Yx/XEG85b+bI+MdU20o5KBWdKmjqOPIre
vDgL3/UXaF3LL1n8rEmsi6lK4bpN94KP/UnMnx5HU//jozeuHao8o1vyygV24nQNVp6lxaPtWlHV
3eUIy/YedlDqua99WZPUEcqQliKaAY72caB5UHawd8Z34j9yWaZv2YnxlfE65829u3/McTFkoibt
afqfzZTNXTCtnJ0lP+QiLu+EtwsusL03lt1YEVeH95d51WYz8UsSFIQiXamnXz1FM04HkvRHjRGw
FhrxU+z5eY8gLkPBwXQW8bZRdjY/dDFSXu4AYpIv4/rA5Az2fvTmFggAlQ/BSxnyVxnlfdvpLRWZ
MFgLoRAzHgpopU25wEL0ifdsLTBSdkLt+LBBbMoxyCzAZ5AJKpFsSwXWo+qgkeEal3PD2mHnKBAQ
cxTUcjBH4gDGBkvALdWOEzKlPq3zIwhrPZExpzP3BX2YNXNfvKFq59Er02V3JLBUh9U+CG/yL4vy
jnxFH91EcKv0M/M5Vk6Et+wxkyHbBPMsLr0wapN5pyQqOIKj2z0qAqS69hG7qDirA1S7/qkw3OsA
XTvraBzxW29zT3Jwz5wa4urIfG3NdM+4HtgjTDDmz+tx4HgyjHBDVZl7IaIukwzR43WSwTEj/SM+
UNdY8pEjhyNaL175D+QF87C+rTtSPoVtUmukYOmOMUxrQH0IeWJ2H+CaeTuSK/GVbILtMVNstLiQ
1nOQko0A6FkBGFGFxkfB2q234qdgdg5W9l77mgG68IVGFJMma0Y510aM3UGoXVKGyIIqLOaJanAA
K6scdjaJkN6xa7WEk8oWUQmX/nSrKWTZr9x9GZ3BjyJuPtxP6Jr1LznIcVz8imU4jNmmu8+0JEE9
Aodfti2O7P3Yk1ELoEr9Gx/kNPzXFkQvGQBuskF3ao8tggohBT8SxhqacOIegWSWk4Ufp5GhCLHf
E0PDa6INCLWM94mCJAXVp+7yzQiZz/7oqDP+9QRhZurTkSyqqLmEMb8xpJ5vkyC6pReq/ntHIAcz
RAtaNt7PyhiNrlhRQ5LnOBv3jm27NSUg6dIDuMpp0iJF34dVnEBiE8bzI6e9W9S+gnhB9Wi28S8x
D2DI/KOKXTAPm1ke++IlJJwqx61YhK+PCRuNU11igRFgUsbk97omumaOuzBb1SvERc1lnzcFXpEU
4B0E/ah8HEagYhpIK4+M9TpUpDGeOG2Mwh26y3vShALnNNYs8IXqvLhLNnaVrSuNz3p2acXotXI4
Pzb0P1wAIVLn8+tof1Gbp+5/0mWIegrqwolP1/VH/qJtQMa3A9aaIa8xP6aoF++Jp3vC3SKVXMnF
Uang9yOZQ0W4AmqKGm76eU7h+VkKys5XzcttoE/eCg+FZ9BvHbhdYx/crJ+WJeL0Z8IBRMHIwWzt
zPi4TSxGQTRY8PA55iCqx0eaNbIZyHqBBQnMtRtkDGPdaxhX+azSbSpIAV1Yj1zfOA91uF0FqADq
zNbKjJcG4ppOfbJmdVgESZ64kT7IgmVVW8etTwBCHaWWoqdi9lXphxqudLY/dZNvWdtwyg12cwaY
g+LNcqtqe39e11yZuTfM6BqCAVwQ5GOJvQZMBt9Hk4oKH3FD3kCsBrpbx3n9v9NwP4tzga+TU5tX
+eHonhHuIaI3JjmBplAMus7Ne3VaKpIXo2g/MhtQMAZ/LWuvXJycxv3d7JwYP09fgg5auZPy6pLK
frFP2UiMxLLu7Bbh6QeH/8Q6eZMpBsJEcQrttAKVBEPuQ19ZsARn5nxRLlljWcSQaCfc6bDkFCWu
KGfZuQ9vN0xB1WOmoKM88juNuqWZNXqaEnpOqExnMcabP8lEY8M4LiNE7O2SEUes47tRWo4WnHsg
gyjpPeblhtwUDN4LN6tQA6koFgBdHgF6/UVKVs6t/+Cnz2DdQtXBm/S+HMP+lpf1MRB1Hjm+lby7
CDKPeDPOd/93a/9jRqeZjng6GUbB+ui79+QyBPvsMxdYKD9euEPMF7S4nOFI1XCuqZMd4l+3dfgo
TFsGeO3K71Lh3AX/b8kyxprdqSOmsI+vs3pBvhGg/GcW1GCEK6iRzpi1S0XgxKJ0SgFJCcXIaqmB
Xw7sR7LiPJdCPQjuAR8/enU8pt45T1aqtsCDP7i0ixAJVQqXFxt5DKXIMBZnLhKaRP6iXghEnmUn
fXAufPfmeMQqRDDGXIIOlquxH8tN5BoNWYJ032N1bLjJbD8yZtTh8Db2JWLWv+y/WoJp4LwGfC3e
2QoVBo5A9kWxDkXOKaIE3mknjnK98xl8L1DPojQSW88mev/BldBX++3h8vyMfuMVfteoCgJvKmmB
AXGtDs1J2UeqHMvXBYdcQn30rJOU7KSkXHUTaFzULzQJ+yGUOcLQ5+5sB/TWDZjvRuYzp+gIjj95
EEYq9kFWlZTI4t4ZU8FC6Qsa+Mp2Wxl2MK1zmxgPho88pZZk7u7iYFIZ2BMqZBhpkr5g9wvzEE7R
mEqy3xPr4eVlDhuidECM1dFrsfKvjGqjWrDQkVsbf4ZPa0dRaNVE09iPIuJ272LRSimWRTEhm6An
A1RLeAlxSTErvw+UoEJrga6lI0GkTxGKVKDFAGHHYzZOL5VdOQQKDOQyRhqIeRopaNANYEKX2K1w
+Dcfk7SPoUEWUkSfZkxeobFrZxROnpwbJFWdtssXxw+/c2YTvRuBqqjLX0FChCAm+5AsgGLBzdT8
X4c7r9eMtHJ7oW9xPmeton9koyzxXYo2G6yNK89dHZBWNIkVfB19ygMANfSmEDV2Is8fiL7mH8rD
NWEwMq2KGi7bAN/pkvXHSEklp4g9ufuDkp0GV1ayLtdQSGs+pdmDPSG4bCYeWRadnYollpBpEDQ7
ZR0Z5cUEW3p9UDvg950TFTHCSAg2eaVMCjZ/7sRjgiy3AQ8PNJfw/spinLHDmysmQoIRcbJHw3VI
f33hQWy+0JvlTXesLK0zSFEfnX+rPTMMsAliUmT573rDuKEM21JiYVuoj1mEHARhiFkTtIITXYaf
9jCUojdTlX5m3mb7VnjEec+j+SorG7YmqQoqCQH4SJKjnoQkjgRDq+2tXDXjQzMzo8mUPdCn9NxG
/BvQkNQkZxqyGLVTvlkHDvkKVoW35H6ke4duWNzBjty+bd7wXBbD5h0b+20qXqtjw/l6XSVl4GOm
y2fNfjTokc4DgRq+SNRyxeqSMIVDAYxaQopKkSYrGTDoH1vS72nO0WNajBhb382bFlNp3HB1XymL
XiJoq93GP9yo5tnAsvCw0mNlvGOLCWf9yrlOpvM2UMYp1YdFdzTfwJK/T8Pojlt+i5bjP7+/GHE8
NZmzmvXtsQYQe0vc5b5XTj7gFvrtf2r21ZbJ4k5CpaDHCLzCPnbY2Nuv2cCgq4atIBlQ1NslvAGN
9QpMvEVSkUOjGKZpe1v7lPzG6LFFIplcch1jsIt5lqROvc/7A092pyF9EeeYIX+mVq6D2q5KLnJR
rZobxJ1adnrZHHiO89hhZCvnbuMN/CGaWfyfAgX+dw2/+vvUj/9ono9MTNFZpEWIVHhBY6qVcwnY
JC7XE7LLmqPVLS8Xgc2aV6P7z1IUuJ1/P+7M1x1Hze8/vIgkz2eJpER0b7GDxyfZA8K1b9LfCRB3
I9mfLCVOFJEbMApjiyEGWs1o1NI4jw2tZeOdTF2eMrAB0HrbpQqsyTqMiKaxb5oHFvkpDfssa+Je
K7NWabhBNGyWvC+rk4GHfHoz+RPbmEm03Zntq+PWLx2COClyrBA+fuB9XioF4JZGd+BZSfU0RsHw
b1bEnZMVvNblcT9lDUjR2kp7BKwOJiEejbOGyLY+yEl8IFncE698v0TAFKBz9LrAY8mrA4Ir06Fo
powWfxrzRAKrBAfPTxYkGy7qYpSnLtAAZGjvFPzAPRH9FjOa0c5uiJNnSQFZzGMJNOehNQUVXAEi
ESPYVFfiilxYJFi+mQObhy+sNNX13f0IX9vCG8/0pEPNMiwC2WZtzJOj8Kf3mUXRkC3eCNN7SBmN
P8xoa8CFIakTl15Oeyp7Q1o1mmimI35Vnoq9dQlnc8IPA5wIiSL0Ere+tCWcwEEyWBq5nHNtR8xn
yGFQOeVCWNt4UmPO3hYq+umRGGIMd1A9bugsGvU/foeUK3uo63jpcM4NJOXLtEpI16mBbH2SecVF
y15jo4eatu0E1siEWZeEpxQ4fhRe5Pacf72govouwYtgdBeUWdhJbvLv0nwCT5RxBevBRLNsYpju
dV1Z7xK41aqUKXcGhpzr2twQI6+mrU9MpmQt53xmJHjibmqPB/dqixCHK8tfd16Lq/Xh51Ddg13Y
4eNrtCtHQFzWhsy3IlSY3R0x6mvEQSK+Rfz7rf8CViK/9WBYeNfw7bwTb9W8yCoYGAXKZ0J6wHY4
/mxue34T2AD6fdWQo/QhziiyUD0hOFU/Za4L0tbrK+hlcWmKAvNHQwHZpYsqKpqDByCAE1K8kqAL
OaUMPR0SUxuiGrXWDRhqtDJEA01M0LzveNaPNMX00aDYx3E1sXbOj1LNEnGmjwdbdaPKmb2GBmYg
LM31mEWvkqHdLaYSVz+HIFN3Y/FZFeU27e9z7Dz/3aM3MSmlorhE6NoGwhLw6k+rUMD5jh2oGllj
bJRWwsMDK9gNkWG+ea/i3C0JbaOYo60JXrlTVWVrOGdt5N/FHizCFFXZmJj53+DOooXQHWsJjpvn
rVe8A51HXDuXPl/65Q5mgVPQmcoGI73njDWijv2NQxT/uI74gD4CcBOXNsEd5fWMWXT4JcZQtVbb
4EG4mMhvqTfDudVvQqkZE/xEmXj33z20HX0RfLAMu0yeJXlWHA28FThK8PnehVn5etkr5rrczKAU
9/BL69d+lhoQvdHGGc1wVs4GgGERJVz5ZgTyZf4QNiqZ6ABmVtl6JOITaaMzHXco35xe9h1Bh5Cw
bUS1hq8DEXJl4bmQ7gkWIrLgOdFLb9+D5NFZhHDQQKVAGDCVNa12Nm9is0jcgpiJ/thfodYZw8r9
SYufoJLq/lcUKaqSG3gyNH1H4/xbFni7KMkAA/1n9QnKekhPfw2mnTOAsSb1x3VsefBjzKuN4yX8
zl0PwO/YYrFxrZSt/pEv4EqtbiBBo446KlyGMM42aZcYn+zOAJ03ZLwRdgRL9x8H0HNBqjm00cuH
iV9GPuO9oJ7CEGKeAUHjJioO3y+AzYAfQnTsKdUMxRB4yjaYeb5hF50IJO5sDKjLd9VhA29FgjR0
eNK7+zCbyfigPV2oetERPHOyeT4QfS1E3QRlhZ4IhtmLLj09+zJzDxTZlCiygcZ6Kc/1nOLflqjC
ksizR7ZXp9iQwMzIls5l8cnYPi2w3qytJEYJXPHNWSXeR+IzlidrxMPCtulreydN2udbBjbyFm2M
BUABreZBHb+XidEU8B34cBlLrKImBqnm1aSy5ZWoKRHyx6qCy+Zq5yaYRkSAhC3PFrfm9p7/zeyM
/uDwc2023u/zmkb5LFWVIhHnIj5hYp70UyjCAo68baAzZy+Vo43p/CFAAy2TspWImtHglBrKySbp
S/9zWwya4o/P/BZAnyhSi2ZZnltJg6A/kM8q1+1s/ke1KLpBIHc5IRypL7JuY96e6eFiwoGo7bMf
HD3+a9KgbrSPvOGDlIYOKLH1ops7ABao5TUvtjSjc64esLe9LUMHrbdbQFUwxRaICQu8MAGMsdnW
pa2vrKRI90rCKvTckzhFYspdMNp7rjLBBrhYbWbIwWvRGcAtQ3vA04siCQoiv+SkjffP6PhqYuiv
BIzo95x6Ny8wVgIK9bZf/TZp4hViP+ImijxWMK4W+aZF4/IRv3PmBrzOIeiY9KCJ6xMZPZG2lEtI
+AQvgmuZ+Vfeu2V1wKnabngSmSkiJiWtUp6R+DZlLRwJmOE24ufbIuIVEYtOCsRs/yTDYKfv00Ui
cXhyQBJfS09AQ03VHzVMpkbDFFWYiEWzdoSt0hsY1fVbYdqLJS/m0ovrSXXOkyaboMMRGjADepIW
CPQZV8MI57sL0Plc2j81ZSf17vejqUnUzkwmJc71WPkumu24tIYpWA4gPSSnuqV7NpClGZUozy/5
Wv6WGmBQO/XJvTfICprkrOyfRzDwdhP/EMD/MaxHSGBUvSjYvpHm8JUn1ZUCymECRTW1K3DjMERV
Q1UeSCIalH/Z7SV5Rg18PaV91pMzJneZjPA6ntsW8jtnRAWH0yWmzveziHndCF3cEBqCJZhYT7d+
S1U+wO9K45SwNgeleLP1hhgEn+oL/S4En9v/8EQui6A6uy8DC7pBHXIaaTrJQtTj7GrFZyHguQ1j
vgPDCeldnJ1wJSIMhgGRo7RmA/zKLhpXxNw4k14k5TaROtnD2BoqiONUCA7lfKk9/TiGbHnZHKJi
rYu/CDAxIXyla5UJQRKCHlhwtMtWMCH4xArvDSCPcEaVs1sQJHt4Pi+0i3z+spunjLn43y21fwSe
m5YzndwlNZNRxCKKxkqxGu/jNSBDKfkKaySsCbfi4nfNEYx6AwGuWMpqVH1e6blSMaoCSgxN4Y1c
/kVwqbyVaGP+PtBjsUdDh/42QVRFeumULKYaIUnKVFIJS9+78kJlDIZ1iRXsJBzXZfU7WNTsCi0b
r4LVgkGLV7tqUEy5CvrQSARw00AzaaYPy/1Nj7vsNBz8v4+85SZvYFjBtz0f/1xy3OqhVznR/Jfr
Ol84SME/zlhv9P2Y64Z0C7vn1/5ymHz24blRpfOcnMCCTQjfeFQGDrgvZUSjhdb+Pmc/65sZFMPH
pgy/XOfaNxqLQw7xugyrviNuWAMEy08IdhwLoZIA1EbEotFOFKYgNaV4w5PgWNzmQS/IiTcU2pES
uB9fuPMzy+DR/Hy3nj0YnSbx2XOkC/e27gBARvqYlgu8y0dFZ1SSZzaoijSpMoHwtCsXWYh3C5NQ
BmdeNLfEqz07yWMspnDrYLwruwb2huJH4HX+6/5KAdfSNYmeS31/FJkI/fe1d7q+oUGhRrWYVRC1
mmDrwDyclGdeek07px8W+qikgnhVVqRfxV7mo1Q/igWOGUCvjbKCt1LsWRtm8khdxzJ50QLuaYTn
enKA1pAmmjJpavSBxoXz02Jx9LsZBRmw+Fi2MALvkfKt3HaNsOTbk1wYMYiNPOp5nJeD6HqWdgXd
kYBK3PaCbcqs4G56tT4IzKgoP73qBRXtQ61tCMXDQqQ1Lzi0CFA8nodLiVbG76EWO14Ex4lAFg/u
VQqHrgsAc/h9b665742JykYbPjQ5Y36xy8ASRwLmZL5jJ0pqfE2OnEcOiM/NiOQ5UsAIPleJaKqw
tye2Nts+4Ju70uUryZ2T7x7nmmtgHSDUVRkVxTo66JlLU/L5NN7Qg15+uIMQZCa8v/bIPMhl0VaM
mehMJ6VGG/qgXfzOK281gJVLEiGpGQB9xmSsfuZykeQJs5xVqkBMtnQpiw2nsotAx0+Uuws1JaUg
QUkElpJ2NkjIudizwPKTha75Lij7HJDoyKNV9k+Li2R6wVHv0YbzGbhobEc+AyjusMtvYOLDzhBf
7PfFgU9KVONeWsL1sP488iQRv+5mMSl6y9Dg0p8WIxu2TH0/qJ8W//f7HQXYpCbecDKFIwOZkK9L
crGohqWhicbZl2YL6Ta2MZwMVg42dC1mexf9DwDwY6JvdUJRBxPmmJ8YBtSHrs1BY2KpB8/gs+59
8eXxMKJ7GUvE24WSIk6JsLzBHRC5m37lkvR0AbnlHX9zjAJkRA5xexFnpf96dhFwvhZd41QHqJga
hZLClQ8lL6nQkl6zoAOIATFPnAti5sDtKZNdCQC36ErqKoh766dsKaFrQPe3td3se6gHlaaIeZiK
0gEnMZb7aYznHYsMPjrs/RyKhV8ZRzVyC/QLNYgLhEShUJKI1tjKJW+/4xcAHQzKVIDMme37mD83
h/egRjekzp91lCmcdTFttHmyrRPuvNopOmEhFIoaTgWMtGGvqH5i/SMXvjhDLMdS/TZYcQHIebuN
mFWiaX2L16+37tZSnLid7YDFrmLGeCwg/xJaJK9+mENA4389iu6pn5l2G9Fm6gN4Y+OhQcFGmdBv
amxl3zNOP7iayzVvSsrTzSWhfijz4GjgEKMIFzSmhkW67u212h/G9eIGrdAQeqJ4GzWlLJ0WjPE7
OJSkPws7WEy5mvbmECxQcVKNLgoi3KJY14zGp0Sz9xGO5Wr/n0rxgrpVPWTSJiqfc/CNCsDh/IZO
WzPc1PeCiJ8YC5/k77TWbW9RJMslp2SEBHELjJAAZQ7DyEbG9t6isPpEmv2uTYi6IUpp8aFfI+gI
XzdN4MSE0+a/8nTqmYHuaLbyZZzb3rrDMR7dBWPjEsk9Kbyhuo+Gv9j102/fOlYj9TJziApc6P5m
jG1CJwNkD0Wzh8UkPRB9sltoAOsAu9eR+qXpR18mO/asIYzVr97TM8L4ODVal12m6kTnaEvAIGcY
hW10sHx7yxjibujZ4jQGcph8CXVnxYYAhqg55U+X+Y90//qCNWlH8K9wZ9Ku2R6OpLwgEMN42aW8
GpYpdU5y58kkucIiU7+fEv2g/8jhZ9DSWIVAqDXchDwT0MOvjw+YfR6t4jB7ePK8iergwOPLKOcZ
mTPcIixochdKDu2xt44A4GQs0eDTh/yzmm6KUqRqiBWERMo0kmm1QNw7iKwZ7opO8zfrUrgBlbHC
ihLde5vvYhjQePyiJpTfDBRYAYi5ZfwM0yOlKU/BECs/Abgmb8hfPH/jSyiqB1a3o53jyewTna1p
DAfAaMlkUjn7BH2AC4b/EI5WxzzpkErHkbaakSkMvGVQDOnqkgjCgdc3SCl2MFswmzAG/eNIzgu3
0nCsk5b3fFPMv/9NJnt+5juSPcaq9X1/JuXpwSLma3Qj07xgSC4LoinDMMrCOD2bioUp5engOK+X
NxquZph5sYOLNYkPM4B6w7Q7uBueYbCGIF5yZvusB+9aN3NEF6YwiWrj++rfaLK+m2cGKEHaU/xI
8BJefSnfcbDWSGFuknoIENi53GLExbWV+NGzfoacLvmpnu9I4N2+OtCStyYaDstO4BPoAQB/rz96
A1pBQY5SDVX/1qUiadgjpNpbmgEKFECnaoq0H18x6s45R2MYfCCODKCkYPqeABhj12xv3Yu62TUk
oqqsOsVpEbyF9nAYa5JMqMrUPpPPvVXZUw2uijMCIQbAilJyP0WgBmG01GwXior5Vaiq7bs5nIl4
JEnZ2Ag/Hp/jHcPtcT1PkpgQ/BEq6E0qotaLkIsdOaqHVs40gPEOA6KfkOmii3KeKYvWcugJvV2Y
riDiyDEyhUoq8tBCEMqgkZXJhcVz/p/k9a7ZGGT75MpxRqbxkgtMHHb3fLKAf/PX2RmM8+baqp2+
pQkyu7v8Wk00SwxxRd1nYE2tHFQYyqzYj9t7QTED+I+e5b4hmbe5ompHdMGW8dNHMG97MKV/+luY
4KtAo8o7/8nMB/FRODwZwSVvpPCPeD7jIpEcjrEpPKhEl+6bIkq27YZqORarune9kvtWevzHfhoe
kg16w522DkzKfkXO6ZgQLuBcTVQXyqyYfKLffYEjdnOKTqEBssf3wTRwhaXrklgyLA2kbxC+YXZ8
phFSTkkTj77wIWdcRkVudwCmdxMuRJPUvDAftmQbqawQD99q24eqpQOnDjKZnYMx1AxOC0gv56H0
8paqgCLw72nPqYjFP7ZRwkrxfa348JsLIol+DabcvFMzjSe76zsdfXXw8uQHTwM02Y/1ffwnybbb
f9etbcdcZoSrjxIZni0emSCAxmzOuOGDeWBtRzlMEBDzM9ntVx6vZBJd2UU4s1jPzqehAhsi4Hr+
uSWD7MjRxlHrfKVUHqfESeDGkQtIxWsEdym+l+42sReJl8ufrA0mGEtwthk6UHhubQgwFPfonPP1
WEzt+bqpnPE6s9rgDk9l6ElGaHd1FJg5QxRGdcj+jMocz5MdmiR0FFZQHCLzXoqB/kF+LN1UGNSV
d67QLkhKFmAr9gVLMvUxSHd0jIDQIumdTAIz8VStDdIcCFM5mASbpNLAztZ32wLSRp0DTI7nrgKe
76E0vOxbcHbZBWvvTvvZeH06qEwvO4o7aw9GCY0Qc1dIgZltuK7PH8pDWyjUCnbFLmDjny+FQvp3
HcAN0S3mrZVKfPGj5SeS18xcaahvh+7fDjCdShQhCJnjbJ5CzkLvsmU1deObUnnAgpgTZ14NFVJq
yyT/m/RXfzCPRlr5XDxgLPBNDHv2LWoUxULV47LEHt6dM/JKgGl3mWA7rJJ7QMYvVnRgvb0F6+vO
XL5NWP+/Iv4903fUfDSuBifqKA+zwOJmKM2RVHhaYaxfjeydQxcoyqe2Jeg63BnRYPESB/D6046A
CC7xD0u53HY44RDvsFJX830CMBwsxIrjeiOwVe1UkaFRWYVwafM3UwfJIuHxCSaaIFzHwUMUASY3
P1SSwIURtxVCEc7MITYJ+tBPFcfl+JAYN9oEV8m32N3cy0xeFuB/Brw4rmyqeSIWN3FcNpOU7+Iy
ddAKS15fJ6pr637t1dL4gIB+CAr1xWGD+7oAhzvjzMEI3ivSW7Q35xxh2mZmTEXQoO2G6EbbJ6ym
GQHcaxq7POqtiGzDQjpn7W7fFKYtHcOmSWmA01Ky6O+iA09kjiMGjL79kWBW6D8tXmAY/kDJgaPT
7zXugbZz74RcbyZr9f0lvJJ1+6NSp4eucC8QiEAjtWufW5rfKGfCGYBc09g7HMssmfpz7bcJi/jg
MqOY0ZMmbf6C5ggWdeZoWeDRhzgjZijHxp1IgpWc4iw8aBlxW2R5FJzRwNtbGB0TaeOkU5T9XXA1
DPLsDpxGGBD7rzr796Hn0RbvlctW1lKXbuJHCytN7gsAM9z/qDWoUi9G+H7xW2ZeIFNWghygn5wP
Zbn1tKazP0pNnPI2LU2p7Slucd4A0B2I+ivPcQT/LXsnnu9gQeyImzqCp36lOthj08ohw3Wb54cw
ZcQru28fZTbeCF8bEU+hL9sj+uAt38+8lIR+ipCoQWZGJnMZ3rhcDHWy9mhfgXrJWzNJsSVp5zgw
B6wriu5gCukaDk3DU0vdscTsvjpv++E+zHpNmDxusl5uJZJPlknOvMG9tKX7yOXD5zFq4JQlxU5+
geq6cb3NOJ7cIC9c5K5tZsl6OL00NKU+enMAmOOxj1iAjIQTYSpa0tHHygUuMA0M5IPPeOh/Gw8J
FNaPUcID8KHAqxz05w+zE+E1/pX9VPnMg6G6t24OL/j6sltNMvNGYfQrCYpXXmDtztzOJN2WAnkw
Gi63c2XMuoP+vcgK89Ix2oXEazi9HBOjdYwUeeOb+apORrfbs2viQqZpCXaM7FcwcQzGlBMpaNBX
h11DtAegRaJgUkZnUWCdSA8kLjt4iTshevzIxCbg0fxmXn2+QI1PFP352Jvvp2XVdkRSmmXp6ZPV
5Ld25Kk3RCSer9hFViAPDBAO73tQ9s9LC8aSykGHXoPN4iOUsXjQSAqhTRDn6/v6WUay1i3eCsvt
vPuLkL6586gV/BQAMf7wYDywo3Yq8VqyWYkJfp+w4TT6li8li2ssp0dqGvOU7bmkhzrrnsH/rQXG
sCK6HDpGnoXJ4ihsxXRJDqJGWDU7W02+u7cuP41pBntVXuu/R4OO2Gk4UpmS/oVfFjpZcRU4xwOJ
quYeu1rfH+Rg2NXIyTIEQArcEQl8STa2pdfa0YD+TCMYbsWKVFvIpPDqLw290SSdNWHkyLuenXrr
0zqyjKkK8LO7oZaFWAhyf9CeMM3X6ubtoZqauCo44YsKT8kQd/zlOM69UqJ3/CqscbPxcUnzJNl1
/bNvPEdRbf+w8huqv71WnZjpmHBc/55mIM+lhJAB6P4q5/cIJGlb/gdfYKHa8CgKsbdNVnoG55Zk
NN8WdmBuiPUXuhKeSVS4TR/mSq9lR1ScfATAlSiElS5k+uZmmCx/InZrwYDykJI22L4d4Bx13gWQ
2zTTnEIVMuAfkcsWRwOPkJ1+UOkJgOHOG/E8Xvyfs2RPFnHDf1lfwK0thKp9WC2wRVC9GVRffCIM
aBuhtURXJ6oWkMeg9vurSWsp7fHTG+/85L0ehJjkLf21XqtCnRvsVky/NU9RalQpiGIboi8p9HwC
+CqMkbL0BtooXibkP22BQBZXTidOaVvB4Q1hKJrd3pnissFvrW6sDxJTsufuL2ju881R4xGhsV49
6kTGcMJG3LGFLS+NcTU3q6kxhiN5yjM7xtRWWD7evCjyNnpJ5uBYUTRBNmZhIpRZfE/mGaqTu1mS
oRQ9uNkNPNrwbncgG0ToCDcY+XJwGYlO4K2UM2WUcdxSoqkALhgNHQRB2N3PEDR8bFPrDyWy1KgX
1n41fQ4DBOy8AQx/TY969HhjrBSI8kLigmPQXO6AEH4hVqWPIANWOIRFTFGFlpLCaaQmC+Or/caJ
ghIRkLv3XX3hryGmXMIjZAuQ/J/vUwq4Lh+8BHplYffuJD34HU/3a3BT44HiIg6hI+KSxMb6UhZG
gBRN6xI9S5zJv4VcLdX5+3bJHkeJIYC3HGuGrJ5nO6LIHLwXp0TUA4EeMG3qZcCfwJZIONgtsdNY
I6u3UUyTpZbkh/9t/XyZI97LISF3LVfWd66L1vcyr8LNu88nT1001xEeIpwrm7SEDSL5bnbeSOcW
KE4yrp95lQi6xpA7OioUKDBXuXt0nVKsrZqVRJoeVBrXaSMrxUTfIekdbJWIIehq09Y/nV5+eMWw
S1yriG71LcvRPnYtuqDwgG0h4Ylb3Y+xvfX8aWcPBP+8yhL0Nhi0VFBFzLCn+K8WTlzTk394RueM
17Svf2hP4ZVNLB7PgEUdugky906FWMcO69fYsG7se64SwlH+HjZGz222i7GySsOylOc996UJvJSZ
pXcFYI+JSHphSTVeVxvng21echC9EypKynTQwdKpucE9IVhnyMFdEy7MXgd1hl+VbMyp4KlcMr2q
ZZmamNLca2T5BVtGeN8Kc76sn0tUh48tFJjK436bWN07uy0SmAH1ldQiSbbxWHY2j6gisOxjCO9u
S7tXDTwcIlhL3uW1LrtEk/EZHGLAmEaZ5hx4lCOTZe4iupAk4rGEbV7FiBsG+GY5ipHl8A6EpG0w
woh//zifyT0d241pdgBWhqckWhtfELdytAGkV7PTrSAWGSNe8SSDT0fF7xGIzfFj1dpLlmTwov1e
q0TJVUMC6AgRywXpFi36FLoIsOTpq1lBAa7QJZcsZWVxJPbCUmESq0J1OcQ+ePd6UrV0ZctfZ9Ef
XdzhP8tqbaQSez0iWEUJyz9LwZn2UmMARHLkBgPorL05iPLlOGmPQGWqIRo8CgeTVsOv8s2Qs2fK
7tUQ9vQlsINT8JR9ySLaHFvmSH+beqdy3rwmYfSdVJDksGI3gZSsWKpAE9P0iGftujzYNHAU/EFd
9PZSxT+wm3UgZID2wi+92vS8Qp0bxJ9hduyyhKuCbyhuRou8k62+peMdWY+pjuiQTW9CkF9REp0b
wZamAFfN/atg8+v/rlrZj54YpfWV84SklRQjbPozXhc5WS9YscLwln4zsVi6E9ZLStjxdYUywbML
o2bVDNvh1gOyRPIIctFIZP8EZt7wkZ5uk+0/RRzq0jghRl7ybySufZppGxgdSetlg8zzdfWIM+vF
UpPxF17aEuizqgViuz9ZZtYrTWKhV4c+RO32tyxxbUjOZSzrAD7TpuAj84PK/SKoJqrOsm4cF77F
wiU8KaHXVVDqpVY8zK2dpPfjOTUWn0c+8+cG1KmPU9j9GYHy2kCNBvCtfxuJR68ZOy4jUetXl3LZ
KmKkSP8nOT4Q9+Y8WT7BqeRoMuHyWcOJKAbbXS4qSohpKhyjSMlps8xkW39y0VjN3yXZobo6Jvsg
Jhbk+IW7o5zYXw5lxwAM0jFm1VANzN/J5iEiqQJDf3Hf9xopabkzZZEpwWHrW9ngRGG5lEjzOJPn
TDakc7ao7fxthX+Da3HR2KuzeZOaMvsSAydEozuRrJxjcQtehVuHfrA+9D0dQf3LYycJJtg77BzI
JW8GEs1eiLx/8+/HS3hCz4YMta60V7BC0TQu6G5r60xKj3ys1wrgnbwF9/96V5OL5htl4C/sJc78
4SBD9a9zmyTgCqAIlSC+2yDx876rnImfs4TzwNLPHNDVBmKvssMRI/8yhQ74C9dmByM7mSx4217N
P1bZGFyrXXo4eB5wG+eiQJj9bVbtYthdOel9JwaTyBK+zC0hyBDdh0biib0GP4oy5Lvi6gIXxYdL
i2b4V4lgWcdyvgEFhlB1TLibumrzzESSjzU9L7Pn+0+LkGNJhYkJFK7P15znZl/be8Mzl1tu1ElS
0zto8uUf6kC3g99huhT6IaLusViu1KHCT8hBJBEoDB2rq2jBL+NkdC4wASP2XhFdcwnbYljgDYid
Wrd5x61DYokGcFaXbpiSPhZcXUxu5ythuMCEm9xtciIkbhbN4JSQWQgY/f2fmDS5VVC1dvOiuMzk
wZS8EqUi9vIhmUU8+vzE5f/MuQBdjBkB7LX1t8U5eWSwhL3+y0MmgD+Iq72LyCHo2KqJ1hvU1562
YKgn91UuxhBp6+owwhP4lCKZYDhRxNKcvBcvQGuCx+rwpwS4SHM881UR893hvyTz5WvYlWwoKJi/
cIQS/cXI5xFjE9r1A1DAriCtm4uvO9HZ0/xt11STRzx48bRTOF9hFh27KQQKunxYT0tFD5uBhNxB
HGfnk71HRfj7Q6TnXvgS838S6QMTEd0GqqVt+qjeNJ2MD5wZ49Wa9TcHXq02X6ZucxabQT4f9mEl
/RbKcdhFbvZT4dNj0lEoAh8B7Wpe+/1WarHuA0DTrLZckUJx0VerRpu8S7DviiEUEEwXF/44s5Hu
ERkbYg3+Dcw4VwRkE02KtXHthfIL86HDcmH4a/0QMF0CYdbtUpCO4Az+qXCTZ8qghXhGtS75X6/Z
Y8QtetCp51wFmSDYnlvqG9IZZlvxvSm4s0td2JKBx2cUGLwks7YPDqNROXvIt9F3HzYRoVxIrvuO
5adAcw/DM8pYGYhdHSKfTz7qmmb6yGvREMSEexbqR0E2esnGfr/T6EpYlnqoirUahvsEFHMj/S+P
tAKGzjrAT+8aLqh8dwdlwJVE7q0rA9YPs0fc4nkKn7xfg8y3Yut/srFSqosk8fi55NvFfNE78hfw
vDiGphng1L0N3r1t9mswlQndebOTfqcZ05IU1/vLI/xsDuxrfce0i7fiDowZFn72X27dKP42vivB
jqZEIL25UFI+bTTlSRn86nEp0awwuXdMPBDAFLagvKLdMjdMTTeKRj7wLaX9qNbWhJm0vv7z7Jgp
pw+5JNFituVqhY+7Bz1UllkiCi/B/J6BZM6Coik1p1+zVhMHeewSuX8+ZxezQwLEsl+MjR3tH9QT
gLbQj23d2/gfLfhMC1dAKJAIwckiN9vVYD5sLduC5qGUMDp+tRLKEcZ0iM7U3beTlnuqS/TdmV4X
jcCsCWfNCGhZfnly7xsHTipf2d+jnSzdbvqH4XahOuq4Y8zoA1B7qEEhR1BNHJD2Zw860/9qCI8t
Etvpf/5xpztnz8nh9Q+V+vyUzlKSz38ql7QiVZ+dY5hyA0KX0oHiuItooIzG9UMIQsrTK0ujawx5
8SJ9qawD25kiuy29H+zkUg+Hw07Jb021Bxk8gjKhDHm0oq7DfjA2fJRG7exsGv6KaF7TzNG4LhaH
sHN6DkB16tltd48b+P5D9GfztPLx8MXWcbEy9HaQ02hwtTP+N0Ec0BfbZsgPpbTpqtUfhlj6IuWj
zPdlIkTSYKEQ9S5PH/hwREJnsgiajHiA8vVmRfmoUftiapIuZ3oy/0UMIIRlh1vatOY63ooUAiHH
ZtF7ClAEyq6Ey7gOzAfam/n419GcTibxFOPCHBfTaKpZ29ilQWaEEVQMV1KuKScr3xRC7rTQueB3
ljInffLtbI0oSBNwS+A0c+WdsOmBr3kBKkfthUcQ86/hPwqT6auSMtNxiJ8evD8M3ql9RRLV7xeX
svNpOwyLifsfZEi/ZlnA0+uM3T5Rtbqjs5BwPzokg6+B3ePbKn0vGWvI2+5dTWp9qGV3g8s6WRBc
MpYgXGebPxz/hXt7XTwwewsklzbnBahxHSFHqHw7KBFROenPCiPGK7TPZd55z3/9ThzCnUL2F835
Hq1qwhbAd6MLm7FA/i/EXBJqZ36bLsN0LA4QD7143t56Y+xBAMTiwpQL1RVfCvmODzIc+hhcz1Zw
W0WeAPBU46xi+0/NvU+c/NnQ40gSErSU4n/4HncjOYb7BLU9KXPIi/+9e69g91Mhnj4Z6MSRqOB0
cjAdZ2vYY8lWH4ATO3L2OdKNYxG/37kkF/jWXFulE+OKlfA15iIiSWrM/IinRYnlDqagWQIcTRd9
8611nan2TRHlD+D0zVCcfuDimm0L4o/cAcRVpAkAZy1UziYupYErBaZt2ZNsfP4PJc66balGuNvg
87yerMYgPv323BxXb1g2tW2Z8RDgoxU92Frj4MqNhCxX6XeGrEjMOdN1i1m0wmAyNUoYvDYWEFvb
sDRp6R7O11MxRG6yT7eKL/vj/PS0kfq07aSFKKLcf7EMGmKFZpyCQFxrW4KOblPSZ48P1Fu1w/BE
yRmKaD6gsTzffYhT7vfzjy9TWJgkP7ChDErhBQyd1fCWGaFJBLP/9Ze8yiHjcjTpcJxoOJvUFUTI
6pnbXd49P/IuMdk3RoSNNEKoS8xIzJcn62+vI627FmKjU6dYSKreFD3xfZyaXmKHfF2umwNRtzJj
/GSY9wk3Y5a1N8P/jNecvmroHuX+D9QrXX4gKELfMlueMPtl1AkfKh/gcgYHa/brUGRQ2BZvq9Cd
hZUi2hZBK+ei1pmazfCdD5qEJRGlmEWduc0yAWr9baRlKS4d+TfUAGQmVZxTMbeWnbvEiDgmDIja
rmwDALqBZNUT9e4Z935yXC/fsbLFibVTVJV1cnnfnrxm6358KocN45ZMuCJ0rNBCNK3279DwWmxj
imcQnfP+E03AbPgXooo8JDDx0AgFa70Sb9HGe2tpAtxRDWwY92nbpJic6XZR4IHJln0Svzyv0wWH
CiZwdMGinq/JKeO+/NxJXV13gzaHt13Ly+MoytmJWeHH3ChMWOGPlWFyzIXw5TTU63DFZ8ZEaSp6
3T9SZxEdAzWr3mYpVxtQdGjRfBYRYHLgyIpsttAg4KMqaMEtQ2rVgMIKDzbKv3mWDCY9w4Wpbhr2
+DIHgHrMXNQRYlb0cq4yUIprYr/+hSYTzvkNSDuG8xUCZ/u1F1LsuHEHjfuE59MYcK25FXTLGQj3
/Ca4lqeSF9q9FMjoJM7JZ0OpJa02s+mK7VWU/G2/3fJZO1Z8AVnVWsCcXA72WfOcx3/Pi3bCGB+W
AJAvlz5e7XfK1YgKM0eZmjeEVbmm277JaQWAM16z/tF1HICTeISHJSv3F84KRTH5IWmphvFhrQLi
hNoSL7FgcV9dMtnrGRJHd9tOsAFuIJVCkKtLtGv43SgiIEfPQLCJRAWlzifuxHwtJpAXeSBOxuFi
vpak9mnCe30LwmHhfnZOZWlJUB3QxzaItdpDaLe2eLTFf9NfobtPbMU6djEpXrlJzK/3fKIdUCl0
cb69ksAdCCF6jtnCgGzZ+v/piBMzJ5bV7QwHmYYrzY0wr3YzRzb3GJba2q9mLLRoaJUA4QovlHeq
BZyFaY3B289cNY4Xk/zGc6aj+0JshqkdV5botRP2DgBhe4mMpiwRpHGv6Ch0VR6mI37IHkkTeihf
wFDnWGZT2xoRFwidaK1Rf5G1FEwWvyR+XymqhjEReE4gGhA3PJRDE9kzQbuvDtyHZX/m5xSbTGrS
E2shZ6hQN8/TZWUy9Z5SDCLSOnG70R3I4iNJDu0XCKVjUtUoOhs/9wsU4fQUxrzorzZscLUES5wZ
C1Hx0xkDe8TsqPvUTlR0RHYoa0mhqxhOxaGKHnliw7Ild+VubrEoaSXiSofD4H0J4bZBSOi8qRv2
iBHQoUs+Et9cayR12eW7rB35BTEt+AwcF/oSVfwu1M9+uZdfj/xKbiSEjlc0fTXX1Qj8cGIzBKi6
ic7wiZIanASBhL3dsLzcGqQ6xeri9f8vniAndoiMfz4/QstKsX4Ieirdm4K5TxUxzEjKsp+2XKgH
ghkYd1kNR+8uNmns77zmKJuAnQEtL1YFLxGxHlgwqIpD7yck3VA5Q4YfMCjcxsghnl/3OCJKnj2D
tNiJWvBX5MpFj70XS5PeXXkcq2YvOFF1nRrAYlr+E1mJvtLr2LdvPtn+Ns/UR8D180+ipwyLQERF
n1SlTVcVeEscHTp/tpfFMfgb3zM+wpbsKG7RsJiJ1FtAoorSdfIW7QxVw7ugEHecXye/KO1nkDHM
HXcQLHdSIV4vHhRzPlAg50aBN2s84nI9DJZ/7M1R/nQTIy2ILmfHQ0CuBXx+lYIZ50tdHPWnfXtu
ZlJjL0pjJbOJLyawFNfm1X2itn7KdY22j2Qlc2izrcYndb3JyuLg3uyTDFHfyWGD6cuuxKFGijEa
TMOqRn6UVTfcfL7KMc/aHs/FrFgMOGM/WP7NIu/FeMgBJsUlfs+cUEBfJqIfXIoY2p7V+6jAH+j/
RNq9rjjyoXWJ2FF1/VhUj8x6kUk/0EyM9hWh30Fd2WeUfR7nTAbLnVtEgYD+OysUK7Qw07cEvUBp
IyAL6uJLTlvE+42AejWw+2nL74Ykcnif40D2lmBz44uyfNRBMjdz03AwpMt9fVevGS+eZZQKyYrM
5TpIb5K8ZkIGFM0de+4Hxs8wwTv02x032q0Cc5oy9LVZBHJVlnBLgdhiaNopRXn0ChP2jY8PHnqQ
etmKlWrBbllANJ28b03ZLS+uTHYFKohw7FH/gJ9LUfjqcqarmyTgSlvCkwCG1oZRq301txMLukbW
tE8/nA2F70HAN2XhpRdURm1PXJBJjklhCeeA3lMFgkkGFjaHpRQwoVJD9S0FTvjryrXj9XPlA1hL
41MgnfuMmMW0vjC8ed74n2LJthJ3DBpJGg0R3PX5Zff4RCZ9mqTUdV7hbTgb9NSVM+8dSj4p8x3x
twIrI7XkdB10UPDjQSqcVjZXOfxp5Azy56LSI89TE5+VSTelLhTnVBvuO4iUrAj04xoEvFU42NEx
op0VX+efQdl/JFjBcpxs6VwQZJAcGkqgLJjEg4tSTvoTcEF3yIwp3YCcsdnWJoBLu3m82UfiUv8T
/Vg+xDXXETMXjV6C5t4oFQNhqXOaMXmrE5RJ2xoei8I45AAmGPzQ8zjgy6w2zAKld0E7GQ9lxTY8
Z0Cjp1feUBKrV4G/k48eo1yLo9tzjIEXEul6wumKwkIB+UC1aaG+ZcEiPr49VuBsIZgYjYvn7vKi
E7UbJmin0ay5/S+08tUjgNUZXId8j5XcdJybCE0CSm+S1qEttsDo0xQrvT0KzlyIe6UefpoWMAp2
cgmqLutiZHuII4xyxsyBUppae2TOIC9gRyzfnnYlBUQoOELZZOEeIXShPNbpwNu6Kh9SOY3cJqEN
0/tHfnn4CEHNVOEml2knbgDrAI0SJBSr134dDXdX9r3MeNns0MEt2A8VwAEbqa849d9ZhZylSnkt
Dsg0OYKPrDiDU87fvEnBusAzVYn60Zk9FaBgcKjAx0K+rk3rvAo2Y117fj/D9Y4vr9itUlFrqvhe
/Ixkh/ccOaX6k5C772al9a7f/xbtSFqdjE+lEIEc5OZFgar+fmLoguASJObnU9MQqBOOW572B4DQ
+Tk0T3Saqe/6hheizx3n/PnrX8vMutZmegrRoEY5y4Lt2ad61oVwbwkCilKwpGwCRLcR5F2Rsff0
EGhf3KfqAToUZHSux5PHk/JaD/wyaf5KV/pnXhiUCqLIPcAG/sdeujQYN46N+kzcmTjl279RFPpv
C0hFxa2s39YExPaI0MYX/cLlFdGlicMX6hVEz5qwC4i1HjNlFyvtbZG19GKfkH/sQ4w/y3PviDc/
oF9ZuVhN86Uy+zxx/hkqtYbe2cdA9ER6yc0a6aX8LaBcpYJSZmQBIs8nicR+0IYYvBUMht8IXu2D
GhxzvahaA8fYFVbjTytk3hLTAJ/9XXFiwq9srY05wuzQJNLU3939uIL7o/wO0aPXQCMMap1P+rsj
CaPZ00JaQhwmLRyQ/pMPyAAbFwLt2IuGUAfvJWhOqWlvl4NPphPB3K5uhIWrGR54P88zwRrclphS
juUB3EeiRb97pP0+vLicLzLnH6k6f5UW4v2Ms7H6BzWqu0MCsNzKy5W+6YdkYL23B3DXiclwe3D5
zq01tWAeXWDh7tH7+TQETDV2sfvyEE2rMdCdD6anIM2BEkEf5ASFYjkqb8U1V9KMCDLbsXKDBVGI
g9FPRgYOmEAB0DX3LUSa4PTjYOS+81Y3z7az3ZR66E0bWd6z+ytv5VtZQJF+HqLO1fxBP1gIORxe
a69mWCG7dXoUjdu7wmo8BhPepMXzMob36pCuHt1FZ6uxMGlTSe6RiUKkoAmPHm1uYueCAmkwHRRZ
5ibmr4YL66PVxmE/K9bvcvUSVO/Vdby2762tmlToEEGapHQerx92mOcOJeeEP4dBqKv20QyxDw9Y
79MGqtJusQCVz3F5tp72rOrKvSEfcC63GH7Au4Q/3DQ8psrQm6yXM7NfGGJGzxNKNvUJOSwR9puD
b/hGRv4KT2vtZGwrdwE2/6i1bu9yxD+JFTDnKBY8ahUwck1i7k9cSFBNAPUN22p+KYB7RbQVz+oj
sCcknFtKHJdrLxVQXempnltpeUmHuOaEKV5Hcx+NhzYFaoNbdvvxIBzPTPAmnQyVHND9i5fIrg3Z
r1McbLMVAK5YMxonAbQLc6ccpDwrgmOhnSGQnKaxqQs49p08DkrwBeyZAZ4qwAmD9EY93w9aMA4p
WtxxtY2oG31EyvXQ3Md+kj/Elq34ozExZF8b0vgCm5t1/sMCkQ5ftBNtjIe6K+U8Iawv1nlP6myd
EzFmR+KYGeBNYb1dUQUBdRoiYtTT9VtKqvE8lwxpOzNHQCHWjkw44bJJkl6uoig5AMX/QQL0gZhi
KyYiuuW87wrQaWGdSrRtGobliSVhsq6PUtG7GP2oAe9EvW9h3GJMuJXSp4ZW3wyMIcPwFeyCl/X/
CwYv30cVP3odIvzd5Ooyi0194tQR3stX8lEv/68OhtI4oZ7Bw3f9ieKOM6KzLbFb7dF0vMilhYCu
j7qCFLbO0TX1tZaiiHAvQXpjlvDjEzEPEalIhevls2aA4gBdOuze1GOXulrDplCXM1AyeYsFrj5r
5Lg01CJkpYtc7ldLDzkqM7H2yetLo0X/hQYDJziUv/LzHzIiY1bipLuEXttb90scWV//3CSSI3JO
2slwhomivezFRlvrAs9LvOL81OIblqI+J6hMzjIPnITRIDjA/UUM6WHTfJ55kHL/3RzfivOk7IGY
iqyhCpuR9yHB4nz7vAR0Cqwwl0CJP+msBOg/mR6IWGtrK4i8cfPN5Gpk9CciTRM0y+xsIeW3TGgt
s8IIoeB6OxvIGR7eW0MvGmnZyiTu9rwEzyikkdR3lyO0vXkyGFjyENQRTWYaRi70zdtaUXO1uL6W
zsDOIuRrAaQSjABzZ7bCxcCTBcrB/yIucgxtlFSE18TI4hNFSQD7rZbjRJlH7iu8fZtgxjCh5XER
vHh6/JM8pznp8ffY23GcveTOR6n/cu23i4OX2f/ZxjHMpCiw1X8liUqPnb9/zt4GEqmX3e8JHMjB
4Jxm7zFTlL6hIqE4DyKaa7EV0ilNVYdy+vDUKj6Dl7waaktojqvYcVWgivgfglzgkeotv9kcwUkU
q3AjhTz2GV8l6ZSsYMuBzv6Kcri6e6z/hGAtyRf+bOVUhqSu6UZWW1zjTMLHRA+MXgj8mz/iVcsV
1I6z96+BeBxTpe+divZqWpMxzkJq4ActfpIu5ueonyEwscrCgV013bl+dQCPs+FFsnAvjHqUDcTN
6wKtC2XCbjYDyRp4Oh+UgAl0PAK38PD7wLhvYAhHqYihpU+L1RQmEqfgDUvk+TJsOhPar6138wvd
8rvGsOteMQPya47R0B7UAs+0MDuz2mCU76F9/M+PoA7QAosLKO5UVjM4eAlyi0/H68KMyLF61+H0
MbUC4ioxpVWSKi1pL/Bu4XinvKaThFc/sXhmMojlvtukigP0WdwKdDt6B3oQsFiQyT0GiSVJud71
N3zs2luXbd37T/ju/F2fR9bkzEv/yo/4M/5H4UpBcYwxxlJxc992sco/EokQXr+Obkr3lL17BUqH
5mfN7l/QxR0QY3pr9E/dDdPlEo+IpVL2eNde4c2pVDqdHn2389MYibV+qOsdW0Idn6sBNApsjIRM
/VphgKL25fx6EUmNWTwy27+phkQGrDEcYvsGAkPVCSh32oqKqjX9jjvPzoR+O/lnmBESDKKMyy97
3ynPWnNnereHcWikA78mqIbn87633M1l2DHRW8KU5BA6YfJQsu6DdD2unnXCSENrFOmr4RIFjWUd
qW+kLeSxnqvnQM1OD3XKbOrU4bcEyk4dhr5cuXcQSEkHdATxHApinaduB3Rtev/1LNyTQBrNtJ78
jmyFIE2XCzfG0Jr2XLklhNBGT6LfcXdg72Rm6QcHnLN85wlRlV/e3vCMfMVgIunyX5B1Hbg6ODkA
QHRv7LxueThFfrO+hSFJaVsE7v35R6yZPKvjlCuXHxHGmEJHjVEHQ1GD5YI+oOznKZZqFqUhTQYY
FeccgEbgNoMJWJwMVKSyr/5TkDJv6yd0LbUDsDrubaSeRCNAeMaWUnCHD1z/kRq5Q9oU2LEsGkLX
E70TZUWW7DIDc+223YpdQWt0HsVjSwVeD1xOeughtEFD/NwyUw+lroWaXMl9f/IwPx+n8IvD//KQ
SLBCTAJV/uBefXlvYofDpAU5LvzjIgmK3EkWSwI3xS4yJ1TrsxT23vhScH297pmrNQRgbY6excTo
7/XcMOD/m0c75Xq00z27M+eisJsh7rD8RVFwiakLLHz6VgRK2Djk+TFEFcyknmsElujRkQ5hUbFm
vm6iO3gCBNc1kBTmEGEk30nN35LuzCl49+VJ7fLhXUfehlJ+Jd2iQJT+kw0Xs9sdEf3boDim1Xav
hnyumf426GnfuHzawyXzFLUnKSkxrFATsK/OOG6atxSOWr7AQR6n2v23xE5G83RFKoj6h9SReANy
K8gb1MO90LayRcxw2EZdT16IdDUNH/495cIjUQBZpzABLicTfdf2IE1n9q/CD8dX2UI836tO5ChN
1H77m2X9BS9QJjckXFqtXCXtNrXajhZ4/MyUWSNp+ocBbdiCEY7HAPJPb1mUt0RLO5PkEsf29xtn
9msAzcrbvc1HrpqEVJTjf2gCWoG0HUCnLZbJG2CoI8HhvUSuPeDQwG76WepI2WcYE6cfZW5CAEXn
apkwbePPrs56CvJd8oFybut083sNRaBu7RTMPK37cQeHitWZ+zwIUk6adKMg2/Vm9qGuVsIYeKBW
2/QPsQtxLCKLSG8f+qTsm6hEjxcabX0qNkyzYHoxvKo2Cf9epdOxtKC0lnjsklufGrDEJjcqW1X+
/Qa8UVwv3uByR19Boin5ERzPVeUh9M8NDB1cn4CYp659npLmNt9gLMNIZBnFwi5d8C7p9In7tsgr
lSGuZw2z2dJvdhD+/KE5aGbXpUI1DKlZ/5pP1Hy9tTLKAxB0ja5YvNUdvjBtT4clllumgMjDVro3
RoEKYxkplFhrFu1C1aUJI0aPrpan5hRWqvxQD2hISJ1vBAa57pow6odEjKkCCXv5lK9WovdK3tVt
+my4pdC6yhwZe68M5ei4eC/NU8K63JMs1LWUdQMmSaYWylYLxxBaQyrwe2GgyT3ooLJ9pcSOFESX
z0RiK76+yHgJj3G10lgxQlEc4ZYkug93viNCzfx625joOezGCTip9Rc9Z345RDt5I03v07o729V5
WIgyQlzkBErempGGoToHyE7K1FbylprUc28p3P4ZHPZlsfoTYG0VtjzYVzIBNieJjcZY6T+WglNN
Wa5ff/XmYgZPmZury1QgfY0ZXW4WIbd60rDpfYTtfoQg1lPZGze3ScQDKA5Qoz/0XSxFrZjzyL31
/t9ojL+cOzJ4P+Ky5yJwlH1FCdstvIasi8ftgQPQ1GIaXtdAiMZ2MiRu5aCTiLofOPY7PDOM7Plo
c5Wwpzzq8qL5k5ia8f4DT3znqRqFTunErQ1SDIkHg9khRpb1IxyWzULY7Ho86rClHn7Et6YmL4Rf
8eoVlU9tWUsseoDxMqBaHWVhXKjIL3V1YNjvK5XQK5/mq66JdMvF8FdDshpIz7tqRR+XX9mkEgjL
KDNFoLJOyabrs0v9rpggSuhoFhsY3/0IhIUqw7eqkr0nwKtAdBLHwn6ZXpkG1Wiv0o7Um8e+87IY
C1DkY+GbMjQeLhD/VoSiO1Zb0KWXQjbuj31rxN99fV+yTjeDG6SRfVTDcIpTt7HMIgs3Qu9AZWQC
x9EJiuiaYeZpQmWSy3Ueb4m/b/SlPf9m2Agtit/nE9mFF9wlozZ/kc29axMpfbmGIY756zqXZOEW
Wg1G7x+7Lv7XB5L8SnTnxXJkX348mVT3Kn6nhloYNVL2jFYNWXb7jJEwTKYgO+vfaw7qWa+VyF/F
P0kPxOYDn/NdR0set8GF+nk8H5h8uHzyr3s/l/kjAxhRIrM5Py30ljFt5ZM5/6PVj7tZ0sLGFgXO
1Oizv3HpKYNIp2u/T+7d9dfnXEAldMJOHUix8c5Qvq8hJy1ZqPJgluXZBeW7+FtygrDpLQsHXt4Q
tk1WAPdnkZHuwaymu9X5X8NTNUJB06zgDenHk1+zXM/V6ilfUVHHqOSXfLc4FsiFatTrlPR2sEc/
0jyc1M3uK9tJOEp8qPgiDX0iXRK54whtbhi9YLzs6V145cXZTd7XvZDZUiVMAlWHQn9VltIHCjHj
DKCrrWb30eUFVCxlPT6/R+cGpWCTFWiiA1CRV1iUe6v1cJcu4gAHJJi+btIA38oLwj+nPEaTqNwI
Gooe42SbYbFnMZ4gdbblusUPHjskbCdYvBqHO1YitHuauQ0zOE0Vo4QQXeK8JB7oLnjY1fUsBsIo
5gjuFtp5oTUnPBO17B/TKcInjTN8RlRviwOPwPXbDYYQLo9QsTER8rdYZhnuxhdZoxpl+Qft4The
0tEjgFQextAVFCacpcp/QsCwfFuUj/lLxQQu75y4VpsprQeg6jUjccYrBR76AgVPbBLb/Dwvxqe/
dicnJfdC5bNhgxzpOUpDJQI8apTrCU9He+OgO+evf/SXQlKkIZjqH4Hn1dsYANQtEEQouu61fe3E
Wk0HtJn1rUN7Zp9XXFJVZHPio/6h+SyLDcg7QIlsnAFuArI7NIghDiKxA2xYOjmDadKnoB/6tZPE
1qEOcDRaRi0hc9lsCBM2Yhj26VUQTIOW57C2HMjq/Jy2pyBeBqbNSvLH7n6DA4QhE6BBjDQhIJR5
rvF/s9UcZr8/6iCamKU3eQ44LV6a7N7esV+Fs3r6gFaP0krjria8KAc85R7O+l/OD/JL4D0k0Lg/
IvpYoX1SWbEB7EpPKABaxLB8fxCJ4uNODVnRpRKNI/dTWjH6Fq7JbGfaCcHooL46lytIxOfF2n57
wau1A/zsjrbPnGWz9rlRABenuVherkIWV6Pvoxeta2GhO7IVjh6L/Bx9fLZjiRpW4RA02x7eM4NS
IYj4lDppcqmW3C0D2ol55jhAh3LPH7vaNKuXdK0P6r1uhUM87EAQUTSydTI57OPKqzGRBUN0TwpB
yfB6ZoEEpOwB70kpCLL3YbDVeHO1SMKB/lScE/gIRrxN064Mo5GCZ2IqlXuXtcO8Xxy7CRTQM175
uGu3arbWJyquoFPaNH3czf9NiGdtXK6iEfeD1w5+G8mfOvEWykGENnhpRQltBFGLsGbUHnrzAu9r
x0u+REcP5vmfouUI8VLQO6tkeRHv2YvNKL1WGEiRblEKY/03OUowcGb7UKZ636h8zlz851w4J4U4
wR6FJF1o/PWZ/jecHUz2/pgJlDmsfIu30ZyCTXXxX/fnrZ3ilGiDuHXmY3i8YDhc42/IkK9rx2ui
wgUq1mbv1h9Q+1SGmSBOgfb4i74HXn+qWgVS6g1hXrcCXYrdg/5CsaRscShbNgCv+eQtjkJkg9Dt
vTUxi/VptAqeGFZIkd8ekgXnmAnF+BAIIl66UE15qrrBF4q2dV+/USsCL9AeGB4HHFT6ENIbGEs+
Wmz02yRTJw1q++kIWmHV2uILJUDNB2va4keHlSdQCaIEyk0RdG+gMY9ji7acTUntaoiEw+xpJbHo
W/GBrly85jZBoqVtsKeVtRHVhDc8kHjY6tgWDwvbwoejosaqCfRYXkvpZENv0VbMJsGnxcZd6zmi
Mjr6ptoPuA57qdylGkWlnGRKRcjQ7+OJu83l7i2DYWFNkXWERZPBG5dwOCsWDH6xC59prrTpFuRy
WuwsOMwRXY/CDgoRwtnc8o80s7MAAK836E86JMcwQOBqjCZImHSVlNeGc3U3CR1WNP8uCHe1nuwO
XcB1Oo9lzQP7pbRT0dH+3OIf2xffnodP268dyecqwNgimxaFccTBcMJH6DOc9aulMUTZnyoGebis
weKwg49elrk3Mvz5ON5HIE/Gnhvf8qOU5brEkfHT8DbYYJLidbYFKWB10h08NzD7UORcd0iBamVi
9p3NhHNTxJIjV3JJvfEAmXhqP/TMR/Zdl57AqwV7P1NSh8MFHOzM+6qXkCTMIBqfxumOc7Fzq67F
NylV8zBEZ29QwXK5OQwFQhylmtp0K6bHV5fcc6zRnzvDsaP4gWsJq5xZOqN8JF0U7sqn3QJeCV+Q
UBs0S3TGyCJutxujiNya8IOJ8bqIU4CUbtyhZgHXfz2IrtCkcapfyioBxOZNS8nRLPuCohOayGcY
5IUQk8N9ujbttLyKKZorQPuk6E5Ts2fBfF33Ti4h5b9GbZXzIsvufnSjYYtzOorFXXkV0DuiYc8y
hqRXL1AyJk+kgfE2wXtQkzwxXBG4KYzZUHQWkPxc9D90Qe6YIkiWn2pc4+De+Zkv2FSXBz8JQzjZ
+3osG/YrV4wvuxp9Om1NS98870+e2aZB8sIWgO6gg+C/JiHHETyj4qIrG8baHQDM1STegql0duQI
/8N5RUDEax3pSQDxo6Vowm6U/9nBucvyC5qqsVk8vVDJ+NH6+h1B+akHQid/PpyXpIBkGiLrRVco
3zCGeS9+mRboYOKV1gxy9+o6WSUrFff62DKNGfD7e4cfuWCqxhi27u2gn5FaWKXMTsQMvrsscKND
hiSZaqV0abhXaUd+lhLgo8z14Il3niaNqicYC3lq1XM+iwkFV8uET+IkSa6yU7VpVu2sbIN6N3Hh
OHZF+vURJbCjV7YrdCpRyEeKgYpuPMKiAiEvsUC13gSPbmff4NlvdfKRMso2Og9EheHqaQIi8qMN
KLhrogfPhx5d6C86xDVsLT+hOvqWGet9n5bB1LF+aK99lBcrUF4/3NPo4FHOGU5ZDyYuMRTu8vop
4vQ/6FO5pw5a4QQ8V+oFdpN4bW8M6ITt4ZOLihT2VGgqgImVwrwjWMPv0zYk/muCJxHhQLkEazz/
xS4lrNJ1G3Z0mFXUKKC0pnHDK+lXSgOpBasyZRxew3dXMhrMW7cNd70HW89cxWdQ3Y3KvnogS6O5
lK9DCrmpH0K5CCumt76qk8/9cNnEHKoMz7GlxR4jFY0rmlxqLToIRda+HdQj7aIClIXFkscBF2t7
dNn0oVg0ZGsX9OlDFJbi95BcNikc3DZeixTLqDWx/RSm40GaAbWlaEzCgRYmmY5iZf08Zt/BPL1n
DHvp7r7h2wlkvMDeyqAi0cb6r9O9QxYW5kLjPHwYENR+17IlmKaYzBQTAFMQcg608hd7FshuRqfi
qBIDxPWRgAFOpN1XE4adsMWqfS6oCn1ykWOQcg5vbPxw7g/FD2pQJT7c/h6bV63//LZ+Zx8IT/Ku
EY75CRYHb/qhjMA35k+C4O8k8vf713s0jhxvumhR4NuvL1bnFUIw3NXX9LaLmnSI9u1wzzB3vXAe
b0XnVGt0agicqJH1RxOOrKW99946YxQLlxJDbaiZq8u/VD0ARx0jHeNLxKWfNlHL7rz6QolbWedM
OWIeeXj2GzD/LU4dDre7Rn1nq7A1eNL3WrOUV4sWL2egwBE0JW3Dvb9tnN1Md/PsyO20PFNJOS/5
gkYVKGwPA56JKeI/qT4uPEcCIjdsFsWyjUckp2w7ulWkT/Z51wCg8d10tsaxLIucPLi45yXOpDtQ
i/vwHyf0k5H8I/lfzMkrGvDzSCSus7NPmh6vYg6IstT4VL3ffAqateM40TBfs/PwyZbJmVx1UWl2
/gz6br1A+ujGa8Wx8jU33HgmrVkwaXvsMGr6ohLO4WX26f23OOQKIfc/V7xavDRc0mjy2VnS9ZX7
MQ5NWC0qZGqRyj8PsqU+1khCc+p6a54BUX+z7hm9rSn3gI3yuAGVLqmO5kx7sW1+OhC180y4xT+5
wk6bpPd/NXh2MOmvVH77m2IHSUz/+rFZAmPDuvGSGkLKp1QM1N+bt/aqRg4H1JxBQpHhUQNqmU83
iMPWSF8nbYaHqZ8cuyy5d16SAu8thdHqGtv3SuX1vIkZwJLA3Zugok9MLiSXtxFXLYh6aTdnIxZq
ql+e5xlpOIPEnJWuQtIZti2QHu1q8GRNP1GeDv3MLGtVWmzA7KLwMSNnqmDDPw+iLx+QTNLbRZG9
Tbmy4xAE4I/gKLQztyZtqDINDAQBg3W3cLx7ZlK1SPciWW0WziH3Ztxx/OnWZ7Cj3qgahLmjbsLi
Wxk/2RQ0Ra0RoopoyGoQgrmkh0Y0RtGCpb0TROd39isH0BViO2dvAvyOkVMnNAijHQpC4Wfo3uX0
I7KBN5NTurHIoY40iGyJpWchFgrIrrCySyzrKsU9Dp3npw3FflcNHBGUisnVGOhpd1M5w6ZJXF2r
gwFb6G+L5MHy/Kh5c+IQ5AqNF7sTdTxsHPx/MqhPtELo+gKyAypdKzgCZphE+dNIU2zxmFbSdYQe
svzoYnG2WErdb8vZbc1nRgQzUkQIGNnXTAAj0cizw6iYHFot5JaltQbRXVrnkVhENiLj41APSvJC
rc6eaZ962D3ptLxmWOX9UGcbjme2xsBl7kmJGhaBNhRkrjJRK9pq8o+tX/fJqzDnXsSsrChIifVx
4YGRIQNe1uFpt51m3Xw3cOXIxxdNrm0CR1V8Ko3d10yovNsAGUsYxelV9fzZREE0c1N0YIvxstM4
vfL4L31NC/7KIfpcW1k8GZo3aIaBJI8VF6ujB9DRQVhqTdl0SqHruH9stLjJ+Mo2xy6cc9b1QOzM
OWoHypJerW/6EIt0JgAVTghyuW0e+ZwFdgXjdPs3HJUi8wPkNpo+yWOZHJXs59cWzeiZIGIu5Q33
QX+YdI5Ibad9QzcyNN+xn8HvzHmuqA1QUZmF1ILmys0XI8V6RFmtI5EYST1R9CnXQsAMyJKZ+JXB
RWdIORefI1JwiStzMDxdT+7ZvYYR2HGMe7WyhZEte7F8xqw8Z3tOPXvrUWczpvxKvWooNQ2bRMzc
+60gUe9QWRZwlxi+jh2/RQRdtOLmlj0t75ThFFgp/OriV04HF1bubgUhQuCH06J5QDI33yvWqDPH
xtk7eiqeXx0zqjKdTinth5ozP8yMBhDIBeoQ9pmrXJpHJj3jhMPIkYtLkId2Onqb/iG9hNkg6714
DhGbLW4A5iW/Y8jO5Ilxsc0gP9iFQZVARkEnAPbuobAgJ9D18c6e/vXwlDM0XwXXk3HAob7GZAKO
oYLxhB1drA9TnvnhAa/Zx0DblKKv/hhMlIrg+SCyVh4cVzd86AZV4KBCP19mO1gs0DBHRVIDb9sF
xVd2NhLrQfjxP6r5K2GI1HGN/OY2tT7CQjxHNa1gi1gbRm5wdNXN9mLLyKb+qPJPLl5iQ9Q5G2co
pg6nAt6C589gi9AL1wjwzjIo8Xq9tGMppfQXj59cy9bTLbpTuDz/QURoVrNagnSvKSzz40uUpzcg
zMaqAEntgwW6uYhBB6JffzjiXpzcFnrdQhIHgN3cACEQnSSdCpsz3HebuZncsX7bRZ6JmZ/HnWgP
L6A4E0V5JA5mP4jrewuXwQU5lh3AahBCvu22Ye1knF/lb4cCAMQSm7HhxU/WYUVm8wgX6YJ7Yql2
6hZTW0Gx2cGeEUv20jO9Z30J8ZH39J1W2/vKC8O5bQGMw7E1SlawaXsDYIkkf6w8IxrI1/EJP5WC
itNpxM0GcbufcGmorBZQEHSJ78P60wt2YneK6asmCUyHq97RzWObHHIvfuepQOrskSXtTZ3nOJTW
qFlJ9eSMQ/RmCk440c09PNSX5nIywcBy8Mia9Ze+uy9Ds/I8jXcWdh3Wvf6e0k8L8rO8DC3zZMGN
ID7FyJ7CCV7XEPhQ2YCT+I1zcf5pB0Ok8AoA8S7ePjI/9sI1WTC8PEkD35QGJN0hs88gIdMzSv4+
NDh5vCcDBycyG3fSU/uMcXOdeBLPY+nm1zBAsGiOrKRFlXORD0UxbnFJQ8oZUc24n2ZBE06s15Xj
OUtHYI/7SzkL1yoC4oTRVoFt3vdnEA+bV0kkoBf/M+w0Ci63GZtYGHzhEJ3ZarVn5hF5lvcT6P8J
CtWVFVkhV+RKXzOwNzhr2ZFf4cYvQcBNWFnan9Xs+jkXzJ1AMQHzeR5ZwStKKGK1lYYNn0s48y32
3rFXGxJtXNJntVsxC69Abt656KeBFMXQvfEIxC2hGIuTNXxghmdgYcDe/DHNSybMK66uimL0DDDA
a93B2xAsxfQO9nsUIbQnjXrf44dURiIkW6Q+rZLqBnM+d7rbTvTaTyvoX4eJDGxVUhRJkG7q9PAf
rjXzr1mCaDpx2tZllExLQoQe+Ppm+kO6uKOUQAw3qWLiv+hNFJp6xiIG7Qe7SBbZKxxZwZiWemb/
fFEVvej+ReM+UPmJ6sS0qhotl+4Agq0VxEsRY0lW6txthF+AauVYDSYo3xNpSl8d8jHYGG05B2oW
ThvLIrY0mGp9USzczzM4dI7Svmm0qpfD68dGYWe5770dr2KC3279N3zpU8yeem/i6zoVVFJBX2Gd
cYmXcThhCaJc0r+o0lygYXVlf1XXc1BdLDJ2iaW+sgXxIgZzdsIbz4YH17MzQTzcqasKUgS/k6Fu
2mkrCFAyz4D3Vie0jDFUScR5pxT9LFHqKkumQPMklAKgNuh+kVDMTm8PzgRjtllS1t/2g5TgLeaR
kkvC84PTp2GGeh6uU90wOxwteE7Qw3VeJCeCDHGQSHaTOXlZNBiyU0hwfjDx15HfA0n/VnaNVLxp
9A7luSIVvIPrHK7VVau9p6IlZsNWo/SPKQrRRS7sRJDEy1jQBH1txYFXPcykk+J7PCIznCKJWB15
FBIAeDDt1QZyyWljX6GOuWhWD1xLZ770UK2YpzDuI7HO7pe506KycNvpB8oSTTzk0KPrcMwKey19
i6gREXAq1wZDFqEdWlpkARI/gw2D3ELNasSl7CWliTr7cVrQn4w/mB0f7TeO2AN0cuuv4moTQE4Q
IJ4fOLBrZleHTaXCUxA+GEqGoCnyUyLARqJBOUZOrmer9evsbh0Q/A3GaVRFUkguDjux/rkobwOE
ZKqn3RQGILfGDbHSPzbhIMPRC4PeqTCxc+lexG0sqWL9NX+XR2khbeZcahanP4orP9/Zh5nTdf14
vyScqGuis3duHGQ0BeZaqQ4wJWhScxFWDC/Dz2GjYVae/SWUpU8lJ+eJ0P8JuPQSCeUPZzIetb0S
19pIGk9/+RoEmaEmjIb2hVBtmF09UMvkdI7nSkCtYOJOeHoB34PqUTdHfaHFS4/J/bp1FjHmEy/b
ICnjkxGlDTW/0EBPFtz0ySe16T7o67JUOZRYpv99D/sdvbt82ZphFT7Ovw7n4iLUsF3yUgpQQxr4
d2JoinbSxtDrzu+fVx0tBdKJQEspyeIFg3w63a1EdAjiim4NmYdSJZhy0j6SLd++dh+C8gWO59yj
fX9F8g3vemlfd/LnfUQ+NbuS0TRRCyhhWGgfIn+PsDlK8FydnwfmDeWxGhywZ/lvdHlKFdYBHM3K
bs0u1S9s+fjWegkkP3OgS6eK3lB+z51YL58qdxpW++r6fFP7ftRkwuoDh4QYWKCaKgUeVVpL6TBl
+XbXUxlu3+TB+jKLXlPufU9mmzJrk9CQcDJEQekeDOXkxIDwdelryvb5633IaWhV0zMOuzNrDmrY
Kih1JIWd9K9LfrL8aS9weAwdKXP7Kec7Rkw6OsAnonuKGETcxTMDtDEEY8yWDQqAURXw7RMRMruI
M3fPfdGnC1OkH1Zk39jwm+rro/dj4ZGJGoOEnEWkJd7/mMhH7h/dGb9seCXSHOLehPNAbop3Qqhg
v1dfawYAZuZf5pARYn7fHo0K4rWmoUUIWpEUrQSaHB4N9X7mAvUiPyQdmDTK41xm7wJdl+WS5x9d
GB1BhjcKacDAdthrb0r+tsAjKqLYBWsEf9k8FokWLZZUng6YEIrRI1Hn1TPcWYrLUfrGYsB1pUeG
tLwws+mHQE1bLzJqxCCZLtui5/T43je1r/d4VRkmqxdatQjNLExbG/0cRN3t5NesoND+oEmmeBRZ
JOdQIOW6tNAWGOyKOfwQ6gyOiRWPfbdKhX/GEHdR7sJYL0pfvC7srcabB+XMOYZDXuD7Q3O9sA9S
ZORUvWqweETwQKIsRvkVBUOsSeIc4nvGEbPrwV/bgziVHVaTbGIWxwg7y/bSlst3yMnvBAq4ftJT
pAGNJXR+ZBKgxm7QTfSaOJCeaeVV27169AASpMyK/v2bdTHXC9JB/au6larRqdQYLYC1amO0gwFv
LnrvoDBJ8QlsGDavd4esWGRlA2vWFi5+KqK15QiDp9I+IEtJVxeeNG4mepyZBCtgTgt7LQ8BA2Lt
XGW9DmoCmCZXela5Mwf5sp1saAR24np6xUf/GGZeDqLlrIl1hl62gbj3QcRed3LmYrwXAgt+xfZo
gqRb37uw9nR5rSZGnlEnzND/7DNAP+p6svw8B1G369L0ZwF4uwGXADHh+IeaqkEs1XqE7O//veMR
hoBNmXiYEgD2xVCq0kQ4a9/gMe2Vhb3Cc1SWZNUBc1kxKhxqGNFU+E6OCLP15EA3H6HSIoWMnCL0
4dupuNr7vbIO9sSXxYB4tlVUh4the7I7WSP5+wjkK2kXXmIu2lE10V/P11We1DyOLNAuKl1z4w5A
9W1w9JTbQhRBrua2zdXHrtPFP4alTyS47bm5y6pIHLplRGfjwUjQNdb5XPgSrOTiCKVIKTeSjNVY
CRLAEiQZMrch7ht9UYeYvK+PRe6o5oE7Eywi9Y0J8qcspLG3QC93YNgl6Bhyo36PCade0UPNojFO
I/mgDH8TPQJyE8TslfC1B9PQTs2HU0Y/PkrY18ExtahXcCCmiuyO177Yr28dbBHd3TbB36SH1Lrj
Pmiz6tM1ngc/C+be7m8RlugKsOy1pZH4/HKLhNyKkODmCQ5eeEod9B0n4H+Q8KauXpTPFTbKV6HW
fDQC/DpMaxOTAHrruVWvs5LGJ88yDIYdxKP/tNYOdW4V+mU0N4WhALK1fTUfBY/oM7t4eWnaJILr
s5G23sLuC+BmLl2t6SjNFIT3Y3CTYYRkueB5nMLMYdRDWigvjMLa4ihICAQMGX5m/Stlx1dSQ/Ig
1H514OQTVojZU2oYjQwOnyQXQDHqmW/4ny/PeqP/JhOIjg9D1VFJoUJtHWCClk8nwjSlcNiDDz4s
DBnsYFiMO3b0GvcRIiFtSRySyRHGUai8k+JCWAxu3jtUMYe06RVo6F2+oUBrVJhjn5L03g7nsf5n
RnMHVGgSFU6btPzijLqWDKAm4sAN1ECmwi2VShLor0gE0Raw1S8HHFVkW7ed6M63DpZsCJGoskbm
PRqc8JFK6DDF6Sj4zBWCmOuU6R7XH3eDa8y1SNVlnQqQbc/7yEleMyR1D9LLQTvMXCJiHCw2JtzU
55hcYQjR+oZmSAzi1mj+Ev8acFV7FrS0zGnp1NeX9shmbL7TJkco+kXW75pNOVD2Qi3QMP7ucSVA
1ByS14k0gSVl6mm9Dvyd4zZQIE3cxATEuSkDYw0g5WD8TqWqXGr9PCgADZMp8TolGjsLJxOHmvkL
AUguftgGyUIgH3Dwm9XTYHF6YQeGBnWnjSeZSu/HlqtCO1f56JlaUf8lf0dyjSJw+0YEv/6vp4lr
8R2HqN+AZpm6M2kxfDHlOhD9qKmKTNCIUopucZNqA2R5Yp+PL8jYEjaMxyBFLwruq2m4p8bnlsX/
puPZiKJSQnT183wwIe86vLp5ePHKM4VduBBEoK79+8cfBFsgD7AwXDvfO+Gw3UwYsG2/8VK9W07Z
GAbrfSf1bFy04kDa2XQimbafl5cLOfpgCHKOdJR1yybkppbdp3SFJXk368rOuiz26UdZZFJvwbEh
fxDmgEcR8gXRNnU7lTe97NDH8zuPSuH8CE4gBUFOfRKqMNbHaGXZ4SiUDY2+Xmy6REoyIGZE7p46
uhJ7Qul3U0AE95N6MgRp/jqb6QbLK6HIneOjvs8mHhQ1R7er/545S2DJvlNgP7d8+xrSFYYVRMnf
dnzRpXktWWzkpMYdInYTR+++M/wdNjvmQ7SskRnjbcszkktNR70FDtOhkfNwPRLlbM05UNltfODN
zmnVkv6hIrKNMhA/r9jCp19Tj6vS/k97I9v7B4MFBAArpDWQXwFM2RdyZ69vx7WKS3ybabTBp2Y6
a8oN57h4N3as4JwiKW+PsefZ0jJf26s1pla5wtoJIJ5zQPSn5QTmjvDWC22KCRmU9b5DdZN24n40
JDJpFHl5dpL51oJs2xKBCGi89ie2IL6gvB+3HGlSgFopIhFHb15IIpJ5dbKOIiaryO5jAWbXThA+
SQfYpiZxW9Qo64s6+hgW6Efri2jLPdEKhGhTqsUA+znCyX5v9m7rWKEhH7hi9XP6w2yTytO1tBaX
Mkx839XF39f6wuTKYQMVS+QUYsGh4Y8l63K4tZw6VCtpRHzIG7TSTeaXfCE9i+RzGcIhG7pTLOQ/
v++M3I2CvU9Auu3B5OVoJ40BKUg9HilkF62iKyU+zFqegxcQzxesi/cnr4LfCtRok+MY7r4f66JW
gxfyxSEAPj3m+31FBBu4iaFdvL+DOc2pUJ4y8SNXJWvm5bQB8mJa7SYgxNOUvQmTa4UFLjY11sVE
RZAOhZVvCzMhTIT0UTuCupp6zH55QRcetgYNSLEUK41lmRjB8td8ZlQ89bApOPJ2WNBBzZxa5y6/
Sh/9RfzrjxP9BR9u9zr34xZFikL87jK44Bh+7xusjBEIf91pp1odox09wywZHTSxsVIgrXpGkAh5
zs1pdT5+LuAtdn9Z3XBgpPmlSkDHzDvA2Y2LMHKe3oqGrEUJdUcPsUjCtcO/MUWHF6DwMEOOqcUk
7q2eqaQoC6BhatmKCExcw69ZH93WxAjwkTesqOAL1l/2DOxtNjXF6FSflB2ipP26P1GOA7p8o7N7
Bj/CjgH/5G+ApdZOZfCVMbijAS5FnJ3wXZkExc225H/O6G/1Xu9pYAOaoNls1PLNp/Ko+q80/opw
lAY6/WO0SHpbXYjzneAfu6yragDL71AxL7qt+vNJT86k6DGtPnxLPdb7B0BQ1gVAiNAS4K1fhuP/
zrUtT2ZxGx7gbDKLxRVOmdWP3NU3H1FvQ0dGIWSuIyvE6IUWJLT/IxLrYqGyoB+/nTEJWsWG1Q9Q
/XvHB21L4YZFB0X7HZjvA1gVN8qd0K9MDJoIEopTikzprUigdv0ZOql/mxqIb+85B6x9WuLlME4W
tjPCx0AfmOmXSSBVUd0nCNBsBIfEgc81iZrQE+uucCxt4AmOnOLsTEZzFQ79N2ViiaNVb16Bc747
gAPgOsEfYkt41pJS6/xkLZI0kErFfEp2s2rxVZ44LzVIBPh0by3y13Pc5w1KeJ2HLcpbrWcS5Zpe
rWkk4CDPKaj6Pe9Jh0uKjoNHp3XoAFFiBs5HU0rphyNRxlexmLfFW207aduvdAY3QBWlLc5tVp2k
s/JgNXc8TsGNDJc8WD/eLpUzOO1hx4gpPxzUHC+P0oWB1LDY4ruSoFZ2IwOkNg0rtNZRX9oHIfMZ
k1TqoQODRhWht0k82eSa6/ol6nVW+13owdzGumWPSWtAMiYVjB4fB7HHutE9en+25wfR6llbcMB6
78co1kPi2ZxRNEuUp4RavRtW2lBBf/5bpVPV99aF+RrEW4xI12tCR2s68R7QEHOg7FUCqNBJS86E
al3/jNOvbj5NmUug70uPucv41AX2R57dInTZ5Mjwg5szZcIkK78hEZq7hK0Raf5GRstZy7L3Ke3B
7XbHOfAo+7xsvQZKjGeUegdyR1y3zYML9beGbfrJcb2jkixPwSkUnFAajoHDkJmfLr7wOeJMdkZd
eERi6iIbLutT4sG/4xTJmHz6JFUzqTawNC87P4CpFmJqkaSSgLucKCQYys25Tf4+4XFdLXDPleRT
culwHMjTy6BLF35ulBY9i81Y6h99WhaxfkpqFNeKtC8MVj6wvywL8nAVWiHN12lTyx6762rBN72H
uQ11UfSOr3FmTp8hEv6uQXP/uXaEndSUC+kE2X008iY8Ir3l1/895faWXssxpN/QnmXm9rJXI6yt
PS9z2nzSW3pjtd7bnTkZ1RMBNmDPJWNnykS7xGpYU6zc0z8jYGAneNwWv8x7oz+p4YRMtd3m91i2
FglHF2MOP9L0dujXo3abS2b2d4lm39CCerbWFcVEHZuRm7GBAmzvdVFhiQIIAMZKkL+PVuIZ+Ptr
p2wSVJJozvQEW3wCP1xb/k9tw15xSJReLswdN4a70/AEqA64yfoQZEMlZ4rY6EoZHOSjaDfzR39/
Hewr6DIlKsSeXpKKc8Ovi1LVL567snqpmh0tjFj3/wz0DDM7l2yYidmbd30T2r/L7+0Dwm28dhEj
srUa7xw6KlopixH4tWxK5ebd06OC5iNVAW6pM1BQF8W0FHbRM8LAL7I6X32DXgfiCf1fxOElnUb6
CtCds2A1oPcQ/KzJ9vI58Qv/XLkdmmuICPgntIAeQmkTqoeq4TZ0iiYkxwU3ZhiB7LAYV3HXHDbj
GjMP3q/Fl0K912cxoUsN/N9pfGDFIO6Z8oaDABmCZrYZt8BM/WFREdVYTXtK9VqASfIi+dJpAjKS
TWwDhde9pXTgZMpFMOMhzfRlUqJyAs9s1Bk12hLXflxIicTcLM3igfySEv4ceBa0jOoxm7z6owSd
C7cr7I5X6p5+IkCkHlCrb9KR4vLAKOzvbtceKIFhjytgbBMfTW8Px1KIJBKOLCUNaWWF5++nIF1V
QpNaCq+mt//OjmC0KVjVgCR4gvx7YYqsPebKtWqmw7nE8mSKZOHOE5oVE/uReZ/WcyCj11crx1k5
PfCFrO0liuNXedNCRWI5A1/Kg+pzCciDzxcqgiN+b57FIdNatq7A71/vaegII48e8IoVmpOyUW/h
c2ehV73222IxqCgHhnRoL4vzYndwIEMRLxHvUB58o4S07dEzBgxA6GlfASyEq4eIeRbBJK9fhrry
J5EuNl5t9pnecPjZX3SXA8rlpxfLvEYOkErNTcu8DtJjHo1WAjtKP1ftCeZz/ipM6L4CfSBwS4yv
bFpfgerxugAYN1/WlnxTYKKRHo5g5e1/jYhAERuNtwwmmRkyybU/yKrbKOWGCwKFYDfPtELED3rF
JkTUfmvRAatczUiMGSNUjWjz6imapUJ0VTrwD3fBsT/GGfg3AHPE2B1COF59+WwsLvmI0ohMxEy7
r9ACLLbXBpsA+1ylfT60JqqWgbv0zcYe6x5tWPa6OzFuArvNjIvqyGZ+/+T5a5ESuP4OP+pc/098
FwUbLlI8xYWKSFYqkvx6/rlOaw0UKmiA00ocQ6olvDY39sEvCiBTsuuLX/a+PiPhGDyDtW3AA6G3
q1iQ0QwL9eGt4uUcspRiU+d4GtMCbZhKXKjOiGIQqEcau2g/r7knqvrCndWYlM+dqR0DanglbpP3
qK1YhI7qV1aVmvdmY2+RVjr0SEuIMzB+HRcpnQDq493hjUuUNAkMeiEeS0I9zqfx1oAz9FCO4doy
UZAsji8eZQo4gwZokglmopHRBeulGAS4mx6gH8zMRzb4EO9F8riCW50IIZcfIkh6s8hYzrj2cslM
a70MJqIQPL7TvAc579UAIVoB54L1Er4XXhi+g9eloacI5T3K77jl0nnbWw5xwv2oyfCyKnZiLenD
tFXs4PPV3IWk/1VHC9aWLIKDmNqv9nvydB0mB545eE4CSK94so1zHJk8LFiRcFPB+Z/BEWpfZtME
4GIItwszxh8LfcaI6DbWS+0ASwIMtwkuoCwP0zXF1wBYuP4j/Cun7X3DGuJ46g5HNhEp6JDRI9e3
pKO/MzyjJZpx7b3CVK8iNQieT3llW5jttXtKr2ZeTVBLsS6FBgBGc//g/KXu1UjFx619kxbY9+50
KITuvW4ODVoPtzgvqa+4IIbfJxv5PjMYLHhbHow3q894KPSL0G7Tgi5aqs/UDUcgFKZGTbUaAZlX
F3zV7u//Nf5ykdSsVOHwz0le63Cx+AsvQrbuQBoeZc1BZik4wHkWRzRGZEhwr2XGJdNYVIfcHDOq
PGP+hxduo2/1qt0M09u1DCOtarChkU4vPtTVZGQconjJYnL0ggoeF41E0+o7QpGJwvLWYFavqzJy
A51D7+DTVcCvLMBAradJCbNDW3JLSi2+Es5zXZ6yoJpeSIUvnCKxetivczBARLb/ILGvW4zrIu/L
L2OjFexlA8fd6QSRquYFQXZ+Y6dBbwGM9gd+wVwl5t/rS4BJR63vJRpPuiSuSSW8FYxmpFHO1Hdo
kfJntkdXJCh/M1MW+80p8vWHiLaAiGn/OXWnhaDLguWHDV/8eQwUGc00Ppb0Dh42g/KI07/yZj5y
LjHVmcBKQnHqCeX148rnpbU7hgCpW1lCRLiwEJjmJ0i98MrTkkWSYpjtr1nXNS7ZgM/S0DTW7rV7
5vPRTiTfsR6ravbL+hm5DGrt8Tc58Q5jQcKuivRq5Rj5WtqDuI7LkWIc5ZZe5yNCjHRXx6y0l02O
BmhulnIQcfDrW+Xf3kiZjMfn73THVFvZo1qe34cidUxJ3f/tvrdvsUJZFtt+JZidU3sA7Oyf234N
J+k6QQy1ByM2w9tQw5HTszul6EgZIal4c0nCuK60HDVyVnWEE2sOd2eSJgg+v6eKEX3SSM1v+5+H
R3HvapdoN8kVgVQPG4+zZfy6M6/X+DFAc4oKuUxrsTqppe+O236L1UjFkubZHOo2Xkt1Sg68LDUA
0vzFIrnwr591IFgZJmFsseewQzu6SVoPDiZY5s6vHmHCK2Ry4OmZWrULA7xynZE1XRvSf4mRVocM
M5gJL6pUwFR/hRl/AjQNfZEdCYR1L2H7eHK2rw+KBq2aNiTEFXWbZuYnmj0zKGlmxHMjP3q0hho5
9BgYg3fnGs3XV9Q+kbrT4oZpIw+mA4M+8EL0j3EBslxvVAi9RrCPer8lsyTA+W0lu1hHRRLHB84u
JJdH039pyXA6ci3oV3gyZShWr4S2qDC9jT/hvaDt/66vajCbPq7A0K7nCX/W4ZV1qa/FE8lMt+Eb
t4zzW8ArjfArODwLIOuLdI15yyrixuj9blIxeSRv1DJZ4KBkIV+x/uGXyvvPGufaKyqFn0ueCneX
YnLeA1cWm5owCsYMPe9jYOO/USxD5NUcI3d+YgWieKWB6AzEfKDGkI1yjP7nJNt6DgHADCS5xbzn
Qh59UOD3cS612STzQAGlP/dfPq71c5TpzkvsfFsJFJlGDA5G410TQUaFA2Qgx0QapM7hB17JpYXY
d/AZgKtGSGcdtz5R7GH4wx7aATSONfJolcVrWuehJoL9gDL6ADDbeNbD5uzW1rNiTvY+rd6uZ4It
nKnhpGvGb667qZNtCYvatuZTRF8MqZCFomj+MFYyCm+MFCNo7jKvqmdBiTUiB1/UWS/iXVczhgTH
zPp7HKeq3hgm0PTGSmh0HiuIXqLaOcy1zcb5ntxQgRVTxdfpWIVWBEngud+rODlpn+o8rVdQGStO
oKqqnjz/ezEYF5tNfuEwOLNu90YKANYeuFgNRPboe50AYgoYaCffNS7DVM5VgwBrU7I9xoQFpqFe
0M0vnrZ8mVYYYiwMNyMYTUVnhY1zEHB5fHbsm82XnEi7tk+Xi0gQRsTxrRfVsOCqxVxL8HaLNLIF
HfsROVCqXGORTTWyxLr2Xo5e+AULdF/5AfTN+VFsgJc4kjxDM65KmJN9figLg6fJWFMvf/0lDcrl
REL8eOVIkwxZO0LBacJQXFhYFWcZrw7yJhcB/zPDD8TUzbGlRYtnchpPusjlfEsCaGzzvrVqvCz6
pVLUJjLhPJJWWbdg/3az4de7XhB/XwZQrjOEJxXQfEzcSbZFyRXxBrrzZrfwKz5Au6V03+oKUhi/
x7UdjNF/nI9HfGzkMu7yJgfA8NVGsRJA5UyaJZXFy2LOtTCI7Z6Zc6gJx3Ygz3G9k/MzQY7paoqA
tFXfsM5PaUKirW6Po0pEFJ16Ssbh4j50KTaUk9W7Ctt3zE0/PA7NXEv2xTKzLaAFOurEHtHdK3kw
f1CUlMqTxNyreUabp7EEhcqhV3uzjxuL3GfTauYnFv20uvc85sOjvk6aJq0VCTZA9ww7VIa8obyG
p4En6CUY02CYE6Gh06uCXJ+UJJrzdQW44Kg3+q05dg5ZSeOFs5xuLPsje+nyo7oQyCoJu4wiAmX3
/1uu9p22PYJJbJiHzHx+oZbsGz/F9k0fDXX7YdCzTYt2N5ZoM+Ck0qPidK/rq/KRxQ9AzPWP6p7d
a7L+xQUMLo9mrkB4hXntEoUJGL8gxSoRSu9vgjcEZWW2xtwZtLwskz361fNhKwKoUTMiYycLD4sH
Gyu0UCCXuLAZxT4XyuBXqG5BUdZVPIT95aMBFNjFVVfRb1CSIgrK5wiicj5sd9BjbmmKvkT0WPI0
Na3mT4poWvEcUz8/Jl4Gdyu21EYxYawsksVjyJopkL0r8Vhh/6xAeSEbTSY5NJZQj+5/XqE36V5J
LCzGIKddKsE4iwPSLIKCbvT5mtIgXe5391AQVMjbaJA+h26liEVIxtZviiMu4xJvwFbeEr1dC17D
54DLRDSuCM3H8hnoeElHWJfGZvhfwXdUsfTqGfyCQ7FT0mmhywurva291GDojrxo7patx8dvrmN9
RH+gMakRdgJGUsskqktkqeeZIq1QM1vJu5eWmsDqsXyHt5TxPg320W9leAMxLvIWJC1lR4Kqc53n
RGumyqz8sKtROJIevBrYq0UlA4a96KnTOWaKUcIdUvZl4TkFB5NtlEpwMhfVPi0SpVgCDq620arj
6kDQHCmgJuw1YaUTY0x8zQOB83kh3P3UrMvOcIU4LA2z+7JIvvjmxgfIfNjNS8I2YDyspuq8D7oB
zzfXrH+WgSpElppTP4B8mwStY0qy7vNqIZ3W0xH0wPBzm909JntkNZyIyz6hn/NCNopH9R7g5ZA2
m1c2Y7y18HRlb8FoEFJj7++Jc24vTwwgFuFNiDAntsgRzR2ck9KWg0C6O4IG6S07hGMh36lrCRl/
4I95P3R8Z6olI7eCUuim8zrcV8LwRgDBa9YbgbEfLFLduqrRrhZ9rRMjUB48pYcv4z/MhOEbTjX8
tpE+okDwVUCCj7TKZU+33NlBFIjK5PSJKnDMW0yIxIg5jXjspiZOGx41vvyoCk64UTSgZFmiUcqA
twrTeoyydziPHQSoQEp3oyV9bW8pJ+24utffqnXMDOCCnOz1tdq39pawzLr7biFXB4tQsezm03Bz
S8vC8Umwk0ZwMKkTBiH6IhCCVojUlVQ8bF6tQ62637nNGkQayrFlAfSQNZsdzcEh31hODmg9NO6s
KkTlkUETlHtjFs9W6Y2NV/a0ZTGPjYRp/LI08KU+n9Xp2Uh0+j1yXzM8Sl5ndljQgMpg+oFjm/d5
+oTuXqD4ZoJ6kKaHJHePa87LwVzIKNH9dP25sb0G/ZsFkmARKCoSiIYivIhfMapPjAISd9QPSvA4
s3B3MIrHzqgRt7jozB/KlaM4VD3FFgOYFHGocHlwb1aMNExBLNM14eog4MXZP/Io3uWP/MP8Mz3I
/rtwpO4/IWDGkptQMSWW4+yagj0wg4QC+MEYi8ozz1Hj7kJjXRqWM5FPR8wXNKKWpzkGbKI4yLZl
8kI1mPv1XlzEkQE/YT+GhGlCSJWKy/JDmlAIXMi9tUTFBa/bNx+m+HQKV39Huud+KfUJCq+MDH4d
Z4IzYKlr7SD8zyfm62D8enm/9l0frwe4Y1bh1wTIB3Pk4woQMu4AWz6JnGYC9O30gUfbkMXsrrwG
/otDcURAEoMl5/zS5Wa6H46RKVFMjFmBiAzehjm+s4ACGK1l2bR57jhN9MS4slODeTidn1rh6OYR
21BQb5ICD25Kf+gCT6VuEhBFl9WbkwR3WX6DAsYO6BJ2Em6dyZ0cGTJIb8Doy19gsVwEZ4x1vpY7
sUtEOPPMGsRzvayrlBVh3vPSHvuuBc/8sAxuRe/i8ToL8/AV7IdoWzQPK06EeBByd5N60i86ik6p
P1UNVAU+AdZaLMswgaq6IlFRQisAjEjbugoYIMp3bkhn4druZFIDZw05YlmWDLrCn0eU519W48tn
lI22aOhfGA1eap5yrfGa9AfVM7GwxQvCaJfaTOtMYlq+G7qdTi+U2SWItmUonLfvw2LUZ0CT0bNr
S0eKZ7N8qo3BhR2vOwxe5VL7whQPj14QMYJN2LBGo1hBCZdttUe2xqtnnbgk/ttAIuPBNUULpiiv
ugekhDjZrho87DnFp+kDfnxH72Vyi/mEFMTTsdfLdEnqH/eSpt80V4QAvq+0RdhpTxdgzVWKnibq
JHYhl0lXHCTPElm0J9bGjG0MVu5b2rPPtKxmxncR6aW5qyvrZmN/5oZO+Bk03l4QjwRMJRttNWWJ
EltS6fwR2mK1gcztStzij8WWxqv8QmDNAqqbSDJCNWXnWdIjRISa4dgsNFdZYW7rf8+2LepTKMIE
5/uJ3XEcQCMJ73irysOV4VjHPBahwLHqjL4Vdw++6KC1q6fj0Sufv/kOV+ZKaPgYUFhXM3U0c8t9
v8XYodOA+kf/616eEJUXznoa1b148YJLmB510hXbNmQj1eHEDSkskhX78K4QVY2Mg7RnphIS0YGb
SXidesah242VH+xCF328gmhZHYS5x+tM7GZU9RqwdoMNaKWt/rnClX3TVWu0xgtLXY631BE49lac
xBlsnlGZTjiSZMtA30b5a0Hb+LFfcBaZR+kZMjiI/ltSceACmAVKPxjbgzfhvwxPgtPmnldj7AQW
As8j+w8J7mnNAfOkVahPAQTvzUyO9cwslQbbN/Yod4605GlGnlGF3hUqJITXHyLkdTpsx/z+nB0w
g00oWnYxRoIDM2GgYp1JxVbHlWeTYuHUB4pG4WNTJyW0qKSO7pXjTHdFzIzPmkgLMvsXmZ5ctRvd
mZDC2dACfaENCFQWYn6tSV+94wbiCV/KKq9s0czYL/3jRTNkvMa7IQi6CeApX0mGILlMav7f0u/W
0Dz5ZXZjbLkWSzsB50XxhtK/YoZcEfzAogPtOWtSHxyBUvA9U4OgOUJgkrt7MyrpcG6fNHnDBAW9
35HvGVQ5+zG1cqUyK96/iAtAHOPi6jcfw60bQGNfqUb28iUil6AgpCwEhC0sCIrCsOOryg4Wz+Cd
OWrZ+2OJpVobaL032O+M0HDKNhoy5Gnv5C+mY2b0IdIHe7JMngXiWUNyk29blx9zUny14m0mkCtu
4GHtlCSGlRl/sZiPy7A0lJuLKe+PaAE1xk1TQl7OlEsZuq+Avf+Vl9CRX0B2k1acfXmJZ926xSfr
e5fgFCmwcGSKNuX30xC/ATTQIWtqjrgKxNRJy3IODP5yX112hXhd+z2esj87Q/zoAB5dNnZaSbw0
+tkqdzwU+HwCInvjLOCmU3b6e6WbphkQFZi4Bh0+sUC70e2nmbuIoSHjVqryfhR6z78k7hqe4tVu
F3m1YuRHgfoA2ULqM4gUnXtywXDTwNcjPmV3MGnK0J/x4p/fcfypFViHx3JDlhuo3Oq/1nsurw63
JBBP7rU2MpQmggNOO85cCsWIgtc3+5f35gyR74Z76sKvr9MVvPzPHJ+I6QL+7GHrRf3FC5SU1pJ/
buFrOjcl86k4FO7u3k+ubj2Nm3qp59vepW6pF+aO2QXAN6QG4RY1QDHY1m83LG3bnO+V06QY2ZAE
ghP1Y5UppslccqDKNMb7TV+U+eqAOzA4gqSJsyAK3VaBy7GiJs+IqqOuoaQNkP7Yi08W74F2mBJe
nFHJZZ1avGCeINZFrrBoyXqMtRUFAbQm+PFR3gVBo5/OZzsU72II204lsmj4AdvslGylkJB1Y4zT
p7aSN61QCR12/zdDzyiOTeocOT5DxzlTOGNfz3Xu8VT4fqgCNp170FYrHgmAWsiQ5qDy4gXXLaYY
xP+F+hKQlZ13/8xsqfPS2He9oX5Ue6XYUZBcBfRU3jur/Pc6T9G/Z1YVrtS3vSTzHBIsnUTNR1qO
1E1evzkB1Cf4TIC2rEkKXPOBaN90r0JiWx6PeG5JNc3dErYI83Nveq/bQ/SyMWJOrHdhfjt8QHmK
T1DoHq1WRwhkXz7MFrlRbNfiDVtBeWPr1G21FrXGU1/GK3xsFZF9HI944oTzP6dbofX1IngEnHRi
nSqSBNuRNXeDADfvxxA/V37Vl01zNBrw4fcptxXQd4fyx93TsjrKmg4uFIjU0k8//DRdbP4eu0HV
uGm+e9VckI+XXQB+tvspYj9PPd1O7I25qscF0uCrPISqbbivjWjZM84vzY89ySMYMnMqZhDxdzJY
3Qn2FpzVSlnQjkNTVqm822Yf8ZwpRo0Oi0X5PD+/kB3/39/e55Tn5HaEy0GSjBfXxR1K96cCef2W
1UUXpqn3Zlf8EnCI5cGqv0don6rMlvyANB2/Mvn9pyzYvkC3Guj5G6u00U0G6g1g7XkECL5HgDy+
sA/Ech4ac+xPNvTKkhbHI3DXNuUQkUpJyGy0ujvAbC6yaRzPVCRo+d9J6M8b4o/r7GEAKpUQuQF8
PE2aKqiyniGqe/IwyMcJpfxjU7qXiyfQFYSQjfdGKHKPF+erzZuiG7Q0hpr1w4KvPYogHAuJ9pBW
dq/bf6hlaJE+J3zARk1wfIsL4+rBQSuHMhT3CcvhgR2pYJjiZadobJVsObBB/LzmCl8Ss61IlNAF
ss7nw7o+2rGB6caNwRwsSdzG4asFWQQVYkf//9MgUqTon7yQYjhWYSaeQ1+tsSyQgvsIi9QAcmJx
crYTBPyhbHqCbYp3vbMuB95NaizWn3rOFNBNUse8U+2A6e05ip+UnI+vLNGurHQtZgtodViGi1FI
7FuPaPw9U8gaco00PiuE36TMC2ledK4Z0MkuiIT/l0sVEH8Thwt9CTBwv+3spJerr6qVvLddXboI
uXYl+0a2/Xu3dPeCwjBH/7QZT2MUdDxzxSBZ8UTM6ypXiO3ni6kCcxSZLRmJ9YCqP1kGgg3VFcXU
hQOnOJytvZAK1TvztQzRw4CJx9X6ycsaWBJQxsPxmS5ATsuTsau5AwSxY1CAXfBCQI1XMi7KqGr0
ppMGNXRRcyQ8tW9Im1JBIVV5kj4lCMCAZZGC8Rn+q2JllQ762MFoh1WjyMJq0pHCgePTLNlZChJP
6ATxynlemqcfXbvo48qdwf9mqKF+oteoVFvP0eveW1YAn47vKLeZrvPV00mAc2f3AW0OrdyG/ew4
eqL3EKiU79tT+rtZfWfOcptvwFKFTXauAc6vqARgOlw8KpXNIRxHicGMGXCntHtc/rje8D3pp9Pw
AiqqM6XadJY0yhyE1Lrl7FndQ21PHWA+qrB6m+uGcaNGGxg6rD3/FMlIkCZ3gaHiaKgQTxgvOYYR
zxKLHB1ArBxyAms/YqzCOeQ5VoqTCjq6/5Spy+/bubvuLIto4ABhOVrJZRVJaUAssB1XkeFGWyZ9
UPvvPBiWRowrztJhpawtobyTx7ucFX20KTU+lxM4cJI/HNYqsSrl/0p+NyPh6mM/oWaxVzkDu6v9
zl9saFV0TtyPG3IQR3u6MG9ku593a3n5HRmMIMnwX+OlrLCnOrVKovH9s/r9PIPhIY5Jul1CK8Vi
WCFuihJngXSaV/+4YWpQBIA45UqHZSxKA6rWo5h8HNjo0yJyXU6JYcRd+vuE2X7M6Nwdagpu1fqf
Dq0modNEivngaVjo4PP4hhib3YdYQbcOw1TMsKkgQAOelOx/axOFuUw6d6mDUKvGPTCd7Epjl7Dy
AECsUDWd2yQ/APdX6BqAyj3q6vzTq//BrbmNuusa8TNwwr7c149zNIr70bD0FpHcfWS9yaq2/OJM
bpYyXfjz3qz+redfq9lhXE/EGHi+c24cI2TBzBl2DicWambsrJvPjzVrRAQMr9WHXGWrtDcslvaQ
rkcW2xmxQQJD3dwcMTebWbj7Y3l2qlDHTRYnjdjJABI6TbsiFwmmWOLuaE0e3r6xVippBT4Natqz
CqdPywybfGeZILgnEsc5hsE8TAC1yQ/jFjpP9lzJDKbSctySIQu6MsulE0RVBpUOytL5PV/UtmWi
MW/JDRKluhJqHHQzYA4YSGYVE0u4YHSD8s3QnAaIcVF8EbY4XdCveh9e/mX9gvzbID6d0wQH6xfp
QNFbSb5KPh6xeIPP5jtHISi2USJw8bSkm5JNqGk4hM9YyOjB5Uvfvab9netbhcVrlA05JXP8hjKJ
bSuHzm0C8hjry6kYwtF7fuSDipF7GwAaZVPXpDJWyjVjimixmZoMPUmDkOYBmYhhp3pHbIrEvg88
Irym7kBYSpRweZkX0sxx/0dyBOQeIjorl9/raPnkOnHVEkHdJ89ElPHxxQbmRrevs9yEqJ8ry6AJ
ow6AOqSIwn1DiecqtnBQwqLrEW6kbX1EKtXXB2za9A33QaCCZzi+BNAW/p00fsiDdrhUnDDXPQik
df8FgLYOTMQU51ugp0ydHclDNUoR0HyRuuchC4uzpiqZr3FNRg7QLz98si0/0ld5UaGA6fXGQ7XD
+c6sPLS44o3x6vAUNfP4UA2TIhHF+BoTKTGZSvElB771Ok47wMxwS9mgveNymCwLFPOzi2l4dMAg
+MpnsFROckwK5OQojRjkKPw/blz7bZ5AbOAoDZ6R0Z/l7FrP33ePW8K5ft3LsAPaLB9lPAvsISy6
nMXzpwNGsdNxclLRZC8VGUr8yAFMgfAukycimFLe3WYarvPTnKwHtg7gcINheSMVgXMBM6s9ZUqH
2WicymxdWzDB738kIiXBlzb87wNH66ujjxDrGcIaFmtEz+FhNwl9GCmlEtqptjK7FSVJeq8z4gzH
pHHtqRFZldKlNeI549205E/FCOpuxp9QGiGx/UuxYn1Naz14BR34syu8W4Yk+ob1G/ZJkMuGkuH7
iABbB6evy1QQbsjvEvELAVg5GjZTJcVS+mndk5d8j9y/jRN0GIvME+iQI7+OMGcobFSl8QlJE1KZ
VixyKVwl+vAOt35TlEFSC9WzXjB4dRkbqcqJgU65t6Huiub5pTyp2O6B6xmNjwQ7bnJhHJx5+7Dk
tHbp6M9cdyAeP9aW/dTM2vRtAOUq0MqM1BkAq9Xl7vVejO8dp6JLK+VOSiRHquPLFFOv8/660v/P
Ch3f9UEHbqm3eJ0x9fj/hSZnGat+AF0bKVX/JWjZWz/XstIy950jon9XLTt+GqkuGjBfkbL9nrc6
MoIf//YMRUG0jrXL0tvdiLEzMeXt5T5OAGu5nMcLFt32eQzAHqNkTHr8i3LUsm1NwUu5JWpneg66
nj1FCxkTnp1s/UcaxINSkZyDFoHlo/FuAG1DWs8AGrYQj/Kpp9l1a7C31r+e+sAunXkSnheWCTKQ
I19/v0le2TietYvoHbqknzBH2hibyVDCKdyzKsqVbulRfHh3CNb8UVDA0eRwuPpLg/4RafSTPZlg
wCsjTfH9ikhaqxhq5188D0gbUNaYnENFJdE2p2NhwpWuazfnlCck4EVgm1PlCAaY/Jp7a2JrkAG7
b6N5q/T8ytHYUsSWB3YhsVVuWVI1KrrjADjNSpdvL4prC75mCf8FA4zgk7JjvYYYYj82vHkyQ7R0
HMeuyPX83B8qwlhLBLvXudvxVXccpvE7rul7oJYb1xHxJU8u5QhmI2RPJ9w02yyirapJxGshf+Aw
549bxqT7vhi6jIQNmtq8LseQRYZnQlpGMUMtxx8Q0JAlLhnBz7e++HUtwSI9nbOaBxfXBdscC504
aX3Wk7fmKTijvhde0i/7V4LNvXrUgKWNKvFI6k6M5Z84bmyC7HFJqvEcL8B19eZbAKq6f5bCyRh7
wF4xjJyliZYi75xiIQHbjd/9jWRvbNnmWp4IumQlBJgvGRQUS9iSVnolOmm2LvqgJCt3v2Rz1gDT
+SugeDhsbheqw3yKYBWPkHenWT4HVbbzRPHFb1CWSZ53fPtk8P4LrLoKWbru0pnIW5AiLrr8GzmE
dI6VUwv7Khv9OPbxPsyuO4EblL+BfJeHOQzDoL/MoD7DaCa+jAVYTdgNHwxzgNVM9jOt8JqiYXjF
u1KsRAcWwzE6UKTnbGKQJ7pcEmsuwYQ7CizZnaoZmFkutRRIzVgIouwDnEUF00sBwvgTxMuYCers
SWv7WAch4ILBw3e55vv90x1UhsVjWIP+RyzhCAT/DiSDfDIRYG25j4d34r/zHxmSv8oGfjE47RGc
F3jYY4o3PjirybaiUZgmkPIvI3QpTcIGWGPr85qdibFWbm/5rJCNpd6hwisd6M3CFg6rmlcxf32B
8ZLj3+VRmlSVhAXg3j3Kj19pu1LjcfwxuDS2yDUoSu3uRaNjJPFPmxBIQJC3fKWwriAQ4TNhGG8X
0o79eezt9zGRAefVUC3MRlQ6mgEOGhilcbKpvS54rNgXzbOf21UR/n+qfw3iUdUQAQf1nC1eZSxc
yXv6G/IOqBHSElI1FAWPU/vpIBrOEiqv62BoQnsqj32rO1R1ojEygBD0iHksXX/ljlPB29Zsnviv
D+nTsTZhb4rZFnx/sr5nf+LcRQ2IGdm+nJ0NJ6PJJUCC1r5NoevIjzwgepP48dvp/o2v3fc2NKKU
NYGEBT6+zYoLc/H/W1fdRHC7nVSzjR6y3LnQS8IMcFJJZoIeL9KumRovFWhS0Hs8O8x88D1NofSO
+8AnnEX+9ZEW5Nw9w7IjPEybUwWXbEIsZsQ9UE8VE8VGYuivtGMO8IiaAUyLiyfHgwL35Y1IODhE
aOy6y7AV7QOmlqthicYJuheVeBtDOClsbDnm8OATdyG/XawHPZfScyM2xV8mAdJF7axgQRZCmNin
iwFc9gnJmj4e9VQwJ1rN0FodOAm12qOTMBUBsSW1i7hYxqbM1kPv3mSAOBrvqChno1+yLE/RSgOm
+QzjMC2VAG+YF6tvQc6y0x4kKbb0GUJ5GVRTx0q5zSgBv56Q2uQGaZvXX1MnYojENgdLX9fNjG9Q
fkaSoLDcMKPBKj8PFuacTGflaApIaDhyctIq4elgx1I2riUUMz191/iYAqn3C5BLQae6cZLe8exh
k8GLY0F2s7543XLg9JqohoJQBNtdcRNWqHc0L0qURJvQpKUFlusQwz9Mwp/WWW77DDE207pefu5o
nMpD1AKQHthiiTFkzwQtJuUD68vPa0BDRaIcqKeruYEpDESX6s1UpBo+sVgSh064B6wHbZQ1NWIc
o7Y3g5VHEpzJAVOST0EEsco9KY4jxl2Zb0muYjlZzQNdHkT2gAJP61K9VV3S772jvA+aymyJiDWw
oz2XGHW9U10bEmXygMy57P/4XvyTcO9ufPNRNcu9Jg+fRgQmdflGw5IzV9R+ABGtznNRAwWY1mKB
7WcagGDGO9tRxEvJA2/f/7D6HISZ2/QGuCl9QSmlRn+V+PCRfMrwHVI3eeeaMYZixYOR1+kQf8JG
VLfvmah/rOCnsDZPiLWv3kIvNnI9Os9GwHG+7Fg/fKqlx7d5zKhm9R0SsU3ZEd3+0vzannE69K+D
Q/MmmWkJYIl9B4uzh8BbYR1dSUKHaUXu77Wl/OIY8INz3BU9g4Br0rv+zfYlE8hGDTyrh/7UadzT
op4Qu/nRqbH09j0R2grzvK1e694Y6xlDGaFNzqRQ7R4jUOXEiEY5i1Hd23r/+c6kgI1fBn7EKs8h
Itrpx7zfoYeynhzb5EjY7tY6ORrmP98l8tXqNiuoDvqoZvosCT4hBHTdEy5cE7UKnM5nF2H7YGy1
3b7UNCaJQjN6y+MwjpjhJRv11TpntlEuVbZwlBJzodcZC57uBaGSJRw9Ns3Ksap1K5a8MPd7C6PZ
gnfE2ncVM5YhjkVgjPyE2Fc6TkWP8b3D6+FOqEW1qRDUTGnzvfF9hHbgsCQiyV1wGKbDbJo1N4PQ
c+Psy6lXh+sV5oIRTrsXH6aeL68NUmsrG8kv8crc85EMqdj6qSI5oArA7Au7UMSit+IOxesKmfAO
DwxkSlp704LsLqGVZvkhkIZ01915Ro6yMU6omZ6q51qaI22ZWJHJBIoaQ0kKsd7UJvACLi2FXDXt
J3ZcfyRMjoXv5KNIZhPsW95rlGsj4DZPj7IsQLQt6+3fVw5ljYvbhjrph7QCoC0yXCmb380ANXpw
ehVWtVHg8cPbklffXgXtNbBwjmSKZBoUK2/9iIAQSjrjY6MsitPo5/cOejvozWuloPsHD/kwJFfz
n0GM5zABmup7lZDmPWMVTpOKepY68eRr7RFKrV+v9uXx1UkvpFjvrjgmpMswhNoLKDF8gU/Ro9tV
z/dw0VgmK4TiSX6Bdw/SYTeKWLDeQD+GSiyoukmqSGjDWLqCdbXKES/26pXui4KPNGoUYDVkMXbA
Tqk4zydauoCazS2n06EU+cRW7/JI0mBiQ8Blq0NdbywmknSETChGv8GdVceqj6Fy01ET3O3IQYHu
ppzQMmJXaahqwkakWF4vY280pGv8oIwDI8ISlIP2ZLq8XZmZDJx2NejK3zALUdTCSTsVrZ8Pk0zp
899hQfzKGiVpsS6SQypnbd8Ux2l6fQh4USFxZylLMRiPIbkBiYEXoNpdCStjUQPKeqVqtPVg48yZ
op1TtueQJdwYttIiy0yAGFowlxoC2X3sE+6tm/UwUwEoUpczCjpAsW3wEC9vQKA5t31C85V0M2/X
+rY6sNkVUZlMxTvcKUJZ4aRe0urIxte8jAKuACC8MBhqW44lSrfdOXk4yY72ehqjjn/Kd4mvRkCr
Nip4Px0LOiwC67lOUSljAbPMz4jSODpzcTmgrAiIcF7jhNMHWGJxSCY+QArkL7JYDtdNSW+3ecSO
NsAYf9RZXAm3GLougAmhw1lTWlOqXXESNv6mK8koJopEmsgMS7fSv5OJLv9tz0NcE8t5hf6hogxP
uw22MOyB+wh61kCpbgxn2li2YGTieBVbJrV6KvSF8AmybHA7Ph+3zJQ0FMR6hOTZuRdcB5h4EI0L
AGQBPHSrKe/paTdgPKrWfdY4kVya9DqDmc8cAjDkQ2cZjmO9Vhri0QuvbALXrSLq6QC9lzZPvqhv
YcFFfWN8HV2n1lvO64Hc8Zjopwd6RSeDEpUxZKEufGEfbvFc2iVqgGxRqA4V0Lw+o96qTlrbogkm
3PZwDwLhqdG0+067kmDw5iHt5I3vxfTPfovq0qYWR/qq91BpvUGt8i0Lq/ZO5wEUNQdT83Q/NPiy
vFcE3FA7gMv4PQR96506SqlF9PMeZOmIvxfdgJJHzdWlhCQKS6eyoEz97/EKrm86eQIBKJm6JAQ+
lBOUh1ua67HOs8Pxz1xewe5Ht1KYmlHolSM5HC90BcLoZeEHZabV+sOgFt3DJBYmg7n7bnMvES3R
5cJxJOf/1mMijuweyfR9k9zV1SRZYtOyt/kBFW+v/wgRTLoYNw/C+sCpgGxXxDEg3S06cq4ikHsq
RYdeNi9jeMECbTJzDywV3Ir36U9suduVPKAn1K91pUaOx5dlrFIQcxC+og1sKIyNKMgFopau5V8L
moKYxVcXt6zpu9UJzjDdZnL7e4zd0cIloGX/hNy5naRWp52atxNKH4YuTq6z1yO2M5SnzNUz6/N2
pByv/Y+zMNWZV2kYl364A9Z1ULcLp6ZjB7+tgPSa4kh2ueKVT0imgwZ/X9gMVyqLPlIhcWq0ul5N
LJfubeX7JIYi32tkJDGAutqgniHSBH/6VqE5xXsfpP4LepxPfEzylM++0WX8MfPbCKZlUpRvyjoX
husgyCt/uNptQ8A0+zYczkha7q9PmpYRbUcyynEnwEoiI+C7YF73pNsnpsvpJ0/VRek+9OY6B/Bv
/SScJtT2RinAwmRtJRVQABfrbo5QHxIeKUtn6LvF+/AixUTK6xH+66BNJ3hXtaS0RFmJ9vKWKk8Y
EUStOvNIbEcYnrc5AJMX+2GGres1C0wkn2JkqzT0gweukYtdgJXj1hOVGoHeUK49lvxfNdyq38yd
foqZ/EYC6O+9oLAAUccpx6Zy17r3sbxWM3ajNIAu4P6W6pwg0/9BV1mEVsfyrU/mPf88S9OvZGhD
zDEUjhwj322EguXaBVSxJIU47n171ZhHZAzDz7yTbgweepgRHfZJiAPTOsaEZjWyFmrQBtLOZY4z
a0lU14IQS/1tIsF5K3GrWrNylr2giNLznlVzoYPetUdhFQyATmRzf2E78vKJ2jjO1dSH/JvvWiZ+
3IjoY4eZpGqTdGbejCGTyfntpenokomuG1ekD95dTBWt9UCmcSejv59szv+Mq4zVRECvSB7mvWW+
heKyokKtPh4N4xJnI+sTXgwmHoHpZcuZlT5YaCgBHJB7r/uUR5lmMroI3T4pPUevjjzCL9bllooZ
wZu0+UscHHYmIbh7iLbO1QhnWcWYGQCXcXSlRbdX+BAADvQmgbbeU/DgxpMjfKOK4n5Ptb520VVJ
BJTEXttic91y194zRyzJWmlsB4Lew9YPkMMQPnjAPfgIUq9Um8UwT37ezeYZIR8rwsoo8bv5grvV
2WIqnKXl0j1ZgrGJ+62lMdLKIgWIty/LMVETfHG2XD7kFy/DDFZO55gDvh1VHJtBqVwGWGEoNAIB
Me1XaWsAtY50srozF8hV6aRrQJMz4L1MDxTIxti1qF7B1J8nIa63pS1YGxYMUyQ+r0bK0QDwJ8Jh
9Fu+Z9IGpp4t2ul8I5wijEVlGqnyz7FqIeKTeN0Z5SVGqM3GW6bVESCs/RH+lWg2ab/FdpQwHuZL
1cwCn+Z/fcm3x4cA7JLuPRnaZf4ESu2mVZ2Hy/ZvKRPz7zqsE2FDkt3DAPhle7eN5IojDVDqiiFG
GbmbuIywa41R44vHQ5szx4eP/0CVCw26Kjz+q1HLKAY122e4++0Y/GYm16In+bASJmHmoEsI7vZ7
ZSlMEuMXVoJYzkbaYApwoPlZuRm5Q18A3hD1+GGngVqT3ZIZEq8+Kjjlu8xqBfLPzZulMwnnxHO/
cgTY9dBQIIcFUkOgp/eBicTsmi+8ggj6S2XRktUSnfB7txy1c1WHdidn8Nu3rYRhABfG4MzSfUZV
OGFNABynPNudEfLibG9zMYNaTCKxOWt7gAt3fYW/8flFDaPONXsYWZzxOhNPxx/72IMCPBoa9Z0S
xZAI+TCYKn3Rp7R7c272fnp6HnDGGbJ0sLLOxDATf7CUfNDA7Oqf3Tl7+9o1II7p5//dCH4d73Vr
/KzNVcEk/CNXTatwQHl9b4VaHj3vmanFTWTC1IfDOaRol9XXZQmGk1tSReaCVP57mTnieG9X82H7
f3EhPokKSeJfsaNqqLi/EUMKw0Mbh02mrYBeR1z8aTPk6/n1ukAAOMDxMG1gmavEI2j9ErGKczDy
s6S4QhCsfcrt1NhUV1N6gb2jE1SYc3xfy4IKLDwjqofSSfksfEj1mGct9CAJ9DsXLyqwUvNo2EvJ
Y5AW7L8U8LQW2iHDHitU7cJHyv9I4rPJSikFtndTp2qM+2bDkqIH91nyIDmS5Z+1TtblZY30CqAY
TTGVCPAJ3A6XSvfwLtmNStb7I7wIdEss+MpJpEAvHFhInvaY1LvODKx3ZncAg0Gkgj0+hiUT2wXF
b++B8QhUoTN7FFqB6lpet+vDZ1GUiHUngoe/BZtwXt9h2g127mAo3iXNPHg4xFEhl6DLcogqDRTX
LtKXZADV8HDdifJ1YtXWlt+BLZKSSm38LcpzV2L0Wj3P4nRQ91nhZPAJtYuGFszKkMWBsOB8PJLC
8/UDWR/Vml/i/q1zDqgj3pLXi6crUSeWMRbwxhbbJ41egcoaIPLyTfNPw/QzrmFaNwE5mFiWpgyv
sRQcz1N9/ELYfmfV/V7FX4lpYyQrwrQULzUvJDTmW1YE360/7nGao51NmbZd+Vce2zVPkle4WLm7
ytSXbz8Tfr/TxLzRDJLKVGvUEr7b6BdxixXH60R5ho6oC47mxORCOwmkLSgaEt1PWL38Z+13pXnr
5I/ZrLgmlvREJUP3VZ2q36ADH9NZxZheh5WqKptyoIOG8jRMG2rl7YKYxIdAnLwvdC6mqapSEGsT
u0L2PM2ZhIQBFNubnxDt/aE95Ih437AzwSm/bClWPPGFJa5udqq5Lvd9/x1OTe5AvFb/FbBKIE1K
SqqJq0jFV6faUCzT1FUFq6Eu2aGZt69RgbPERglGXznv+0bgwbpuTZLACsfvJo7pnfTLvza3EkMb
sQg6XCfVJYcUOvufN4pd0yAT4wOuvrLJgE3utn9U2WEaEKj1ihOk8qytrMpB4Xbryohyziiy9GcX
ER+umAkUyAJ6zlJoTR/4sxhoWUBa10UDj1f5eNgzV4qTpxqTokVyXDVn19NVwjMGuj30C5pfNrJB
FJWuUTDIxz04+tr12oe7Iz0lOk6yorfBewGMR8K99muH0gap87BbRFzs/QiQSMVSvYgOUH6+szKo
mkBypP4UA8FubmmIXP1E/FLbiI11Rby2NizKdoaZxLlgECfmdClSSm2SL39Ffa68dv/+01vRBPn+
Ox2s0mqG7EcCzX8lLE5d3q1+Mr3Jq+r+Ey/b6GvV1mrhPb0uTs7AuBG3ro/Jp5r9uyhTdnr81Skp
cOjqldwGWW/6FCI1NN9l6uZZtsoVFeBNHL1mzLnsnk4K6jHiRpEDvPcTRfFzFUwTwZOIBLdlXkcZ
RLSaiT7Ocv5Ku0Vm1IqtiJ0rMUKI9ungoUpNMApl6eF72nWebn/lwGnrYqUipmIJARk/D+sYJHWg
M+Jej7mpPt/gdu6wHE8nf3wBq7eiD81J8ZdtNIFhdyE7mr+wnjKkMYxsx6lxcLcHIxmImfEzlAsI
WjjTFHMbNGm1PUVDK6VCFLNjCro/+Mpms8cGXwXNSTQ/xexof0eBjzSuLWSWDg262K3zkiTSUzzW
6xpWOUZO6nki1/E2vzXGVBOlMqm7H4JUWD4ddZm4SPynbaveFGwszG5e0iiXfvxWutdzkXEhE2Mw
bq8zTt1KRXZ3BwGA857sXa571JsufSUgoMPIvSfIE7B9kInS4bwrZVufyd/SRp/o7ZRUX0B3h8Ty
u0ptNDUG4Vm+fNFTiZm0VtSEEUYZNmCrJ5oQKB1/ougYNAlqunxuN9hIFzd5owVRxifAgmXR8fmt
8Ru6cN6TRoPgf0KHE+C2C49aHJXgfDv9KmkHwZdrk2IzstxQzUcYHP6iZhIspOsLORnD9i6zl0l3
t3DX2R2vn37r6ZPt9qbYrF3AHLkNj5D/GKZN9lcm/EQz7DYRaknkhvbRZDHGaP+B4qddqhLbW36K
qioZY6J+ejpkKy8hpCk5j5d/FV4FmHvRfEZuPLKKUxeIyFRRX6s0NurH6AqOcWwIsUmfJ0geF65D
7RxE3G2kZb47slzYsA6jAOn8y3+bl/aVgpSSCcoi+ZDTZAWGkbPdYzqedHYxcfsBXdSWzTjnfMcY
wkrU7WEs9vdmIVd0lTMQdQcTWKxVNDOrdc2tBg8qFNnRfyDVXMiHlT3T52nPeKE5GgY9ycY6evs6
xciiCV5KWIUt/lYXi+kxFiqa87nWcUEpRICuG0A9h2hNtnGcibsAnJENpA7SktfVGSm7aeuUO8Z3
KTNTcQZn/ImA91kClXS0yIX7i9ARONv5EJPBThP0aDBNs1wj/6qLGGXjpjZcqeFSQTqZJfWb0KH1
luxwtX4PRTxr9nYFoWIXJNrsA6p0vQdrH+6CG/tZMkXR6yweDbMaKy/Jfu0r6jXKw1EpAtl2GUXc
Hb8e9hWN+vwobFN+nYu2/F8AkdCcp1SV+PFKm+9JeE8ac2EhS1pq8Q2aiZ/UoMrf7NgmQBtYbb6V
TFX5hhi+Erad3wM2lA8X7bAG8cbVQU4FltOWfZVQlPyxzsP+VcsZntItIBse1PFkd3x/gJbTIlL3
wnQ6G3Qm7zN7QfZif/tLcX8oebGPlitY2EmcycSYpNkfrRDIy/ye2Sh71bNC5U18PizD5+W08C9o
RPD5eXV4hCI3vB657jdP43R93Pm2XxlIpKs1X9k//aBFz7L1aCmf8fuc2jOGad3AVL5E0t5wMNxc
WNpxGqsR0/HpbXpOkNwVoOpktGSp4BSGBNmDOJghzVqEsI6dxcPFWDw21t2iitKmj09Rh3imYqtR
pNIZpO5gJ+yc94mSgX3VZ7aZZbBzT6HtMmPU0H04hME1nSUX90iVUjprg556NRqKe9Bx9Gqn1t/R
6VuiXiVujzIClzU+v9P6+cmclZfp9NtJpryFRRnUnLy/jeCWG0dAsxmtEb/bT/1IE9uak9y47geJ
Wr5gSjaGHGmLvDKmibxHBKyPZ7qizyohWM6pl8LMluUifwnnJDvHayUXgJ7JFPgiWAfgzv65TYnP
gpQFH/9Rav7nMehU/4TvNTs4p+Pzsp82OH3DVk22p9IBrarHf7dwUeO/4et2A3C6ne3jWO51an2L
ThGt8JTWCFAi4N8WI8aEjXOBecjs7+sZyZBfryvNlfB6NYct41N1IN1vy67ePfNUpMKkZiXGcR63
grMwC94U3uqMx/Z7NpoM5bgmU8JP1j6WbXQYQaGNBFZ2KyEKRJtKm9NlfmSkC7KXx/axPuRBqMko
SkM4MgPka+TKhMSB65+BOFuYrHkAn2Lpqv7v7ret54TESuw9SXZMiokpWf5bozLqWcOG+UhsacKa
TYPyqpld2C3COrDK1gVsA2eg0x9nEMhgoWkg3DMwGGhwzQNMUR1b9Boqc+NUvlwI1m+66MWkaVFe
gTHg0Mf+SvtMOo2WTgOiUp6miw9NeeaNlsqnUcr81h0/MbPyRI+naBiDtQvnB5dbgzoY/di2bd+m
X9XevBW1WAMCR3k9SKT959gpTw3xHTLFWroCFzoaREl2GUR5SGv65mDIfPo1bZsN847NeQwUG42b
hk3D6C5s7KPAzL8NjFCjWI1l8Sb9JGgCJMEJSJzGrqu4BbWF8UK6wsqjttj2h2pcSOMlzOsK/sga
joKMq+o1b925DxNwOR6L5Ph/jLZ7vSUgDqaBcykbFRAvruCADG2LRsrypLFossJm7UnfDLwq/+5K
5PDGuyQeVRlCIJPBQaCSSVLOCBVlPwGJYLbHwioZMQX75qgIMPiYmnGPSpt8I1LyWDg7OSDm8YF8
Sa+iKAa97NavWYy93OjEWSvFEzbmy2L5aOkUUmyrNADXKMcmJJ/Cmd+8+97zNMLWj3DjbEUOLB9u
BwunjkX94sfrg631Bz9wFSvt9KSlMrUVMNRpZIjivbhxu8nJKfLTwuQBsEabmgyVzl7jEIjFA1IW
CyfpY6o1c1cvosrYpdD6lkib2+m31r+Hnr8zmGb3OdbXpQMLQYPF+vz7aZhEC9FhSmZYdrC/tdjZ
IghZfHBA5Le0MUhFGyF5bQ/RENzQmmMmdCv3FUh/lUJEt9T7TAm4QqlOCsP0mQwfheQLXzdmmnMm
B24gPj2GMJJD4vwmWAVgUm91Og8xaBN7MIVdFCfv6zwHuZ58ojRbzTwYlh6vZDtnl5qsWIUe5ngN
hJZ3svV73BIYFGW7JZrVaClLxoRUrOzVkOFNl+X9RuyRpnJxJKP7it+i2hXLLakiqdII9JozCb9d
Yz9E428Jhpa/HKKla5Mxia/idAxuTxRvWYjZ9E9TCt52+oGQ0FxQcVjZRLUiZKuhCaLqT6MWwHrr
PCEqlNZ2x+b/COLVO8cFn8Jl1sCbmqNqIrFfhzpEyEUNRPt6oBlOdrTsNkUqAtvsE+Z9frRorFoO
zjTIeAY8yu1fhVCQdq3jvZc42eAYLu1Pb9tkFgm2ceghr37hwftc8tC9cxGIhl9lXqQzEfwamdJW
sRScvWmFz+n3JBuAqRZtP01+CDNx2puaE6AcyjL1nBZWL9kMAu3Ab1/R9+SwPh2ElRxTNUGF8lvW
f4WVexPDQcVHl6qgGT34A911Yd1/JLbX5W4GcjcdHxT6ShsqkemTf/oxyVzR06yyTzbvOfcs304s
8lKWWoO67or1aJaAO/fGTjkV87MALVfe2XrkT5QdQUeqe/818Ouciv1nmfnaoqqTKhSgzauQISHc
tFCwhibfJ8EJdvGgnSFrO3AHtrqtF87hYSN1oV+G1OCsNs0Lci2iplbrZlffcndVmNVF+h2JDJ//
1j/Q/dhdulahz8x7BFa96VWllnzfJOHrUq9akkbByco+99FvHZblfnMIZtVcd8xwoqm/V/V31GCj
xsQVSW/NAShJMUnCyo9VwY+yVqFlp/kYqsNnI/AT8P9XH85MEkxQ2j9MJ958k2hzXWScBtYsCXni
myal6S+raRcupQUHUBsjFNrmKqiy2uhEV7fEUnpn2KZ1ue3WOI821G9A449cNgEVtLj7tQ/mytfd
brK8ke/u+Pag8ixNEC/5Yj0ZG7CR4n/H42h6wHj6GHCXKdYFZqQtOSam0hHONixGyd7uwobG1oBJ
DbHKYqbiQTcv+QT12WHJtE8mkPaIUVJhMaPluMWhVtVe/otsucvKY8kzVa/jLdWmHNJqSqcpK9Pu
y1g8VY2/pmlRpxUZNzjh+3KNooykx23iuY38j9gWLf1KkZ6qyoR1TTeUBgffGZznRqRl+fssHmer
rTm1qKbknOo6aZD8v1mHZgkHXzHHuyArbRUzYn19tuVO0rNePPnwGDddMiLm5Rs3uChjLqUR3hkN
tk8uRdH+w+KlqZBj5KP01+t0KwXfif0Stl/ALaG7E9DS6eCCSQWwUUkmnXfQj6LZ4anKExKPqciz
HHd5y1EbNax1B8qbEm7Bd4bfaK7fvX3G6M8hes+v8vdbuqG0KIIOVTaLCINoJv2pyOygXUi+fk6b
7/6ZKw5t3jHwMKdWK0R/CK8efa7LwefHCs8NI3BBKfc2IrZSkCR8ioNXB+oa+iU5bTME9EMO0YGk
ju3RwWfLjadsDzr6u8+N0o6VrXyJLKXjU1iz7LCfOESd0cssNoj9LiqSbQnqgZaZ+1xjjlQlqZqr
VT8hmA5c5N3gZ6nDZvIzoXEch1rGywgpQ4wQ/43uN31V22hS6kClCKJR68oIor+IcEzyaIfvoNih
cvnjFa5F5/mjwh3KpygecVj3PygydJ1kQhBpbeYYpC6k1SNDwIhaK9dz5UE2894cW0gbqMWwSyZQ
E7fwYfpQYhm04HQn345QGntQuTrzNCYKFqARHUweyV9SXX3c3hacfnZt0GPzBPr/KZv7/8Sx/xv0
XY6EllMRItI3/18QDLAYIiJaVcQD3AMTyECu2w3AWE/izBkV///qI0qo0CxTacNCcchGyEYvEkTK
w4mLhEvSzNLi+akfZhsnOK408qPhyhmfGkfKti3rXdnvLJu6UUUjyOlvUgy+MKCkXx2Y9KKDmfUr
KlnykX4U17eIK1RIhO20ySDh+Jfq3OT18iqPNJjofehHHVXHMoMCJ1X4YsHNKGy7Uqf+7OgRYlSf
T24ekJk5yU03erzFBOf8Lb72n6otovHbfKvUZv1Pv0+lYoGUChbVXZVnDLVoOGZdtP+lZp2DT3ey
4eclBl/ZezW69jhyC1Zbrf6qWhCSJN7Hg2vsvqj6cIGKIG2iSrVH24zPKFTKGgX3k8KgGNbpqfEj
2knh2bE4gddaKVymYkvqKb3w898xGKpUO11wp0eqhRqED3Xgur6NDewImLdpsUNE0R9gUiuRLQ+S
BbLcfx1CTFe/vPV8XjjSnROGLqM94U2OJ27KhPwAzGDbhIVzcfLSAeRm7otkWmn48L+eTyNSvfjq
al/atWgKyA9kefjD1s+fHw386/wCtB+zWLfrZ65gGc1sbCLeHMowDylMNIvAk/Qxd6GekSQFrnfj
dn2N97tpSfSnmcybrabEUPpOrgzktez5qRTvHERhsxP/Jp77pbyV1GjrnLRkqx+F/Bj4HUqCp6e7
lZ5DcoEt5bzcng4Kyp5kylOZiI+IVtxr80J2FHCXHZOsw9QRiDr0P75ZeYF7tbNfxrn6Z2oZgYD7
0KA4Y+42/aFNtiEV4LgKxlUYX48ueAyqnXiXli1nwUToBYMajbU1oB3ohKycmrh4z5sdcSNkupZ8
nr6P2XnXoR21fy35e3A7y7/9D3xRo8Mkwe8wlnrysP4u8GnBp+5vN/2Eg2J4VPGdy/HyXuglXN8n
jryWgpwBHSr74qQO6XWphSeZxnmg8Wfv/qFNsDwEu7D1/Ct+qVPRpbwGqDUKq3quQ25TPNGi1XkE
WW6Ds8H6OQcqZmQ1geIxz0AYr5GYGGMJILBn3yeRHFcEFDCfLTapwmWYfAhWygNCK7DZJIn8LivV
easSGkeGKf8dPTY+ZgJqp/U+FlRd+AAjDitHaMlNiY7o5esbaPB6Evmhn2X+fUoSCnSgfhLBE+V8
nXmethQVP18asMGRqfL2mchmeVNePJviDgg1Zcl1mtg/eLkfzK1Db6N6L2KEyKRSAiW9t5U71o/S
zkd7Z/71nMiLqmjrl8nnEYLnM6IzlD8iF/DTRT8iNBSMPb/NBZpVP8bGJOEMgVRESNQC+4ST58ZS
0kXZFRZkL3vizE0ujS6ad/qP7MoyqFSdAf6gz4XfL3ArR4j1Pd2JabsdjTOkwCRKdiFR6wuZjOH1
wYiVBbAnpqElhbXjy/p7eAud4w5WrazeQb6vjY/rQp7oTZlAHrvTUuaIZb/G2q/obbS/xYmhJ1b5
buBVADmzEDUMFJM/3RwVUGVIiJbvusyCQLJA9c7Ka6k0P9wHGZKg8dJoA2ztJB3XJv3wEveGlAU/
VSvpNc+YWWRrn992iNR+g31F6IwNE1msFcZtpC4S9lCPvxMC/396Brl7GtEIxN6/cD3BN/qjtSee
uVTMA025Qv8Tw/UvK7aK/Z0nMNzOS4/CnHOjpb2/sa/OhDPrfcsy5ffm58UGpW53BfNDZEaCdE6C
hEIAPkzQFW9FJkrf/IcDutAcM9isp4hb9I9gQCMoAAuB35aKsVAl4njj6qOXJN7lLWDV9R6MbFiM
Oyls4IM/G/6nkIHgmN/zQ/D0XWOGgOO6+uvbQx3NPVSrjSBSLqqpR6k2t3irz/9bj5XR3y3B4H+q
SD9KFPSCEH8cna7HQdJqVxLh1uXU6bu1U6N/UUqHFpBE87/NuOBN+LRAHW0P5hbxfn5B7lZmOY8S
MwNP5drzbm0oczC9+0X8UZlADVaYZPVnpuUR9SoeeQGuvPVe/qitgx2yjkP5bIwaw04V+xtU3TuE
eEom8J4A0uLY0OgIHBu1fnWJm9iAIR8liILxRXDne3tj9DPVXrAWU8Ml2SuLNoowtQzirmJCEZ+2
2QD/UK6cZe5LNDPR14Ln86KuEnNP3h6l08dvX/s++PQgC99ffrPYvTXeKNKXq8w56TjuMk+lOIWC
NxiGcXfBMZtF6LcEPp6gwd9V+E+VmLTsr6Fc2HcgkuIzgWqPAqJErV58B9Jqtc4nEx7ty06JZ5vW
CGRdnNdvlCujgLMv+6LU515wa9n0voKOLUW6vyenQN4U6Ky2HIotqFftome/7+hisVrXHczEnT9h
mrQ5j3Wc8NiKZehTMA0ii2JJFFV36VPbXzAhdyq7elcc386D4BPEje3UO6mgh4zDPlVrS4uDyByb
HUXD1pGGzaJ7sOMhc+fdEyZ9H9gNGBq32XeWOo8tm6NEpN2HsKYelhjBgQSuJGcI3u9af4NVaHkS
etfLyiiEA71mj9MooCqN2zI8Lpy+CId04J4LThvho3eFIUhlX9Cxb+gURrh2m1q8HO5+VgE4OzwD
HdlXsP06urYuQkTbwRWzvn9s4qDPVg2/ddpBmPNfZt31GFsjB+J+ylcM34k5K7JCsTuNsOHpyix7
UGt6XqK8/h3BqsTiTnaZaTt7OiEM6sGiEgjO0M3+8NttE/VaO3xmKCcqFJZT8JoAzagbn2HAgRjc
t1AH7JyomTvgbRNkPohOMSPhM6VBUKnk3i3ucvYQnf6m5ekdOGRb6NiFDV2LcgSKu/ujuj/3MNWq
IbU5XFwbBZropH3ljJZh9Sb+Z9AtsdKdYZAlSTGKjyKyinreH8AUxP540RbMYYrF2fsIT2HdKcbA
Kpq98+670OMHUzK6doW9ir5o/cHg3Klit9qTRLEF0zkXUlsHpLVHAEsMvw227WZ0kMgRkEjJYVOX
D+2CmmyA3DllgIMZno9fOqzsBIxw1sf6Lskxeg9ZrbJbPnDcc+harLjYeVEGGPIZVtDXRFHViJwW
WcnSJbfA2UL1e351CqkFJMngFQ3EE4VlFj0sLkdrQT6aEUAkFaJB2fBx6egkqOFLMEfGdsp47lU9
b3rmPNBqqUS2pEE09RARZcg84dbJApFBCCUkE+oodvcWlRNwypCMt3B8uC20SsnTP0fWuaudKHL2
3QQNJIiZ34CvZeNBny0qxZT0unDyrmrmi7uZNJWJvDbQWLxNQyhS3pCWFp4r49Tf/hTsTmlGcatt
NpvEtYGfqWsoLWv7Z+Y45Bu/A9FCVg0d36HDFPvQ2mHaST+YctROO38UCtCzUls00rqaogcVO0dy
/snN/nq8W/SRameTu0kYssH0Dg1QUOyBF9ZUN/KFuWwyBN8FQGEQG+3UbSc71TpwuiqFm5QLVux/
wxkBJDKUSegobaPIPLQ25Z59iuSU5/tSR790o1evbEobhP8nDuSZstizEeE6fS2lVwaqkSozDij1
y5Q0UWJOch3XsThujmWaNfU+94mQEtYSVf2e9XJyaoeJFY7EzJddDL5CNOFoGa4+7t74Uo4vJ/WZ
EmGaDXM96l5p/uFcBxGeuLdZ5QVlwflZGy2WkJ+VBWdUinMUSdz7zFmLivmbDFPmevXFU4/YlHZp
0eJLgWJabc3TiZhIVSNYnfuTLA1Mz+YAIBluwMYuHO6xZag1Lj/Ih2fUoVCXdhD6G5DMPeGvmSeg
voKsYmIFu49RLt7w3YHgZlrcziLV/ypnQ1v0B+V0fSX5EkBR65kQINrmEt3ZgD7swO+Aldvcu2Hq
fpbfNm5MgK8nKCLQQKv8EVv9UJL2PjHRyVw6ZUMU5Ll/DHYXcV09j1wYQzeayN+6nWqjiLABoMk5
O74JNlB75hPU6pvhet5hMZ39XoNMjVkl+G0YSDsiRqKfV37JkaW5+f591X0X/0kSH/UIXSBT5K+8
C6ofBslnG/NLXc/BFuqFm8jGVgK8l64+XTFqSfdZ2vASX5kOq+myB58RU32A9GYAYMl2FcNlsAsd
2QCxsjynaFj4WIfrz5G8k8+XM60afTsgb+KA8shv/yyaCfA1SmESDWHO0IQJ8IePxysR4ZaquPrL
YF2Drxpk2aGDf/AV2AZpAoxl+hCSxlW/kfkj1H7aHpNRhkGYdejUSLoo2qq2wUjFYLY+Z57MvqwB
R8//DCv4YW+9Sl9gfBnMusD59Z22yFNyAMbciCcuh2ge2wMjpF6XTY2nIgpiuqlfEuFznunauubp
YuctMJJNGX7LmHrMgrnPe1tSC0VOAjilavN0/FZLe9GtXQH2T8mnhzkfmz+5rIEpyIHGSes5Tsdg
5BWRYbzkIgWQ7iBP/vSBomAN88NMAVosiGrY+N8AWMEiaBKa4lAqG5Bheh0xxFMEoFyhCtHlUSQr
fIzfIus8j+O9GrsECbopAmaKSeDeq5tsZLM1uVaGrZ+FM5WZxZnCeiuSOOVWJsXJK6FE2sAH/V83
/yoZhnim/rUvGOVc/nd9PwlIa5RlVL+SwzwWkL8elQXFx2tYZbfO+7/pgOWmY9PnVMl330GmvQdh
7xGgKqBe6M6eN6jVU6QPdx6TkwINIYPuUO2rxQi/PcTR7dQyCCDSX5lMTcg+8HsovSz4P6fHZSFg
KFwY9sm+9C4GMDEINnhbDdVROBIrpHzfraTdobcI9b4QDt380DKl+zrULnAjKj2uRRidbtr8QSKO
tQqwHSeARmDOcLHKqFuvc0iTZN2Xv0g/9cLBpbtGEdua8Lg2j92toRWnbvB40pucf7nMKLXekRRw
5iVCBXkeFzX6MzaG0lW4Jn1HBmn+cV3UD+wqE73U8E3C5LlPYuV74EI+83FqwcD+bDz1TfUqt5ea
IE3jSqQcf46FQYCiAwQwU/hVGX7mIGN6F2KTnKRI5CAZHaxWE58t0iVqAZo/0DmuvE97NITISF2s
++HOkcWaOw9Q5Gi2a0UwG/Vm7TILNXJRX2qxhPqDeCc0sfUXzXnoSn0j1/JmxhNi52R7DxzDax5G
nu+GepLueTsdOvf6Vm/9DAu98gwt+BdX/hmzz/8s6m+Mq34k3etOkFVgQqpXfD7Zq4/VS04iXdKU
T9HE28EeiDl37qkvZvqOFIKEXi311TjcXy4AqBFBVDlPlhvHO0wsManXyClttipLNUi65+8wj8KQ
k5inOUYs0yP2TqaYNS+c0l5D1sKyKXwPhwsk9hzYL+GMcRtrqTB/torkY1jeNkRHBz780iZSmbiW
wfnwprQB2bp5IAictOD+mvYlEip7f6VWMONoDV4+FGXRxAd17ehqDUqKtPX371k0gDVwH4j7q7sS
4WYdnOECUbV2ItWOVSKTRJdyLJcWTrONMBAR9/VAeXIADP56J22o3ARchXIOnbXxgIgvkEHpz32z
ekvgbVrP+U5jnZcaxwR6kvkY5VNUygfbqnKZw/XzWgYIu3PpIgrgX3kAYcXUp52NMec2Jz5RcKtl
RnoKAi7LBzbqkmu4OBVHeW4JiYBbdO2xxR22bi+Xf5ZJLRHceStuZE8iKSpvrocH7WKShj2h3IKZ
WQ8K3IEVNhTway6B8TP8L5KjGbSF4Wc5Ya7ouLtJM6O7EBk8bvahmiCXo2ZIBjQBM4iO41XVFT1i
3uu1omxbZc0fw5BhFJGNtvFzin7G8R7DVnyBitpuBicbK/6tzTkZO1DKMUoEYuMwdj6qrxycm+iV
TJhVA3ne4D5zmPRfLPGeUhaMFUAuG5Up8Kp39WXTlY9X5h0Ls40yulr2Th3igUboaqOKtJdnS37b
0gLRfHb3H3mJHBTLTfNSQl+cuQ0IWldVsshwOptdXQG7oAXyMF3Q+q+t28TKY1htU6Cw3ZyAbzse
eXBdrUtHlOR7amsGH8Rtu8G/QC+NsEn07Hju31tGf3nbHM2jAqxcMOAZ1QY186PAZ9QMsp16lwR4
QbSbTX58P1o98tBLpJqJz2GuIKvrNqLI9Dya/kf16sGNmaPgcqTLhJbSLe+cfl7WSyzILJnrJO55
xTcoo5Ty1pkuizH/3Gk+3rQvNrg3WQ66guWvM+YsF/fNa/VDh88oDWE2YI3NZzXKXD59eKxxpbqH
MnALXiNyyqiZW3zCVQR6g1GUkFJvwUlpmc18nIi5tJ1llUPgYUI3T8rEX1ndbPYmV1jBhhLVUyHJ
T4dSoEXzcESvtHcebjevB8X9wpJpk5okgbXXXJeRNPUd8WMX5GZ1yTc9lSO4Am3vnaU9rnWIANJn
IpbqThXrI1MwpnOOrNZCdG93rFL2whLfvUrFU/dPgtjhn/yNV5NOjvYVIBqFi4BwCSGjvZpjs++N
whvSQs6DzHc8W2OE2HF23Rt2C5u6mFFP1XgBXDo9CyoSbYrFVPT7n4xztZqTzhRgqLn2xEE33m/O
LI+e0XELRl0E/WwHW2+lv5SvC03WBx4Y4XlDxux/+4apbQGNnKtAR6jzUlV8VwtzlcoQUqGeemSC
gCUpEKOjxntW3l2jIUOgm7PdC8d2lkoWxMwdz8odwB1yjKHYZxMkFuTPJdvNL/cWwfxigY7+iCbW
Z9iyg3H7HvBilhDLTjEesDqLbq/rFwYXwW7USzJ5u3uJsvKoWteTYNRK+CCsOua8BbLywjPTwo0t
yLp3ow+UohR7E215InGjHSHkTj2IIIo88ILZPSOLIB/YgujZQy1A7yvGvdZDAnXVi5/4KEKFcf5v
V/FVz9AtvOf5EpSFy72SmYsZeMCZGwoatAodtuU4swp3VrYsaDmVEyJcDKN7B8zJiCKT+AEi6P67
Sj6RTQLKGwgGph1Fca3UfTTewsmBBYQ5UArQahuLZku0KOs0E0vGMsn05wZs7ZQtTLHQcr7ZrPIJ
uzwimg7PYAe1OlzMHGHMM9KJBrM9cA2S6yLaA5lfgUjGhK8SFWvgsxMKK8agC8LgqMMuzYTV2Ky4
mHqdCBhJJSGpm4SZJjdtG9bHw/lwiYj0720zErSMNZ7JIia29Q74Ax9C+5EG43i2ZO2utNts0WAG
wjDDcokHtGD/inCZCkKcwh/if1+QpsORf/LCGITywq4pNVYoSfGRAwEnuDsWojPE0mzYH0qCpgFw
+gjl1uA2SEGibKHKSQtXmmIm9Zjridzd2KA0DUZ/ZfkdvZvRpxrTSIcW9IGgnwuoXHNkl+LLRjCY
msyCGLd+mW21S3QU4Ge0tYX8KBOkyqklm/PiIMNa+4OIUwdHUZOyLGrlHYbcEqnndXyGbJ9j/jqc
kI7clJGkc4hNGkMtrNl7cDsG42sek+/2QclrdQVJEqZy0aNcQGmL6oO/SXHuM7TAgN0KNaEzzwFM
0yt17G0S1M3VKzRXkhPiwTOiZYYKn1vN0XcYugJWk8l7adM+4tlnpyH0cO4YlT4JelEY9ZfeW1Y3
2BC2tSTP4XPwMXkTbQMhp2bztsP1ICEPkPIrCZeK/byGtZP/tzqHYxki0REldFEsIum4leCaX9EN
ib8vcRfR6gKj5iuEMHiJxqWZkqUyaLWI00GDm+53IwrYHEnCrvUQU+Mn3rv1AwcYqYMd6apDe5z5
0xYet1cuB5VseGpYkUmmSZx4eSAw1DFzFx6E5MSXruVXwAgJyPBXWRD08zTtEOPQQ2H5MXvwftAD
DwLkC3iQixyJRJ62pADEMRt54k9jQ631RcNfNtDN2GWFe11Q02r2AXc5U1VaROcMGOUcVJhC3tIb
AmcC6haSJr1MgzNXDRLT+7szXSXh88fe2dMh0pVfNvcJUlJB6ocFQ7hrqy+rXqb8S6CzUtZ25Pz2
P6d9t2cf0fsCf1E4d6Huas4EUi5/UNnfo+i36kicZfT0H4gJHxw5R5EgguKdPheUcWv75CnJhHDu
GXIw02Zj9awMaJYOWW5qGxXQBq+MeiV6o6bJslsp/GInVw0y1rn5CX1DLBfxcHK9Ff330dFSuyry
o222lzg6IVcvb3Zq0RnQUgbkrVHDVtMcLCMxmmyYgUDjX3aNX93daty8iZpXgPjuQ5GZov2HcHB9
p/5I8zwXw/Mq60KdOfy0x1lcDwrV5Yfw41VEWZ6iCbfCNZC1FBlpkzUL7aINeVAe0qJCnyFifYPq
IAUy8tU22Qe1ZIoFlLaKtrB6CiXjWfvjWfAcs/o01o8EjEUQdANIEDJmZVSvM2EwwAUpAiiyLBBb
0PLfrrCcA1R4uszUfI4NxZr1vJp7B2IorgE91ienLihPrKyt4CyZgsDirrN74KRFU2AEQzYCO8I9
gGwo2FhdFz7wyLcLMTcaPCiNMZwmf8q8l/4gTMuMGi0q8TvQExDhAEOTYPfebI76YsPbKNV9Dv9W
p4+6qAIqRaVh1b0q9cvUzhlb+ITNIvOIlLkBq7SA7+R1fj71Gtv/QSHaEbHJ3vjTkrgbe5mfadta
VpD46jTu/GEQyDdjjsE1Xd9kUeKq//5qtlwZdSUOuYewmWuodRuJbGr1cFyrCM1GW6nY2GF/9CKk
shWiQVOuCe9cPG1EKupKX0C5HgJdOM+xe1OEhr0kkmFF6NArDHc2T3U0ytfA1qTVPl4s0BSxqzi7
ze2tw5jv2bP3woKaX4DH132hBST766rBJn21CGixq0ijlUE20L+6CHd9sIsig9iPkt7j4fIp6vFd
TnW7k0ATDQeF6q+1RAOKPwXuHG1nySCVrShe0hjXD7IvY5Gv7lEtBttDMm7ZV8aeJMtjtJ0Bu5Vh
bY+Y+9verjgib+t4kaZ1cIEcH7rUGfnoV6h12wi18Ot57iQGo1LUIPSUE6UgTPDnrqAitGTStRZS
6U8TQ5f1WCciZEkRYd6JckZq1bWq2+PkqzrETogFdIDTJUlqrYACXjouQQX34CtV2F2SEwBKXhyb
hbOKSx9kVdoe923TwCdvCU+CwF3AD+yf6CXnUE8exMSu1vQpWug/W8DDOPlr0nqZR1HKjDqAPAdp
hKgLAsxKO1QtS0ldN4C9lvgJn6BZXfPHNzaRdl/62ztRDyzLutATrSnrM8et8YbS86GzkCCzkYN8
5xn0GHbSwDa5fjeaTQeM6wSiw8k6jpxrT8NkylKJz/nz5cvyEZIpg2pnM9M3XWwcqXbZ+QphhlLw
WBN9zZsZqGtrlF+323tJnRyAWgE3nIxs2s5snk/mj7KiPeDzy82b9PrUav7Jpa5Qf7843AO89qzM
0YvLmIb3HLnr8ws+YW1OLeYIl1L6kj2Z2qm1uAFYMnlfh95dRa8HTuYMOoZCzUuA0eBo8y0bXXm6
+vu0FNpwElVwEPr5pgpUBvOlu85cvJnGJaBQH1Hib58ff0CiTn9LPzS0wLQNgKRh8d0ASDpuBYyo
pH4U6qrYbshvU/c03AGWZ58RWCwsLYHWpy7m55c4Uw6U882mjM8AM2Vx+XkbjUrhguclrw1WIAos
B4EMMcLOVjco+Zm38ILJDqlHrcmMuKiAPLysflamvGr2o+6SnDDIXAFRVAbgYFgv5O/APyZf6Eqj
IoIPdZn0Tq2esft2jJ9zBdgccIvtf6YCe1DUR/oMdCghbX5Du01Slizy11NyOqgAOzWcHoG7X/C3
hzZOH8cA7LS3YumioFtj+CU6fDJmjiYCeLcAWsUyimmGsYBqMtGVU14FmVCbU+MIslgDGEWr8dgk
le0U6OWEI7yJ/EKO9tNu2rX1bKK4xIwGQYaqrYkdVYjIf4YxBuLfCw/3D9ufC5PdFdO8Eww+lnS2
kqf6z/2Di2z/4nVgggpHKP88io5Pto/mNwZz2ijVigWDKcWy8PG7OxU7VPeD7FWcwkTqy4R/RhPm
3EU7zO28fLbKe7DHA58IZUNHgouyvEobYTkzgRIO14jdMFkrdu6sYwGAZFN9ZklsJtsthNd5D3eJ
6nORE4fd6zVSq252JgW8d5qbDds3LHHbU1B7CcD9MSVUdyyfddYqjCkH6r26p7pYs1AXoH1mIoD6
8x1KVX9wOkktQqwO49nuXUhdq68muEHk60t4uqUe26f1mo2ddsVz0Ysk+vQ3U+nI9WfI8AM2VYSu
lmujj3qV1Q4El2xtvtLM5ueI17mZ0B7o0trNMxYVhfz3PcRFgWGBKNcOn0NIo/vd6Mes1QTQuSIN
gBXFzey5z+3b+RSTSmmzOUpWkoCMVYbOqyBvLYVHlL7xVOtV+oD4CPN2wwv+noL7zTykd0vwS/yi
L7IdWcurIuAeqNCx/a2qczlzUYD5Udoh/pLdhB/BN9GTN8qy1wK0Aa0a0g3C6npv/4QwT0EpxZQC
TPqTrNBrMPX9HknyNJxAqFRcd74cGka1EEYl4xIOA678PvDp13BSVAP5VXMBYE8xyYtJmC+dNR1g
jXn+4ac1J8GqqFDAoJQKsU4JTdl4ItEpP6zceKfjTI5P/jOOskLh7U5wtlSoSmnuEpuGeGcS8AD4
D3LjGfyWOIX84huy8W/iXAViGjkyJmuElEpkBH5gs9sBRL6IC3q6Uf1JSA+hk4GHr4pfR4717MLi
953wnMw1+E+jI/c5qDMRs4g1WtqCh86X8ZgIDw4NL2bgePmZh0MSpHUrTpREwApGz90GMAzS8RVq
HUkXodvy2PcD6FHivjBz7r2pwEA1c3MbiMLv8QMzMfjhVKtJD60UXf0gNw+bAKbomzZ2kDCNdMgW
evw5PpGxlbocLL5IvXWp/H93Is8A0A3s9oFUB6kWACXN2SlUe7VYSs/UECfL7vCTRAmzWIpzuOZS
GoasF41Mrqmfmmt+LzGF6CdhPTglJCPRK5MMmmSXDXtroPSuxU5Q5urZwKjgymHjSXh8CZuZFsd2
+5MOkpEmy8fRvSVlO7hTMj/hSYRtygOeKWgd/tBR97f0aahsKu7ElqykATAgZ1mHSVAf38ThGsrB
x9RsCM3grmokFOfjOIDqEFGe8yHRi2Pe2JL40o0UlKS1O/ROSM/nhLih5ukH/4qsjL3Neetvo8Vo
MGEK75qldR1nmRKfl3ZtW9dBHoDMOO8CBAqjHISIiurxMLqqDArEU94oFG4Mu6yJ240fFQfh4aV1
rzaQhiJfLihj3jDmNqZyxYRt61MUmiR2fEW+AJv9jlNZIRLkrB6UGgUEcZoP37hawStFP5ldk4sl
LXDo6byFovwRRf1zBPA3xDKMyAcRbdQYp5CVqCnJ9T/mcXEj925KEWLbMq/ruNGGXAva457X88W3
BHdIFPKlEWTvn2soKtPZsEIkTI3wmzIt3QsI4tgdDRuP2KIuTR7zH4RGxRilNZubhmcOIbtr91Sv
PUtPGH7G7fnaWm/NExwB9dvDimAr1J3hUS+DJGIx9PfjYRR2YywJ8RJrvV8iFl18m2OKKFwnJ6vD
gyvgbBwu3qkTQ++xs0dbaC9kBCU+SoZnHDGYMpT3tP7WJIdxT82lCtNSsRh3FfCoPWOlKk8xbmew
sVAOhwZYWKJmwreHkUMzsQP1rdMLJd0yFs5yEBXUIShwE9ypMalGq/t+oHKR24BB7cGGwlGGMICj
ZCsbKX5/uTnDP7ZBBpl4HuXt9uU+hEKy+Ccfi4nn3dvZkZfShNshGUZ5j44udBrLs4F9XrAjCGYh
MojJI3uJih8MHRRzJJPHq3YF1LkEh5MGkgmFgikwBhKHvPzE/UNFkinwL4X3E388C8dCMoG7cgMu
KejsDI+NU5qbggcE1D2I/FXBKldBTVGqF0jrZkWG6wAcyQUE/r32xyJXHNTOtB2AJY0QfqAtvYPH
yfGSW7k4nBUjTxxxpGAMBfCaMR+1PZJhSOLAX4wypVNqDS+C2p37PA1b6LtHrxgy3xgL7/5+664l
gvz89fsdW1FFtLwByeKxNPGcZ2RRXWqwe7WEhOmFwptEG4SGbwOPZe3vqvM5L6tFue9oBcpAYDc/
Ja0nw+3Il+mNzD0IxnIqX56PnqM01X9Ss6bt7Pwc/gPlGW35wcx/1SSpGE1Myp2+O4YyR6iFVB1n
+86Eof+z8cy8aH0ZJ2q8EdgWLBYc8HFI0YBXqk930n6Y+rMfw51ItlRI4M70etogsDOlqM3E/hKL
7AP1pW6Th5kxa39sXWqVbMwMR9tvLnFrBrPPiPZ2NlUlcK64oRdh/7lkly81WlztAQVd6/NZ2b/W
ujHEUvu3OmJjuRgYlRDx2+SEVivmnZh5i3AqQ2NhO/uAIllW+R7hEDIpqPTK0bZ8l4VWtscA+3Nt
uBtpTpUnJ/S6+rHraazwnWdrIE2ZpLg/F47UiTH1SQuriWLbVP5+n41tHgUJu+O6s1Q8d4vDe4kd
eN4NrnEiTkZvnRJq5XPZQytf2huOIbhoi++dd7BfZy/o7MN+pwCtmwZU+sIgaN9Kx2mONoJA07pQ
qZEGb2TNuefOQ4P8YNDLgxyO6lASD/YBhpsVKaCRTDscI2AJqoF9EH2gDxbmnglRmb3POBAR3DWk
Fukp8qH2w6ksHOfkbSy333oGhanS7OFrXVhr7M34HUx6wLC7qE35iQdNSs1+Bqm7wmgW8vB2f1Ss
QCl0xqeWO8saUZf2aoZWqt5RYKVr1BjaKdI/24f5Fzb0+dXNnpvkcQOu4TOgsnVmXVLIAIJsWw4c
2eDu+OJ3nzv4qruo8W7yKfDrbA1caMJQD1/+zRo4f6BzKeF3/YEhVP0ezgxKBgeF/cw2NmNsTSts
fY+vGe+m6XpwPmyTKPWa5jJTj2U5dJrSk2tD3mGO+hJV9GWUjUOZTozQgkZc56cTf7l/FtELDHfc
d2jVpHCsz4Xeljvd/2kby4sqKul1nPCFL1DGwrgRiS11aKxyEWJExegp02xJNmbF1n8w9GhEJdrU
B34gySZGSryxQCOxRJ5OTKyetTnsxZ+gJ/e1I+Z4+xjm39/ttOUlsTjhSkTQWpOoVcU6bNEGBrVx
YASxLRw+7B9jpFdJCs+zeatZ1Z+Nm4W9YNTXLNyup0DXz5SBNy5sGKvxYapMGDxp9QX2ceBcPdws
wHSd6SRxvBOIMgFOKT7pa2MkSfHhxE1z5IIR4p+X3nu1MyyIPWvU1+AE0eE4rgiJTnFJcvUNm06i
9jTp50UH3yKN5J9VBxPpMyMdgwGAHZnKtwpq562pj/VA099jjb61LnfSix/GuTz39SNz5PCTUJXP
UCJbN6oBYpzm18AZfcl6o/BNRz2fLnH30l0qNhQ6YExrHHsAW/SXbd68OYSQnt5LnsM+OAzVDyj5
HtTPlRaIQpn2Z/qzK0IGsrBMUWBuU56atzenXNB1hYY73pPUOzVDDKu2ldYtoMe3C/87tp4WYMLl
7bX57nqZJysnEOtOcxfl0rVYfMl3vewd8IX8OHS/gcWyGrn1VUz/huKWd2e9Tw0D43NiK+H9lfwb
+g1MEUNkHEIimL3GX++ET0VMyognW7wn49UFY3A0F8miCowEOPBEWg3t9qLR61CVm/93nIcSKb9p
gTX+sjQJPNU5nyqJotT9gjynbyVAT03eGYK2eemrcaXZZSjDitqkQGF6aTUfhmL0jc8yaTVDa3Q8
BfeEqonORBbXFcwd0jBsD1ikX7D123sbHf2YFLIx1MIAmCIsZVhojw0krYpgzZ+BbpEsqvH/w4uZ
9tkSJTmO6uhTfp0gCbdeyaFbg1jbcbumYLF5FCMyJwPguBqZ8fo2vsZxkTYUuYvqxredhw3XmzfN
iAQ4IoiRk6qJqEag/qqYcrjdj9J9fKz7wb9eAbklMRZ5+4Ov3VoYZOpcNMX6MEXDGThLMhwtGFwA
fPdt7yoMNF/vhX7Di9TVIW1CWH1xSsWRYYY3uOuo78lIl23RX5xZWBAotMy2LraH03ELKwXC92+6
WF6eDYp7DYF86Y3NLItrcQ/jHeQuXSJ2dPW+8vQmg/lVfURhbBgnPil99Yj8R8hsKnbFegGVr0ei
cM7FqeKwHkTmACGuOVfvOj5/zPjHVfHeSfgyXd6z+oFS/+RFBWf3/GhJx1yRk0CgUifQEODyqPOi
oTiklNvW8xN76Z3rBIC4AkIvRZDOW2DeAuW0dTpg+JpIbJfyE9MqboBxvIR/WG9O+CnHo5zVDL9y
rMr5WSRHHMNRmdikORxZ2ZSJYji+7mTbk59W0moTLOgb1vZ8gqsBkiWLa8gZHJVjMGjwyer5HsmU
rNKclshTnzdOo3T4BHbvte4M6i3Vwf40WN3E1T/VX6wlfEVeZ799rxYuH0KBVGoAaaENZDpQTOvI
Im2XPdb8iMHcfnkPm4PDOQhjnDIlyprvt+jNDoZqVCD4mtHpOLDO+eDT2GeJtYS5aLDIxl4THRH0
Tw9cojfGBd1h32l3JB2IDeld8W0aKbFt5qCGktkvRrSjdBqKouilOldXRX3uPxEp1Q5UHXrgPvF4
jU1MZTXt5NiJPS6tu/QWrfxj6YqRxCy2h8LiW0qohO668ykHgozmfOBSWiKxYl6QiUFCil0+BSxf
v13HwqWVhn1AHXug3Ep0P96FxkDNTva7yDVy0qIg+DokH4oIcMh+pNqLGUf6EhwNt+mzHBa5UznA
kIQWVZRZO9bWZslNyiNGZr2a9tdgPJVlM7o/3pZctQZKUCXL2TPGkmUSkAI8mXGPdC0RLxFloWqw
REgHHinWlESVAtqDJDW+sEefEVd66i4uQLa0e3d5nSUt4M2WGoIouoF1sQvXT8EKTTz/Y2iMpxal
WqJPp2GidqBySUdNYQD3tytxVLXhILuMwUg1bZWPIf831HKmSYDORZ0YCYDThNO6uoRH9nKrzO9g
2CXEhayXK45sXS06UOXwuV8p1bnsYDVULqNPj/yV61KPfv2Yde24L+3Npt+JCfTPjZn2lVVOcmrU
1ZQ9pV+DALcl21/Mfu7th+0CljuWJJ+5BKEVawYvZWoOObRfHiTxyBdtMBV/EZpBEVSX21HMSkEl
iw+CrrCNlERUSEMKXEpjR2BsVz96+4tgqbVYzvG/VUmpm+C+Qc7ALGMpFr5V4l8SeT/tm1c48arm
jT8JsDYmEVlYzS5PUXAPzNtDGT69XnyzrhMErIfKzMQ3WhBwPwGZuH1iE/8QtTtXOpCir2e4LXYo
cXpJReclBY/xB50PHnXD7zTl6e4I1PAHzo+z5DYFhMiIQKF8qrEfHmFMVWPA4IgWtDJD6ty14x1n
7nNNxgpfHUg01OFojmFDzAYA3C2mWQIky1o2hKC9DJ15najLP9kBULFzFHRaTY+T9qq8H2RRa5Ww
1XKNolaNfbORIfbDVNHet3IEU9nKFo39S7L/AZWaINnUyV9poMEe7ArFzvXUKhovy3dT4lvSTDa/
1+7wM973CI7i0k2BMDPQZmDI26Vm8KVZrrCddf+tHzhjuQKhyFRu72kpCfipHHGZh/aqirN4V+73
BC4EdFYTLnLLJGYuR6vVESMjIKCTkcJYFhAI5APyC1+cNSRl/08gRjzsofipl5lABfhx2zYOmnPk
CaInegkVlXBa9sh88Yq8xRO9hix+ReMA65yllYet4P7rV4PO/KuQal4InEaaqttc0yZWxG91tj78
EF6rMVlA3r8ireRek/Ef82J6d2f3rLWUKp+upu1KTtJvAn5VjATneP3Kgy7LAceoHZ/bh7gOpZKe
+rpyWcCz8Y59VsSzG8QOCTlFKhGZkHEkrk6pHertXCSRYxjGLO3szzyxSzkdujDwJF41g9GNbl+j
HTgIbtEM/QLsW/SjEit7WKmaXjpcu07MGuhlfFTTUNC4LRzb+SyyUFaDHGRHduYGmeQyZX+8YFzA
eedcl9Na/NY6aGVvXi8zjwTY+p8vn12zVH4AeoK9LaL+VJNZdg1h5hMbQqQpzH3yG/SbzOXj/z8i
dRmlBHlhzR7C0ZBqtKEr5CY/ByEWI94f+naYb5qid5nxRgrSXkFN3NeIX4RGVXuaEQrW9Makp7dp
PUv24x8ntXlBv3+k2ZDDGvLY5x69fpuySiO+qXbYSfFoQSUZ++K9MFqA3GezmOuGXunhaRap//Zp
vieYaEkSyz+93AZ4mJiI2sxCtqwng3xgMKhGllujcH3Q9AyJuRZFZDD8WcqDpQ/WahMGxEMhHQha
FCUQk8/w7akBRwnz+T/wqPpF4Wj1AzsEr+PQ2LESDeGzwDBk50xM4s0L1GUEabvsJNdt4Wd4/3MT
pm1GBDYAuxUh5rtLy2VNHu8KSY2Ipuj0dDSE+kvrNoz07jeLeuvHCdDUMvpnNsWO/niGLuPFPmlV
Xfiyt0S2IKQgm1YggfCrgDl+1cpVogj6qPwEtUf8K8wLFpMf0iALsoKJLqILDuiIVC+YCX15K7V9
Luqx1IggQ/2ToDBF41rKQrJZ0ilZ6ac8bMHFNFSygj2jX+gBKoA5Hyturb0stiMWNlLmB2umpVAS
6R7aWbcUuScT9UVEo7F2GMc5tSMrUU9qOuhU/DPGgBHgkHPNnHKctkooKqJrJQbiHxLq8BBqBh9R
K0ozdqv2+LRuENB0dkdr/LBSFiuqPdFuk4UHnMfTlD6UpdM5UlTdL3jkAXTq17RaHiNaIClcdkk3
aS94x1yKK/hyy1WvX6MPw8i0eAEnlezrKLUo3+G6fqpCWhvl+o1Jt2MMhDkJt8q5rP4/zFldIrmk
RHAwknHbi8InldTrMrSA1AYPazFcuz9JdH2giiBMmosLv3AMnqtwDR94bYY5ARVwlAVMsVslXtoR
wm62NhWciBKUXYU1BEWR4n/ZJ04iyq6QOcKCtDRO82gC4NtMXm0kQvK5Z/+AX3Xzd2URtzY4MQBx
mGIMEGwTrFayCj6JuQRQ/ozqihSc+oJlVYSf0JDWuLPM9+o8W88BDj5Py+pzTZNw750gZ45RMBud
4MHmSh/fv7MV7ZCmqk+PT1htY6U1wOc6f5dm7JhDVmRtQ6ABdZ3WkCxAUh8VvgzNFk+b/1hl2ypJ
aDs/fCuTFx7E8pZWttnN08O1YKHTli7K96c/lNj1XwIc/zRiOlItSgG88fEAXoyXmrE7usA+7wPH
hmPzAHvUP9oA3e/HaZSeyFvWiYNm7WqElUi8m/7CrwZcxgx+knZJutL1VMz78h0OluBQNdV1Cx0Z
Ou+V1FKmJfH32icJWBpmxDTzXkEgj80ktWifDFnf3qb0Xi3juZaORK6x1rb1rx09Yck9A0us1ZMV
XdF4hDWa1y5SJK14qVeaTmwBmFywJ0yQkTORg7WyboYCsfqThkJKElZ2V4U44Z8FqJFofsbtAEGj
sKIxLNnVQwPatHrKdJ9wLKWx3eFaBtzQllJtElLtpLKh4HzRtT8r6uIMQlp8nqcSmJ85XMkICjeh
kqlenlk6ZZax5Sg34lLc/+M+lTrqimhmlzzeOvfkkIpwf6mHy/nMgmBtxvVkbLyT5FDukei/97fa
O9f7bUItHpOauK8K3VP3Tc5hdR8wyZ7x96Kcg/szeOdMoyj7cI2DRJM4n39QGULeWBOtjRqdOELl
MEy2XGBNBfS9uvEyGpJT7NeRinfcGYRbvFTZRzppOnSxCNcjZz780Ofp64PJm9tJwJMY8DVkOINZ
MIjRcu6C+V7q71wExDZ8Upv1RBC1BWInGwm3wLogp5yeVsmMFNKfeMIt+5zEg7/in2eG47LCb0U1
MPtaQr3h7+zx98zDLWK3v90dnCRLE5MvQ80kzlLoS2w9YSLEHSUcsX3nZGGO9K6lwht+zmm+3k95
YSv4YWG0Tt+fvAE3iehaN2joEd1GAMWkLsVM19hV+BENkNHtKy0VPq55Uw7h2S1li02YuOUyPVnM
1Mxpn9rqpYWsrBf06SRCv47epVLTX5eyNzYi8wfWmAbYkV2hbFty/fBnwZJ5C2FEIxQzAw03OkM0
+DKTqb2uZrsiAYVpVKOWmXTvlubjvzXM4iy7W178onLx9T/26x/PQ0pCzeF4qCp4JdsoOXXn4xBh
6vAZjF9JdGndwfRlUf2NnAK9KAsTJGdkEYrKQfsI8ILGIKl5C6frrn6I2Bm8Mgkqgxo3tSXk4gZc
UF7J8arsGUWhvcvfzVTQ9dDSwggd0hgt8zImtbbGBYCowSKfU2awG3dSOQJomnpM8BkCPnXxilqM
eaJF5dC6wWi3ut0i/nLqO8zsGfaSKb8yrP9kGmrEEM6zBUsJJ+UHkNKqiRaap4KPFqqeWpRh0QJc
UBNREk1jB0u6NF9vwzh3Ve3BSxwUMj0WFtxG+8nDu4wsRgkDt5GpbvnoBy/MtxpxLeENlu0ecNXA
Lm5xLHvPG+UZoZQeEy2OXnHjeD0flpHnARL/6E3i7glUAgAI0mKPS64d/jepeJ9YaOv4bTvgkz5x
fQez0QyGfuvC5YN+BnHBnVD3RoTZzk6y24mfWuf1LCL+FXiEdI1T03eTLardud9Wg/APJkzv4r9f
Iw+fi8m8AyUBEeGOry3BmT23OKS+k9n7DpVxglnDQp9rdXmdyovyfQ6PmVTAUajTeiFrR+Kd9NhD
ma60rmud0Z3DByx5TOPSItakfXz9PnpuXZE4ahD/Qc9PqOwPZwhfoMD0d3z06asq/Is2fNuEKNyj
anryLkulegpHVIrzSog+CxDNaSMwDe+01Plv8i7sZndz8MOM40KU0bdjF1IAIbPSizLmpYRPq/iU
/rSMVw8w5H2TByri7x2o797WLIgc6/oxQAGn7Xs/biJJnw8SV6pHH+bp/2qwusvqB/4SSLHPuZGo
jsCXiEVUddDKyH8JMZj/y+a3xk9D8W/tp80F3ydnqpbtKQfIm3GfgSyfxQcCGRpAExAKE6Q+sXic
ABxxej63sicN+0BVsPVLbuMXOBz4w8gqhXQiiUwtnVcaIOb3QOzjQvRpXcEkcVbsTcpsLmuMoMcQ
VvAZ0YR4GBcMw2SPtBJqEEU0PA6+Arphar7at6c3nVIzg5O03CUoaCblwHOASiyeRSjLKm9lQBio
R4xw4X8xYnW96gssEtITS+LAtR/YyFMqCJMeo7jiDXr3xHK3hkM3ng5Y4UrqyC23vE43uRUsbK3P
FBE8Uid7/YKLb1bIlay7dZi5qemFO1CLGeQSmd3u8ch25dWRrj+gM/Nq1FIejuutDRCySYVLb5Yl
GvZzE2jYL+d3zMcA+eTOqyQL81Vv+1DtGd/oDtZQ+kEWwl6zeLNU0BhhkQRz06TCNWspGpGcKmpr
+pFxk9WXTkX5cf8Xu28Hzn0iIZEDzWUIxqhgTRzZl7mShibtx9JyNzH/wGm1g5cYb+CY22qgnd7z
LMJxhKMZGNjAzZMsKAJ7IzLOK2c/LqXVqCE41huVdOpe5ivzI5VDPxXURrOw5zHweXgm+HXhKc4M
hjZ6bTYcZIO3A82Np2CIp7Y5pjeEftZlIlPDZ4hWPww/VgwzOcFRdvlfDhVNnZQrc+b/Gh0Sn3Su
vNVgZLJNXbxsMiKKXlU2AH0Zj09KJwSoXBx2g/pY7W0YVcoLTJ9g7lSxlBwh8NPikPzEzztdjrFK
vEdVrrtVKfYNylM7w4IL6MZmA1RQ+8PCipcsV4hn+b0BD+rS8jffwPni1OtuyA84X/YWg+mTNpB8
tIu35EIkmZ2BZtYYB3B9FvzsEs+azkotfrFiNkvGGXfDeYWyfCzQcZUFFSrK3LFJk3ubJCIsXeAJ
cTbcRNpRrU+Z1SHwyURbgLQ865w90X8upxX5TalnnFt7HpdFecZV+hZyjRzGhPv17R8ePO2Ruo0/
WsebgVYO+sFefRd23+O3owt8BTFbBXZxh7ub5LYkuHEyve1T31VyxO2lIvXjDfu+GkUtIODyRLWu
S9p+ZKc6kChmA8in6Ua9kon3ZiDrWrYifdOin74SZ1o2P91aw0vIc6EombE6jS+NtdKRYG9i6dE1
aFzQw93Hx/vm9z6+LalIa6Q+WGJ4SR5sEu9PHP66wjLhcW6krtpXLizfzZ0tPqtNy0otORso8RNV
1BP5iUy1U1vcWy9YyIqqZga/PBaZH7tUpVJiy30Ih1IN11dIZ8Pl278pdE8kKqT0KN3IoAsBIqam
7u/XrO+lj41upxpNrOVnHEeNNZdKnQMXfbREWbOWSfcC5hL5k4CBJFiLaYDM1h/7ra/ZJ3oFzwge
IxNFPnp0740x8eTuvIKgpu1Cd/We5XZLNVhykdFDxUIInDd1IJL9BAZa5HmVp8/0ijW7UgNAjPQo
8kiY56L57Iv9vH6t8YMSEwMAxWA6NOCrYPLeOgjecnW5ljjYkV1762wVWUepCljM4Gl6YPQR3WOG
Gvj2QNJE4pbJBSE6jKoocqnaM61cdW0xcaIF7+nTWPSLzrU8aDqGb3n6qF/ZgNOCFjV8BJFUUx2A
FneO3J9zqX2azyJTsM/CXBeU7qws/FkfNHWkTZqIKswk2KoDyra9Dj58m4yHtcUpWgU2KO7+9CoK
gxqpHCuoq5Ae8csHzK31YF6yDVNQVDtdr2uX8zY4NSHBWDIE6TQ3wt1xRGmP82UFrk/megLcCO2w
6JW0wa1pDUpXQtNALaFMf/JQA9DAUuPrAqbxeCDrVWQ1brE4UAlR5b7q7Np6oVSOl/L4/bi8KGbc
S9/tYiuzQ3Upwd0TW9zelae5241g6GPU3uubEAtbcPKrmn16JB4rqJNOdt7lb+d6sB0FnOrRS9nc
/rF4NVLHBVLllro8LKICFiTbvUTHCzUvZ+VcEfa9sk7APom3dbDi1J+DNsKSG+Wk+si/27OKOzDj
rMGBRkCf3vZQc5vkvLO3ASHOmZTnDeiF6wo4q8cLoE5wwgCOlNI+Vk78g/NLDcsX+PZq59cRJFjE
AvP3KN6s1bui+7aWCU7GuxxI2nIknDtS2npp8GNfWXHJmWe6f+DD98EVAuAAl/pXOi4ICcGhEamB
tI2yAgiTOkz6A80VL/PWTHmtMoQ4A/DaK16Qu9fiIR+sJgYxbqqRc3h6ivdcCR08lM1QQNU8hzwr
ByZ+Gqhm9XHJIy8FteRyNCSSyAL++FtihBg6r+2s9/hsSGkKgJcmuHs1SuQVR/HEovpeSZGTITB2
bPAzRh6Gc70nKNWiTcvs8ZznYUY/oOv9nvjmPACVkn08VUdEieQDEGFG/WKBUAa53EFK1CvJRsq8
ivFSXiiPkwS799ncD8nmmJu9pEhhCbaI3r56niV7DBM45c0rIwSxPDsNGl/VBPlbtE7vopXVyi20
7fHeOJWNPmNQkJB6cWw0X45LeJs096x9bScdhBsbruD93guzC+m+LuGZVuRx8foLd5ABz+tZGyDA
oz5wYCbMjPIW4LSc94BgKW8aLAxqiE/tu7gjwMRoumXCy1t44RAOV6r0sJp8OG6stF0Sy6XpTCnH
nT+35Y0hEitUtvDizLYqkxckeKI8Zaeo2GFf5rp5iNX5RKv/GHQXDDeu5YXShE+wA1CgwSOWQVIu
nqaGFqsc+UoUj9dQ4/+xJ3cfNkWnXkVGqaxcOQAIaEdL9uJ/UomH13zLiT9R9PlK1k9q5uoQOfls
Un4jiDFaN7UQ2utsceIqga1UQxky2h6UyA15bUXgjdyVjkQsz1k8GDQ1elg6RkD2zmAkx5sdf9lj
sr275qXlI82CJmhAyANRoIblnbe5fIPz1FNwKGlhTw/UeGvegLTaYqoLcJUHQYWjx4qds0ZpTpyF
x188OO3hO7Cm/Gm3PEDC/Kt+LfpKsi6nXnWVawz78QdzXV/dXSskdXp4HVTZoT5hIIDoweYCM6Qs
XYKr27kCRYXrZQp+cGZHv7zwvY96+wrGl2Y6TGEXuMMILAUGvEcLQ9u8H+8pbCGM0Vr+brpsvTGI
qUwMzLlWLRv+VX5VcxMHtOJamqqjVELPBwsqNSEYuXLqBnugcT6Lvt6nQnJvnnE9JPmGc80GPGA9
GcPMHLkWYGy4FopI3NpYt/LhR625akmsgM4Wh5eONuWUmwaNjPmcQjKyCo95IqtOAudIsH9eLTBn
CzfX/ukpAp9+VaJaKi4sP036UwHnWzaIzv3+p3dGWmpTUHc2kydHGUoGUSA1gNzag0PXU4lG4VAE
FAkJV6hk3cSrVdtUWbgDXgDtBtXunDrVTK4cWVJ0VhFdQuO94I1t3fHqeejcp51pXHD0JJEXI4+z
R6Ztv+YgP5ffe4CusfwaDtYx7alscraxEW0AUnjB2sk1Ti1T/Ci5SmZydyoazd3R/1jk9g5J4YwK
9JSlawy54qNxVbC3V9k2KAToj4iagVu+TUJm8frmS6Vgt84ow5o7VX1X02kqJBWHxwdF3tHSs98r
kmHaKnxqPLwVXoQ0chE6yXmTwTjIiJQ1tPoIUtiDGVUarNMaqzQ5uO6B3+9E5ISijwjwEzb+PMQX
LHIJBNPkmavfrp59duU2uOQZvUaJ3Ukj1ToYWB/TMdgoH2l+7vN/fegQ3D3Ajbn8u8qnLJTmO/Ct
dml0b4O5nmNB4QW8xeM9HCUdkAzuTzuc+2QaYKdF7Y352Oa3QWS2MQxotJ2n+JOg+YiRbJvCrufW
dy+mOQdec89p4d1l+YvxB644TQPZxvhZaSrz+P4EExebRysph48lqzEyYWzzGTqtLrypnjM6go7G
m3CheMhBQbe2vPvCCqDTL+dVIghgsS9S+BRU3P/MsRK4wRUxD9aObksweITXZVw5ZcblzQM6+vKa
nr1ZULxnmZlDbKSabi0P8Sr5haCzGuc4Y8W17IbwrUTRzJmM+vk3jtTQE3xU4bECHfS7lBar4QRN
G/1wtgcuubmvCRLMUclJN6D9GlQIOFQDbt8lFTaVuBalghZ+DVo2weBTE1er7F7dwH/FhkI2zCbf
dqwHRu0QgFEyOwCs7oFWvlA579wneFS/E/GhRIW3m104AXV64/bhvFftBwqTaEnvGdIhz2WQQWIg
cFnz432MXXcLuDiagu0tJbQQtgfB1qk8JrB2VpdsvlaqJy3+mLd414uJ1CLrtJ+ZzGszm9KOBCUO
jLmFXEp94gaQM6uoQApPDhvHTtcmBnjltzmW9X6EBLvCjsNi1DDGovvZLFVVcQN7+TuHZPYOkwtA
vLHbBR4QTY2EXhRc793tRenufqcw/QDn8AlKyLteuYtrn8GoJjiVLzSOVSY0959IHqQkGInpAnye
jzKN34vO2rw4jKo9b7E9WRJT3r/5lLFWwqyJz0E9IaVgB3Dc1w+i8jchYjh0OTrgSWU1vWcd+u6U
AkUgU7xfskBLSH6Av5imXY8Wv6i9tAI9lebNMFtAT3udy25CgCFAa/IUeOsI9FT2tWvdhEonnCCp
nrHNklQSqSuZdxha6xHlUwx2IyLpaOCHjaS2IIukyxjTtv+mPN54o3USFuJoPiZq8w/7Qmt0bGu4
pRPrHyQrSTztqofB4Wg7stWy9u5WtQReTFzGRPTAjH3sOBheAlexY/+BYU57YovLTRvwzV3AWREo
qrxUk9jRgCYwhYdX2o21x060VxyPDmCgpqftYOLDmCA4/XyAtPdE078EHXEEe+I513kyk9fU3J6w
t13YRn8upfbKc/E9lZMAFa/irqDy2DWBKLNUEREBieFTFi9aMTjW0vFfaNM4x8TLIgANKuOWnNbR
AEyAEMaAgmfuJxlt425e2IRe/WTN8BoRehs33DDdO2WsVwN6ph7+D+h068DwgKFB6kt6P41ZDzy1
p53IID5Eptyr7PNvOfBT0AQHeAtDBFYse/sB7odISFvb7ZyZky916265AqcmvKiC6kVQ70IRug2y
bacjougTJ1q5QU8QqZDJat2YRiW+ir8hQs/uMCn5qIiFUNVBziQSDeDw1PzQqZplD4T6jk25fEnD
dMKWnmEOyo7s6A23U4ryPxmykB44nQ6tr5GKd2bqKYyITrGipMvID2biR6tiCvLXsBzVSgxpxfgu
DHH2MuRWO0j+FWRhKHY9Q7wxp9TXQ7TFaXLNva+q4FiaRx6PfAndzMlMV+/uGDqrCNEB1MUs+Z7m
13xl9L6poXFN6CBfUMsRGePV8TbfFAllAgA/UZfW0vpwIfYtdDm9vqcSSpPGxyGkP8iJqXGq0OsR
ViI4HKwS5QaF4kWGat6UGNuHBquZFy1+Ej2Pt+MNPewkqz9RM9MvNMjkZOYtq9UAtKqkDb3CSZSs
ye9Gbf2Z4qSaMnuRWRRFlQs0q3s+vNtDPMpJj3JJyYNM1qAa/jRAD8wFZjO4sazoYJj1r6Bce0fr
iDDAkx+xK7+zpPzzWhzk6+Wds7OBCspmwvkHtZUSVmDoDh1L6JnZ4mTTc+jSf1lELvJ/o/DHD6Qq
UUN+/iWSL+L/n79imCObMubgbp2eO5KT8smGgeLStP3yfkDy9jz0mi8XHfNxdD60rwMLh99V/54/
1zFNnxh/h+QhtLURcY9sbpEyukHNKRx4e4Py0WKgSGRSypi8kpdxswNhUGAHTftvFPPM2Z2p8KNm
4deC58p6pol8V2TW6I9TfT54Z/d7rWlWhdNV5OWJl/oB/cdvHSjjewzCHFq8YJeTBvNXWwfzyAbh
6SdsGqya69w+BhbvGuUdj9kE3NC6xwr2S9YmAt75f1qHwwmTY68SHAfsRwfvoqKoz71RowOk4ipP
kBttdWomA8XQ/ekSBAWCGMdVxb94ynkV3DuDuh+JfcJDD3fS9ksyaRq1r6WDVE6Z6XK1dEsHUQGq
ESHxkuYBV4Aun9TmGc0alUgFToSn/wOBiBX813XI0eC20rbtN6D16kSyl8EtYrjQrDPbcAlt45MK
NJpAZXiOV6KggSeV3FIEx3tf2l2K1jJ7uGHm6wVoQpNVId7Zg4XMrxSiFgHLM6LG5AIwFLTX4CzU
eHDcT6qg0vNr4Fr9W5FClV9qnoHPFHq4xZaLPG6VLo9P5zx1eyrpNAjEPqNj0LlmERoJk26aK1La
u76YzEEhWjzP0O5Sk53RcrR1nMvV8IWpPLm+LlTXsoxZUbC6ojxxOcYQL8efCP2Vau2nWA4lptEj
0Pn8DfV2C7hFdu/wJjrvu2Eau2ODVU8/vmBEn4aZNRJOjtCaMghCNK9bG3WhnZXNJB6AVhw6pg+P
gA/NwgH2DWMKLjFuDQ6EsQKjufEdP6l8PcsAjRDNCFPn+iWcg6CSMTQO3vVl1d1mIfaywQRiWs2D
uGaZQ6rCMcuDUAJ7D28ipk8twq+NvDnf1gw0AE0WKLU4sOge7ZwzTmVe2ugKFeOk75FHBAVwgaie
mDtnV1bA6SxzM2FsVSaminClLtPmBYp9kJX0cuvmoKGxlFO4+rsavIKIgIO2Gs2SUC14KQwUt58d
9EQL9pLXZBKiWeC4xyNPuwQRvgPcw6DJHPs5FF4rAvIbIJ7kCB6sdj7/14mkJj/Y3oC6qy6wdpKR
Wt8KSuZCUqXhSYYC/5gezsgQh+0Fc2Xjs0eXT0CA9pKe6VsD4+05wMGa9MejMjx2FauyIkB4FHMX
bp+/2tV0S4MWlNu1nYabJzJgHfxL243JRm4ZHA+URswPRpXohanQRzWUPscR4wQWrcKA/FBcYRr9
sTtnd7HtrqQZjcnPctUTXpD1WZr84AhIWKsk2k67NvuRYKW8bhhCjVHuGpOTUD/0nAZ7XRSnoJZ2
oXd6a7nFTsC3EZPkrS5PdB5S48iMt9RUU4CYy8bWHCaAR7linESEUKWKYOyiDNppo5MGwGs3DEPW
DDCKCYaVCVQUNGNoeJYHUdkckclV1posQau898UkpndmUsXtXsf3yQQ8V2z9FY2pScv6WTj57RyV
jqnbV583b9g2o/VCt2QVZNSVvg099rtgzRE2WdeeSmWXLh9rHzLArh1VoEnKGxplxTGJOcdi1qQw
yHJyB0iPKTcJVyUMkjOua6qwxPxAAGBH61s96GETHSikFVXZ0aKT5+8GOLGX15Dm8EO13Xdegc73
qyE717Mv4u5VC5hjzp/gETVoox+q3dFNwaklmunfV6tTVp3KNYm0oXZIee3tLno6lK9lYhAyyWdW
q+tdo2prY6r/4AIseTVzwt3jR4KG3IKkPrZ0i1UMAVUXc/8WGaJtzV/YT59bIu8NF7lhKGUImjXr
zfe1y2lz7YVwORVa59loZ2p1MB1+c2wilTvdmEVV4HpbgPiE3cYITRn0n+N4F/DOx/g7Jz+yIcZZ
g8SDyVWPOtMbKa9Kda9cvU+g9PFOMYjO4rVWGMuQmhA5HN/6qA9dPMvADryfay4+bs2E3i5nLilA
r64A49+gNMWrB/owfGwleVep7L3pYqv/N+StlZ4daLJPg0OCDWPlvLC9J2HC43UK/r4ZO2A2gQQd
EezyZW4tsMuXChDSycujzuL90TEKr85cdFPDdI/u6ZJL/+g7zZyawLPKwqefzCY6wTCmoBRDP6Af
78Hcbfo0MTOnGYI7CPoO+eobufZ3Xl5TkTgzGptf8fBfBtS+3j/Znq5rWjHPFezo82jMZUPLc7fe
kKJdy1soaOgrm/yy9cf9rODhYtZVSdldSj6eCmZPiCDAAFfUrxS6KylVgSXEYWhMYm93pmvTttgl
tTHKeZPArjrTdOCk26O2Y8WMViISxWbPPMKYwp6vJqoywc3+P4wK5BJEnIMpeTKXLmw6+SDGhszO
a0TkgjZCu81NALxT+elYghfyBAl9Bpc4f6S7K+8KVeiVFdhm+Dr7l0ktfkVwOLb5dbd6GT69SBUz
IO07ZDBAX/nSRTWPJWA4WkB04YqR0zSgwZH1BLi9Fh2YoaiL6MOTyA5A2tATQnrzJWuT67JXcgn8
6zZJaIwk+O7A/22sGkCuNJdoDqvyCfvnVp7acSSkNrOZszTVqkHeIvKQeLf+c+Wwnncn1AwxsC+U
w8SDNhHYZZuGO/foQZyXwIBrNVCLXI/HJUXdb5Ve+uVRtnxLu86YPkCJnqp7Wxdg9dtlL376QHFN
zqG8gWFDY5QtZAAOrZmRh2f3XpVVqcVdgHs9sbOxMXvTetI2d6nAlVtaq+3kR4MAe6+u8z+pLyeY
cwrAu1lbrvo2NQHDsFHwSHJB/4+ulEBUMm2Ea02u9YrKH7kVwm3iPD0tL6TUT340iX9TbBanrSKE
xiMomJdmF6hCI9Lw27nFphrXsHbUbO19nBLAJPHvkiBYUnT1BMuLjGE6U+/6MmmozWhPYIksK96a
C7tUc/kPuz18h/sMsPNP0e2+tHeRz/lvuohuuKmMiEnHxsfvjaeAv8cbPY3YfK4QD9xJCYfP/0kV
VS2Yy3BywYbXI4DTLwfXVju7eon396zRxC+yjs+7gLzzqk7TMXuVte4mtcZLNxb20hokdpYaCqX0
sOSbluadfnjTR3QjTVLztDKaNQVp3GH6QEn++Dz4Uz60Sz34gor/qnRTXuAdBYJ+6Bhf48tdI+Lh
DAT/raAwSqX8n3BtthkcEJcG+SnDkOyuXkrhHRHmm0aBGptUNWuw4+rpsiNH1eQn1pAZ1K6jN+xZ
z+ngouSvDkbTCY6FTi+AIC18e414H6RWrDG+SsXZzIWrWjHhzWEXLUFs1gowoujO7VacMqrYgSkq
lZRcYY+bj+rUksN9Yo2BlF8n6Z7T9gPYLZSH1j57Nb/Hx/EGv1JDcovI0vs73OMJFoCWiJ7ez9Me
7xF5N9xeJKhAPGf+dtetloPVY4KXFOE9cg9HnSzA7BcqKWCLBfEqi5P9+4Ab8GsCMQz8sSItrbp6
Pcmhq1A1LYVG1TDjr5US3NUEzdVPDrtJVH80HarzOM6Utq7q2XAcJAiMwLst/fSR7/mTyrxzQqQy
wVZT4NVZxCce7cjh+Gk6kcFlB3HN0qbX4o39rYibJ2NMmQ0I7snApTWqNLOGsMezDmPn0SS71w0n
3QDcolgtDX0qDclgUV31ywAZ64bv8FzAvZZ09c4RPGZ/Kd/U7FkSzQ9hhllS2XBUewxnL7D+paIy
WT3sglxO8giec8LMTXQezT3/M0cHwlQXY/kBNquz99hC0zewwEGxPp/pH1/bevydyFNOQ1TC+nFQ
iEKw9kDHLrGhhNB7Ox2YcaBw6Ho5RSuFYvGX4d/Ih+kQDWZb1LGv+f7c9dcgPsm0R0EYcT7RvT6K
Hv+8uvwIHLt1ACpKlVfNjjs/JGK534pQ39Wl2PBjc6BCwedi7V/Ril7Mncpdov+bs5HcQBP8oE3p
cv//V3WCDXalt0XNZ72IcLvnYz2y4hHB8+VZQvU9r23vLAXCaS+oeqkr7Ar1Y8Dafw2IeYpfxeIo
rHx+NZJ8Q38WpdCYUPE2QfiMoZ0wYiC6z00dj8zFJPMmLjTU3aF25tfd6VTOkCtGrgPr53OvsO/Q
y+UfSOvCxJMKNqJ8guDKbi3cAfb9AwHx6tiXkVSSWu5tImsN27gJKH6aV8OMkCFS1uFCYoDx7FyV
Ba3stlmaI2Xh5UyPC7mPmaEtrB1ycZ/eiCWi7GmcS4oXeHaYa7klzpcwg7d0Qqo8YhqytkIXe2xj
/LaffP3doFQchVtzTVcAR9AmYcay7Ar8s0R0tkJyRpqvbevkiy6incmAnYkMYPsnKQLs9XYSrG6H
ruz04UJwN37OxKWhnFsWppzC3yw+ByI+SUk34fLG0h7hjq1tg9JUku3X1yC/Krjmw83S4mwlX7Bw
BN7mVkBAxBF3S5BRkC8+fFgL501ZddUnbMLSRm9qRW2qijz44YvkPqbo/7fYEO0Z6uODVaXILlTB
aGadD+/0pvwV/2NMvHY8yiHEqwY9xP6h8Fl9XTGUJIGZ4xJJC/7bcwAUVqpHM94dj2oe54ZPVQpd
SZaWidW/TTempkEM1oabwMNctUVzK4YaBplmNlo2O3jOa8xpxruUNcoTTZ3Baf18+MegPF5zKRXw
r6jbC9ZHv/hCOVhWsbltJWAHfT7YxerX48XUG9uIBJaJcyaAgB0vmiKO9Nq9V5EM5R3/byv2rMsd
BLfa4kgP9ALGAs/QKF01z+7WY9e7kSbI1ZTsI+TodGGzwO+Op31rhlIcYtXZ7+R9kAcD8zlEeIwJ
tmZo2T2ZFNAvLcy4bx3P4dooANi283fZqlN8H0bI0KIhATNbBUu2c06WrT2KgXXjJABfH784joXr
DWKJqseEgd+n64R3Knd1vLyR4aZ0JN1ccH0/ULJ3KjlTf+1m3HZSQtDLvx6G6Oxqj0StkmpLlA9q
ZJu2ca4henKjd4SP9bu/0xW+nCu2+VXp2bGi8knTT5fNf+ZaIm9wvjDRnbkDwMbnTI5b25udDa9J
vRP8dnPWnQkCQ1ndy0iIy/k/zn3gi7+J8V0p0K8nYpGclxIp+misix2q4Ddc/rbidLPupiGFumKH
ukeUf13+pU+szwFwnKPA1GpfsHr4jFj4zRNuVX+0iuNxTnMc5dKV+ookl6yxgNra8cqZWwYpys5P
dSgT9fYIBG7HQF4KJKbek5s9SH6tqsqMWbwngehyZHmrNBV43oDmuFVo36ZrZyabgM7jGsDMnU/Q
L7hFi+FXOEMqg6+JO0dy6fr8+j+IIG9U7Vz0ARf5pRlxdQ9+uqxdaU1uJf3X3mxYQH91qhKHQgs3
4BQ8yYr84ae7BvrKLAxwBe14cAKaYftK01QUgyKdi1MfqjE3iq4rwBERZ0NXlVwu/JAoJCNWID9A
0UN1feDZ6HBQzwgDLAno96G93W1LUxSKOdqnUM/VMx2Ph9EfEyg8HpBwdnIiIDpx7jVrPV5GsvCy
W8sXITHMOhEmXKU0GuKtqRz3YaESeqGgepgv5WNXwGq6Ap58j2kzplbJzXoqc9FwRdx3926EeUJm
/e7H8rbtykTH8BdTi2aMSLOdcg4sUmkIdfuzBTJC5O/OziFG2mftkS8HR9FlmojPMUMDuT8XUu4b
bzL03swt6VZQjLXrRMIwTV9aXXbe6+2yl59W8oS4lzohobefs4VYgMhZgwbWTLKj4K7/O3DF8+jU
2ExBAe6J73EM+FSDZeNyUb9/Hxs53WImUp+ojvR9vba0QOQua+c1/Zj2KgQTwE8jNxnlWfyNfy2B
RVnU9J6Xn494cj2D32/5EpBhbriEJz+DTlbTjrgZ8pR39KeA13T1XIWtkzVmF33VJBJ1+4cH2kMl
0xUxXKtHIdu8FZmbyWQZdS6uZVsyeOTKbtfbN7qcEbqmpP6hyLe7OiMPFa0Qavp7kVOoU2YhB+uh
s9E8gQIEUjK+VEmdBXSH8d/fEHWOIdPJ5e+L5OfzNR7Ez/g/acIACj6Wnu/UktESKBADr+ECuKSh
Q7fNgDeGYGcCuPkJM5Q54+IId3kcO2BiZjl/DkXsRyGEBLujXPO325tr2eSlVTqZJYuvNcLAskPq
636928ZJzxgiJ2P3mx9SImyX26bmbiq4uKPyL73oD+rxDja298BYrsdrb4HDQKnJCfYF4NjexfGK
ziAdexxTBHvES3KTpMYyKisp46v3m8YQccV94keguZRPOexObjb/1OJMK2pmojMfFiPInGEKWPgd
WkCIpw6TKp1Hti2pps9UCRP54wW66vEYNd8gJhSTs9WQwgluqgbhVWPJXDvLQn0tnQ669EDA8Dab
JWkEbpal/+OEAhYh1jKdJJvTxNmxUhIBkUitX8cETThz1oBxFJgUr1whBPGj5CRmree4F4CbDsYX
B+9pvTHeVh0WsojVm86w9oU6FS2Jzup+U7jind8eupyxihNBPqnR+BX4kOAg6bfvdES9XV+3OkYl
7RNgUK0CNLWBbd5ZlJMCE+84aBv5MXk3ZhcufnQrPOGj35PrAhNOWko6Ipxin6cB/utnyer1p23B
ova38sCpE9op+BgBc3O7g73tDaUmhmZZQvlW0ktCJK03VK2kTouuvCiUibJU6xpDoRhLm5OXzrx8
BNDctnGutz5Jus8fnU0usdxUBwYZH7qmPNpmmsUZ02KiIKSNA9wPt/Cl5CcFdCz1i8CXsHbESUkD
JD3cGrHN4aK7zvz0MFj3pypSX+YiYSNHaouaizjxcgd9UUpeNJLlV3uBM/V0JMSOO3p62xgL0lDF
CHhbvFYfKfI+4FSB/jh0CS86eRToyfcS2dF62iLfjp+9BqDHHAlMFGWjeUo69+o6CdKDL0ZlCj3K
FDehKkYW7aV8DZPwj6FAKhtTZ2tkubtK7CffnT1NnTiZM2QS+NER4W9VU9YQWnx61YQtpxKjgN+P
LshFQqBvs6tco1Yn4CyWybJbt+t0qF7JZxHP+jdVunlV+fviDLjvBaDp50hfxz1v0KgPmUaiCXsE
+UxSpvbatDr7smBrnRvAHDnyMUGIfUGMxUWaGjPQZknfpnjKGSaB7fpPoKcpcqq2JD2bh3GjOc7w
m2tIp9qxmCJICSTiXeRLWaFKFsWDPPp2AE5tW84q+3l29OiDUcTY0bg2z1OzJH0rfNCkpmFSgLTu
dU9gN9X+vvxdquAk4BTnS2RMJVlxUO2Gz4p7AIxGtvwEEKpx4noOjeVKXiWJZxN8533E/GPx1Met
la6dZlgUCSXC24R26hUw+Dxz1djPZhUUcJl9lixDviIYzB2gjpvOoKs6Kq1ppnJbwMxXMjEKY2ZL
/cj2FuMcPz0soTzt0FpYw8WbPlWaZeCAp+c0I0YLGL038ORex5zHhpBG/mU35CKH6mFjkVe/nJ3c
bLTG2SyOYexiMlU5komMbQsjpyI49tdKoRevtFzkfxX24nZhdBflG1+mvUAZzmNTuKw6kplI3F8u
S/UmAuXariKLCg2lukeiyuzUu/IA8xR84pn2aLt5RqklrWV/f/Wm/sN1H5IgAA5MdumhGBFKPCNP
ALlnak9pBJ4av+W7B8tF3qDmRSDweGuiHSOAXJmB6SMiubL4FMCl+vKIW8RWAxKZqHG3gNay+lfB
mSomfdM/eW2F6IL1jo9Da0RWoss/hx8IgmPwtNaEAIM85nxiYS+tHI2A8e1XJMoLY2/evnkHNt3F
mCbUHKttqst4YLzy7Yt5xkhpN6s4tQ3okmek606+ptzJit7kkH0AzGQNuhURGkZ2W4KYVqDYIp+d
dmcceItBJe2Fj9dDhH0GrxwFX4phnUbJU6OP5NPeXxwvLAn2NG7txTN4PPxRLha8iZRRBF1kM7/a
7mlG9F9nj8FZKYT/YEtGiy0lZq/VCMlr2uvYRprTPt4uq5btzcwFCz6aHts47SQldaxnVFl60JQh
Gkgk7jRRXdWAJF7mlkUmoZhXSzwudyoypNJ02NluzB//lh0yODza4itqL5umSHqIl8mTPqziVv8d
gpWgHFRjcA0EOdFce+Okh0X5OdNp3kHJuUy+b9dWorx8H6cQKbat5/YfAiqS+mxwosyIRWsr5yyB
aA4gcQ2DRDgVLfDOU29PJd4RQDGYgSqJpwQZ27OFXr5RB9OfalLd3mPWwQUnL3C/3Adq+rwuDe2X
JsSQZ95SttATF7isgz/Di8NQ5lcIyVewMBHNIZmZOz7BbeUSnrjUfYI8MY2mSzcUYQqYEv6llsyf
t3Qaz+ElVk7XSX4ir9h0v6gOEmQxphSH8wrLev4mQeykzTpgYHGOgweKREd7aWmgXn4n0ABHVGAI
9IuY2dA6M3TxLS+uV9xLMDd8KX3hUnHoeptbRwaq7xBU9U2rd5L0QyF2FDKLHjPItQ3lB+h2rcT6
wQaBoMRtfGARfi+VmnxXxC9RDndkD3dDWBttYXFaanyLOVBjT7pCLrQQn4CeNKYrkNf0nIdZgCZc
lVlpey5WiPCMYKkE9WfyebT8EuxTonSl9KBNHOySMPZqrH7SAfEjgx5Af7FdFbkM7Cx1sMQCQA3g
luTDUci1zMAFox/uBDm+c2Jrbi41o5dAEA3ILV3X3MdfQWNyavKabbNJmtAoiJDMYdwu6JRELZ8M
r8JKQQhF6IplOPvkDcfqmCovofVw8sXfjgheogSGNLJEkNFXgyq9lLetqzR/Im96Edju1ty5eEeE
hd//CQMHjP6/yZ70djccgCAudQZtpUWom6dnYYX7Qhahkqnv7QTzRE8WDt8IN1ZBWh7mf7MGeaxe
1v1WClMIijYxkpK+Uo92zExa9EtQD82BRa63FKf0bNVrVUZCcr8RSchpoA6MW1o0Z0hnxwL1kKeu
r3VPaz5V0t93JW82Az6gmFpn7zquHjjEHsbUZLiJoLU63iyssH3lEE/1/hYk6FZKBxqcq1dJnDUi
PTA2mvXbU9571HbLddb6X3mBqP3Lfp5IU5SA+HypwyKsR7h3EtvC4ZMvVaEol5N8fl1RsqxhYzIq
zsVFYQwTV0bGUX8qjN2AbSEKAlbxc30W85Pe6O3VOFTZrzTaBL35k69YG50ExhGSWgRLyX17aqJj
wlPJZK42MISVLhVtgjZSKhh/6i4YC3pKT0Uz9gGFfEkDyM7OVSEY+vwNvfUZfHTiji5yBIyhYY1v
0TcuY610PzA4RUNI3+w4WZCpt6gYIinWi69mGwijowZWiaGX6ZC30UsiV5nlYLotA8/6hzK2gbig
mXP+7wgOo3mr0yxIfl9zlLRSWaaVIgJo1ObjRMCiRxWKMW4rKTL3IwxB7x9C526iNgQqPOJk59FZ
6yYu972B6/HuRHyI3/9z2/5PevUpkAB8Ks0mLIQcqD865+c2JOzPtStIzgOFpP4dvJ4jJkwt8ORh
0U0FXMXXbm+qkWAqWt0zMcQM2DcUncYKQGpQ0qPfo5rh01W1FfgkRp86X44Hyt+ovi/L+5dWOSmI
kR3RMrIhB3MV/Sf4D+lgryF6IGsZf6EKvq2QpyXjiiCW1/t0YQk3vt8HxkU6vLWTlnjUo/ySK9Hf
FKZmGkBBlaQcFO59SdGQK9x+tQ4yE3d8Ez+/VCITcShcY5JxPDBHoNiWF6OQYvImCZTrG2txBeHO
npxzu6iehT8b1beKXFftg3Ez/t2c8IE9PDc1/wZCwAj8Ox9zUYOBn0fTNUf16YUhkW8vWt5kT8T+
8RzwwhixubCo1yV3F+zjFfxyibE7GvBwrohb4lfLjVlZmVlAPlgCjIq6awtdfEua2c8vigjgMoS7
kF+T7KjNNs//m3u401xhvLZMhu5U8tc7J3J2Xrj7NtexWV3RC8NYhxlAbYkW9rjUCWJsbb+if1MC
J5LcJVQcZvDUEWL5dV0Q+O9jEQIJvhV/7fBwYvEu3u6T7bqopDaGFlVkS2qMfoMXOKWXRE20/di7
m/s57wyLkvLJdoCTplronAkR0pFyjnkT+YOQYu2BwrRVh84tB4pS5xeXUqn6JRYjxHZ9nj02NcUD
G0wX4ttf5AnGJoC3+SgASnJdmdAEJnf+H0+D4wA4LBoNqGj22EtaUxpLcOuHa7kqVd6UX3u7bJ09
Hlb1YGNGJCo2JE3eyDVgRa7XpNniWAQbELEBPJGD+sir5GHHMj3Sv+P7TT63dRZgIvZhZmlnRQ2u
DsxHLVYcnhZB+Sdg1TEa17CFWIdvDGuexbKWRAwHcM5nZFy+cqF3O/jFW3UvjSFQsdCVY4L8novt
+Fi6PT/ZbS1uEAdN/dMMDQWZ1P873fhABnvpmjOH8W2gYhFYEuauDtvqYJlmqxajRhFwCqInz3RJ
HSL5yvFel+0bwYle18jakjj71z35O1xqVf2OzcyXnAI7dzJ1lr/ptJa9Y3t5p4F3WAIpxsigRqkU
aXkXICo6VdimZf6yLnl2RuRJdAISLtPUzmE6HMvAtlICrSkVlqdnUfsrY0ur/FbFNf4o2nU6ERRH
bI9uu60cBD4OsqmwQrLRJPqSXaAl135kkarqbKKwJALwTi5WBjqy08e2HpSfrvPsrNkxX2OOSVTW
QstWM8wekTVSEA1BRNEDe2QuSqARNCl724oTBZUID5zQC9Ajkhwi9G61eXnxJ6TGy2Dpz+mPLMA6
8MFye5L83G6iNKH76LLLf/e+pNOlZu0QDey3PYtEqXrwn1jiWRZhEP/Scr2Sv1X8XAfolKvSQFW4
fXVzMioOEU7O0BN9tCgHmu+i7qprJet7w+PyjfOaLAxSkjO2ifEw+HW5PosATG4zGB7tNG3WfSOS
ZC6V1l97KBNycu0njvM7afx0mpHXxUbiJqwvSeU34UXj3sw0QvmIxZrqJVDiLDvhxBk3heRSCEEH
fmRmVVup+VbTD8DjQhiTnNmFhVY/BeN/rAyiIVFrgOOk8URUijkye8bo+GGIdR+Gonz8uOUm20ll
lJh6Aa6pR2sUGO9GIHO+K9ykFIk+ScnjsA+mk0l1UYv8FunVGhXe4a+OiVcy2aT+9XlQ4FdZqytQ
Yx3anwiiGWnEvb0UR4QN/sU55jye8k+emA42fcjRaLlgzrzW6BSzsMWtmL8KuQi4xLoNopkV5ch1
SCnvR6P6owpOO/mFbHItnvGHVs3Ymc3sAof8Vk7HEDyzugpiH8cyLGHyCGQEH/Glvf4KmBUUFOMz
TGVxgGnVH4BAHmGgXXJ2WBHW4DZ6pLvM529IPQh5l8BBJjpwqOSXxFcmlMnFqTaV4/necNg0v1ul
+W7Px5xfbJKik7aXIZvBQmhTb+GB3DcRlSWiXZQnlUzx7LDC8k0n3B1Ih37bbVxyUFn/mHMUQZN1
mAPZzPGPWDKy6A0xbSH+yvUn8tOtGXyXocry1D3YdlkMQmTORrzWNZLdJSlqvSOHUNLVSIUDAthv
jMLJQrfDUtOnqCyXBzcOJ59znP/hT82XqxCsOEd2XNgTOEIbz3L+wZfpD2z/4Tw6/RK1va2DM2d0
nAld55gO4PormuPh88q1qQYkVoW1l3RJan74PxhBiVOtsKwt/PBmmTogyelx6oE1ul/M4yVvYGuO
JhguhTxLAdW7m2zw9ZeYS8gEv2ZC5MXQQjZ6Rld/sPeP04BiJOZoXx81NqsdgVjZDHRq/JPbzWtr
3yKxv7KIOmIwpCPkzMjSd3UIMtP0FyCvA3iWBNx+sR/EpjkOeH2JPagCsuwp/XDD7jiQ95rE5hD7
il/zP5uAKHNJEagdNz5siyq2YrytVeZADuOCc2p4LQ5InCQj0a6CqDhwqodUnvtB1BjwykCXevy/
pLfEJ80WpbkvPuAvLsviHQei74ttG3mmfwYmHw2pP1myoFG926XoQIXYorp8hru2bkQVvuGmMpWK
iwDR5YMCL0WGJgNy/N2IxKSJOBLVw33374ay8KwjVZTGhIoa6WI589KCYr3wlQfv+5apILVmh/KP
sY16yy6n3p7W41qjoFSJMruzZalgAz9ZHO33fqjNoWHun/mW6+lVnyhiZaFDXGxXrjopSOTQ0u9q
tWCLg2df4tB6mm5FGuSPGOsMcZcl2hQap2m4NnYv6ayfhtihCCvMObzlLq9F5A+fvPy/uEa11HwJ
/OWsluxgEBU2k5Ydshsv8dzErxnDoBOncJz+j2Z8NBva1bfcg7M3z0VkjWKP1/f6F8MX6D3tGyN0
d5ksY40d5A1OtMJC55iuY088ZOphwIiHWZahoQmP81rFiYt0Xz+ioW1QC0zvXI+Wgs/QcxvADnO2
UjYtK8LV9pcs1YB4OpD52rx0nJ6Si1k4Y6f/nSRkdSjQmbUJ2tRCDsfdOziwg7zHBLoY6oUmVajt
9mmd0LH3of9jwZjGxv4RKz3qs/vxW3wdL89AJWqmQGpPTADNKj7c8Jy+JY23ppdkgHXlBjQQhVmT
aAgyEbUU2s6CXbW8je+xLdt49V5xtLDPpQhof99eLpPWMJ9d14JbCzO/TBvolnNO8GNkPlBb2gl3
Atnwu0SQU7RNxwH7OPzGeOKRE/sk9b3lk4UL8dj8spFblAeIODmOOnMRN+FESx/cOnTrmPuzLbQ0
CW733DW8pZQO8CX41jRAXs/BCHXDdBi+rAHkXa+4CsXx4Ti0GqfFuykGiev8UKuF7EJQoSePNZ4V
X5B7Z0Ou3mFhQKWBV3InoHZT4qVG4xN3WpzPJLs9uVJ+6Ezhdf/C+aPMcOY/nCjg+olhbw02Q9Tb
gLj0LCDVZHmMGcje8lSooiHie4HhRVpxbHGxJYhTJEtjCri3Ri+TAvsl4gAbn2EqSI167tzQzoEx
lJoM/kTB28zZvAzPFw3hGuOU2F539xOKYoARsrYmWL3FiSkOHoERq3yhYC/kuvbUq2hkPly5zOw/
LhWqMg9eVt2zH2S+T2mZt4/fqoMHfdz6IKZ8YCQmNWzdK4udI+kXTd63GgrASdE7H2pPVbTYt1Cy
NeCC5fwX7pnM4/OL1vH0YAEIWdU2zUcNWfG/cRsPst0Qvf0dxUqy129gR06ZBP9t5cE050xxfUzx
CGdRgGJUl28esVIUsJWgDxylH0DKo1w1KbsKzOZrui4BJR9em7KH2r5NQsVthELr2pxz0LG5SBE+
Xb7XVn0bS7MW4GSXx2yXX9Yg/o8fFFCga3jOW36wU6qyXb25/tI4VHlkppLDYG/F5FRVym5lxpsr
hupnqR6me2wb4AYQ9uRCtAOlg930eavTjCgovUFeHgv2qH6KDUHT7HGuA7jQQ7HhY3WBdjcEv8xe
Wzmy5r4iS2ExIHVvQwCtXrsx1IOaT0Ebvj8IWigM4Tnbjqkt3NR9Ie0rW0pDE6CSOeZsFYCyI8im
77LHZXKj0Pl5jhHXKkPv4ld4lbhDj92c0mBmkUG9cpgb+xLbw/pSnwENBvhskoLUWJ2j8jc/7o7h
NzhpkKgMH7AIczDmaRGUoB1kwfX7pEi2gQLuzv6RR5qu7kyWjQB/ItMVymuoHqznM7VMMI5DvRCQ
6ZWq8a1GT3q6CiMSfeFyTTw7RZ3Q4BSYMOlqPHztEAIX1/LGo2e//uIWA6aomz7cItv1ggAbtbLZ
prdQ9NFeZ+0VwYY3eW+r2kf1kkzKlAYY1FxDxMz6UrbRjE+QYmiWOMqQKzl87BwClIbgoO+W22Xe
wuZDOAyCd7G5/wdqYalXHhiN/1dDMpxVDwhT3g2NDOGaIlBXHo04a+nIreMulvOrWMXfgXNl7O0f
e24Q2I4LL5WNbD3Qk4WiZSwn2DLVPT1fZzo4hu3bMu8mN1ac/zLQl+Ezh3inciJDaVFbwZttgcp3
oYnQhfQDqgXw3qt6msbLcp2mFdxERqXMJch1mfesI+SACxXEm5djVEZ4XGccw/OXwq3Yxo1gN8hb
Xge73CBHngJl3h2z74LU0K9h51Jzn4xpwc6ULMyRF++HSSv0ZIoCJ0A/WyAujETnuknkjUzb70k6
Pt2UcwP+jd0Xu8TuEgIE03jxAURbfHdXmPkliZfiyOYFRejZGBXYWe5zCMz8yPmtYtm+mY/zLsbg
C5OUKtmM4qPEl2U0BB92nJBDbI7AoRQe0DyPAl9ZGHrBxj8rUXntFcuP1mfhQNdZQTEI3U9Wsj4d
ucEs33/PZZHWHLUKjrKT114g0C1Zt2coSMI6iKZx5fRT+o02G1evEBKUK466GpKnydLbaINtXZtK
wJXhPI2HWDCBzvX/3m+a/vI72JZb1VhRzcyNJng37rJvTGyy7rULVhndSUpgV4v0nWLFvBCSN6nO
Y1vJvqCGb7wr8/U3SX/FneEnNjl16BrWe7detF8tlNJYW5rzxmYuWY5MFtJWurrYbNH8Zs8eQZYD
VxJy53aWFEgCmNt262PDZy7uh37SmW8HwgjKh8SV2aJHPL20cucsMIbMhjQA/s/WZNYQi9r2xoQo
F6fjj5bTGZ08dMaQKqUzuoGdg8i0ufJgwvAJ+Iys2Y48tXsgo56N8Lqdz0Q6v0HirBSJbvApWiXo
/qKI23p+49wRVD7R6v12pqqMnA+4ViwCk9OQVnHXmGggR+7OHPd/k7ZLWQnh3fo+B+Za///i268b
HxDgOFhWBGUMasJp2i0MnMmQbPabpBRvNUoIDu+suNq8mk/IWjbB22fNJWbf5Y3/JnmSgEYLhjkc
pEVKOp47VBYfWTWvwU8w9JkDrH37CGZ+idgKnPK1KPL2WluBsh1RZWNVwbh1EC8PK0FKyGOHncBV
HEgZB8+GrquQRJc1UJj2g8qld/mtioLNchwHjylgjw3+2Dpzc2APwYb0MAwxcRFJ+ane1Nfuc2Pb
0Wv03pLYPTdjegTd6e8SebnKaXwA8fjUkUzPAjOjRr0CDvB/YTNoPkDyf6VVzFFN3kkdcq1I7N21
GBcBO/d6ug6t6pvq1poCTjNqwEre5qRkkX8sIRtKonwTFkpEu4ig504dUn8K+CfGKBxOjFT/WBeg
OaWEz4SlzPLBAha+es9VPqt/mcmm/m/1WIlFyFm3YCsXuXPjv048hAlwV8DLOkBh/oYmP4D6iURz
PYxVtkamHiwGKt2FvBiRK4L8n1sannvHWknI3W9luvg8VLwPBTpZ632VeQAgOtIt/XK4EnJGY/An
iW7XFdKOhrgeXNjHgKd0HvBx/R0ehyx5Ls5C0UahU5I7IMNutOqPDUL2BrVMM6gH4S0Dh1D3r3EX
R1BtVQjQlm6Nz053EcbE0vo3hpaD9eY2DRaQQUKPNWEAiOhrPay315XSCpWKBsHc9Xvq+5WpRvoF
ZOwmjhRg2Rzqu3GJP3aCVGOSeHSzursqToBLEu3gYH5f4QnDx10ilpcBQSchcYFX3khjiCVchfs+
cIa81OiJhPULAv9v4dKsbM7EZQg8ZQhyOcwrKxD+s4xB9APZrwOKGGSfvM7mT693a4Qodqq52d21
sLESPnF5j+i4p1Ui2Svo8u+5i31/U8W/kWv+3UZOr2m4jt3g3hgKCxYozqplPCdpcrNEkxIBDuhI
MIyVmvMAm1lTe9wZXgFUmaMxvGKnleQxlEUfsAOYkbFYW9hD2dauDckQu0eTMfef3C/Z039ee0+b
sRyGP3hPOEUx6AnWlOa5FjQf6jYabsyTO4PFTj6jliPrQUFIjH/zVs+3W8igQHA1dQt1TssGBgmv
ILgKqKLEyO5RsviFr/pzIa4niXK5gbWdvtdC6Q8TFNsq3ZeDxkKFfl2CDwoo+fCHftgfl4TgILef
O+3mGyi4LtaSWneFR+tfN0fBDn3bq14zHdPB9e4eMHYAtV9SQ/Ju7xX0ldaUX+y+OCkZmb1Nluok
Rsojcwid2/d+dlCGAKx/PiRmBbaCpeBu6LMzSBqiK4WoYU5lEmWQBc2q+meTv7T0P6aPVz7TIVe1
qb6k8OT+8xlK71G4TG/ix4tBupGyeExJ/GH2ZjedO8wG5Nozf24HPXx8w7sYFssqiJyV25NZnMAG
k37wfNkwDhRtocr4eX2S35zh1yU0lNO/KMs09bgZMWpCzDYddKLolsbZKkFXLSqAjsuBxtSu9FUG
/h0dGaZ5PMeOCeuZUx6Sd2MtcYEL3ws37EVf73xYgCVyy1RbCQplVWiiqFaqc8TyrZHoaCW/5Jir
4wYNOM1TH0PTUviGGMNHrAUPbDakZoK5RV9VRLM1ILKE0bwNylCGRx8FdrbM4Q3E3QA/tbusio7+
wto2aDdamcd9ZOEH1tKNMf4Su3mSQxviY5oSoUHvcQIBoO+gE8gNnldzKy8kj3CB++h8aojZdlhm
qllOFWqYu6CMBtrf7TYlo1wMKfYcsP7ch1COU++uM5suQy2L1OYM4yl0GZbcikVihX/NXlq2vSwF
/3Jyqox7b1PO0v5TU8TWl5MP1ZRZpBCxL3dj2Lckt4tQovk1Z+7kJcYxDGWHNfxQfT83wriRdId0
CL/tjVHJgryeRrpTAe2H7sjzf58cr4qbpwbiDj0RrRBdo04tqpvrq3UUlEFvgRTw+TJ0+MHevryQ
REY45nm8ALae64JUnmMl6UE/dfLRjFLyt/9q+cKBx7jftLSpvG0KMrbtC+qAFpQrtgS7s4NKWpKA
+c4f9ac5Vf8bV0XpDJKh7eIdbZ8MVX4AopDCTywMvE9N0llV/B+cVhoJxCUT//9C/NlLGXc5blwZ
0uRN579FEMuzvc5R1VDE2N1oiDTpOfp0xvfX/7isqihMYjCOZLM3k4uXnA3187DYFq+dmKM/O12F
s8JmitnKvlL9loKY9wCE35/vxW+maXl/L7WvKNZWPE0RYqIBc6RWoUqbhXrrd8cbuj6qOwEjhNtC
BcrDqWzBqoi/k3LrLMIC9ayAjUcLC6Q39XTccUMpJL1dzgaXHArGdXNV8TTkmapYygjXDcaswqDI
t8lDt1wGlhZwJvba8l4829RovzaFIcxDPrRpPaJFSd+iVh15041iHI3sAcazSLB0uIK1BRvGaiB9
/EbEYZIt0Ycb2mCqDX4PMCqMM9eJAuoshtnxG9nI4kVvt5uvh4rf1PupFzMCJ1tfrbIykC/76LW2
TB49KeH/hMCG83oyR5WNqnGMPB1yQSfkostipOhYMNeMtlRCCUS2EZ8/IaDNSIXgTVnvuewHWs47
u+4mOljhlnAg5JOtiByYY+l5sbekMicN0+h3HPK9oANhBRgDt0UuRLlhyUc5h7sE713iQfPySv04
G7v57p7+m3nw2d69GcQbW8t+YhDKdktUh1AWDnFIKfXYks8eS52mUm3lRkySodfovHLzWGhe5KqS
kLNpnI6vlZ/B3LNctv3Mtga9ygWBTGd5FWRRk9MYkkQZzVNF339WOHpQJNnPbz9Um8Nqx2Lwj43h
eurKSK+CA8srY8mCoWEBnXUMaFXSUU0LOV5wTT9c4/qNbgtR9+EygfnnupmamwfSIBuY2mycwrCT
3shiY1fXZQLDh0MX+FZQ+v4CBLj3avzxNIykgojWz75wM+ChkICQVhazIu0CbzdY0ddjA5l9rMY6
FLnYsYpA8w8U5igxZHdj7a5V1dB5EkTC0LitKtBnVcG0vSxk2o674r0rIkOkR2Kb7e1RMtXcP4fw
fOX2c/F+qCWu6dzWCy9s01uWCgEpbozzRyX6dylyHS6MUo/ebGGFCeUd8Ezk889rZb83CxT4ojZD
dU3BELjrKJusif8ywvcFl3eX91vkKYC+tSWzxKqzViGCEaxavslH2Ex0CqyqV6Zcmf2WramYRcxZ
TGRlESLdAvZLdzygBo4hLhDpv/l4wGGpJwRGgOecshhs9VEcUwbppwnfvLsXOTB4b/73BuJlugSl
8Ug9/IPTyoccuWtFk5+qTUeYXbPlT3ULa4qvX8qAEvXcPY28wNLkSMVZXQTpxk3dQc2zILCp4jCd
bYev2bCXvXNGJRXgv3701A1+wsUQvN2vlK2H82uLYGSkNNEbf8oYk/bUM7Ljbah70r8dhj8z1sAR
yT05QVdVAvaauR3wU3C9nn8tGQJHyIvQ5qvt63QS6sZ2lWVbioDpDSLmwosJLVfcygqTqYabaOnV
+mGtBV4qoiR+6qfLJCjj/Zslioq4peErOtOsyaxoYL6Q9gtx7D1zT5YsF71dpBPvIyKEpjbqsSN8
1cVvmW2RtIpA7baeAJ8bSjNMNJsrW3HN0yBdq49A2Ht5+x1fpw3IYFj+PRYbIUcITpo00p83OWXU
X8JgNyA1F5tHmm/lnLKC0gzjd6M3NmO7JPLNY/pcwcCp2qx+oVDG6fQ/UI67w22vAVHt/Ejg1O52
aYEFZRgVfKKKRQ8nQvIh+Zst/qSsi7TXYnO3SB6MnSmjZNoYQIyLMo+AxWwZ0PL239S13cvtqvt8
dTTyYDF3GMTO2mDbz3By7onh4/WmPy2D8SL5KwOFiFiWpdDmWojIsXuM54cK8oGvs8BnblXoqZab
Zg3Z36x+2kcldGIBZVEJN2+bDNx2fBXetJjeyxKURaYcTZy9XGufd29P26F+UTI+kewsNwqESMxE
EjEuQXzRfBm6ydA4tGE3vue4d8qw78wB8Xst8S//pxTWlUpZLHFMIS+l5vsfIldC07ZaDeNYbFhC
nQ4LwtVlZxm5WWQfJG3JwPcgy5f36CDkv7YoMJV0E+L8eOf7AcY8kDkFHn5A/l+gw76NUsIBQcYn
WzmREJjCooCZkp7DAq19M5GJa+IDpsRSKMMD9AX7zZG2Ld5kiIuDAv/NfhEDrdKe2VVS/BnYQuZV
47IAEvOXwot/Nw42w54PH7YGSSAXbrPOM/R2hq5YBUhhNSwK4leBqkVbn7mM4icsfCUXRxHCOWBV
ARKHUPxUHSB5gyViKG6xqhIEqGhMUERYSaO3lrX/Q3OmlUYsBSRzU48qyk8R2Sr3SpU06hqMmdAz
Gb+7eNJDj3ZVy9iX+vkcpjCYXtkRq+bpXwgQRWowOaIK5MiIdXd2IdoIx7WWX8MX+tEPoT5VjX+O
fPWCDQk5OXYUv25S5V/omYnvIItzq5ugnhLJujGIrjYClU7HFpeoyxVNrutWBdTu5eHIj4r4PHHv
ydEceqjaNaxyif/h71w/yUAozHjHJykxaXXRgxN5LsvvT7x1OLPK7PINnev685NiOy3M4QrIiM15
BzZdwzsqYSNINdTDwBzOP9fYt+6LinYN5EYVHgNTwmEhV8cjI1jRoilKCkfyWQ91QQ5qCOPMKBo/
621Nl34nS14plXwcnhsluy4nyuv8U3h+DUvoEPJt3yCAECfM4b2WN9VREANkq7WC9+B615gXq2q1
7SAhElrdviGufuZv2YQBP2JHA5M8esINgu1v8tDBA5h1fMNngypUJG8Ivky7eZNBticzQYoi6O9r
AjJ1atvSwko1cWci6tX7MMyhVxaIMeib6z63KUMkFA8K/HuOTEYdcv3TDW8NyMaB9w2LlEhYNdOS
+lOxUGO6yKpdxH+w04rNU8kXz0Qv0CXWZg496Btd19Q/WT6uh5/pKyrVYodxYe3/9vgt0q6uYxQC
Bg6KSlY0MKH1GAFdktxlxsAWD65dVfl4nsYAcLSpMh2IpfwaE6sGY0jZaQhojRMeezH9Gt1tyeZm
l+S76Kco30E6HovjL8uSzML2AdMcTVI9sYV7/lrmnVtIuR0EiFfITvhtHBUgHjjZYVG+UPi4B3fQ
zq1IcS+lRR6H5gE3yFn9NLbkSm0VYwoIkmCp3+Obd3LODbDUz6ZP0lU+2xSFsEcY2gzK3v0IYBCo
A7wXlInM59IOrd2nzrN8vCoTOP+Y1xFj8tRVReTb+jsNnwZiSo19IkVlmMrNfyiqpkAJNxHbaY+M
7dFZqd78+ooop30hNbaKcgvBHo4IpuG7u20BppgeAE0oEs7viQtrGMFhsBFdRdLxFxHKIvXMhOcR
v7fa//bF9wQ4GleymYn5jst4RHizdw4rvicZsh2tI94euIBhN1O+iqm6f3yvseo6FJV7xUmnzFmP
x/iVSUPhShrepkPpIKpqT+GuQdmA3sVfGg9FIuBThHg9OZUz624UQWBkMCG1mZUoTv8Kx/j593AO
OZ3sJNz1lBav99wUOUPeL70BafgSSPMOglio1x7T5MjRvC8Ncpg5He7NiXmJxAQrLrzZ1rC+/vb9
II52SXKIxD+lsZe4zjV5fzF7caKcnt5+1lN71V3UbJBnEhFVreSjNY1LfBtW4nPXebqEkBI55qRC
HrRwL3lAnizpNs6ST6TbE/a9gZI+aiR2uiE7zwQ44U7irctP0fiI/rG6+u2EvLiMN9tdt+T/6MdK
9rNbRUWdGWOlkdfGFQ7di1QuJaEsxRR+OL8YPmAmfYSvjccaIIMUgVsYLf5lVtdGevr/NbDZn0JS
dJ0m67uzQocqC9ZkmyZxzGFOsNChMRJYKOlSSw94FLMfdry1rOZKBejiIskVTy+fFPAY4kZVb96t
girJYWx/HYPEamiMqu/JE9PNX4RxDWOsmH0LrAvRkdIJAegxk2ANYNlTF8vT6QdI8veoiIJ/pJx+
56tb/umt2x+fw9tjVpw6W/XBzKFADX3aTPbSjOAnZCnslg0Q1M9UV1IIBt8FXLa2P/wyYlmMbh8+
YnHmAfuWJ1iRTdfoqkxL4rCyEP7x59bI7FnYjiDhr5WCG0SksMTEcMcqnKh8whwuXnqzvz3lzxCl
O6Hbu5hlj0nSB2YrmW4R8vpx3XGEWg7m3QQ80G/zmJpOdGCYD9HZPeWO11PQqqOc+Udx89zN/6Kf
HNGKeX0pD6gdGt5y2KZ8qojpuk1qifaTmxC0bjG0o4hLoTWJ9nnmvLDoH8Mp1BD4iz259OSof7vk
LQT7c9yILhq++2XZUN7X5WRvQsjcaCDraPJkzockPKwuSbzdpeegv26mDhLmKruhzXIvbBCkYzeW
PWFtVSQPlS5KMttxieiN04o+ImKUnNnf8DhPjys87zstNQRPGEDY6Iq1m19ugbJTV5XgHD/9vxq5
acZ5gKzVnoQUTl6xHH9Na757VX95DYrW8kGV4IhEiHZ/CK+sw2fgZSRrKdMAFvyFlc58aFmXO+wW
tFpyCGczkgLxYJ4oQzrYSd1KGaJ7I1qiCwi7a0ldNDvsa4/9o8LAecxMr4W01irJb/w8pY6Sc+PO
TH6FiFmsGdYk24gj9tHDlDP+YN+pzeDnEmvUQX+WNnbB68GUBtRHaqCJNY14Ma0J8db521ZftFeH
9/S5MyH7ZHlQKJGAi9n8XDZbxFzS6rma3gvhms+l+KsH4NXrjYCMO6GELwEGctU+ufMQFknb9drF
pYsEZwC9bHRPe9Rv4yDuyRdK1D1R7dkyI915LdDQhuOFwFGYCB063vP1CEIPFtEjYd7IxPKyMP1W
WkWd6+fPlSoou7MU3+C2V0OrQhNeCShiQvq6n1iMOEeO7aAmzQo59j6bGS4pUl7utrZIM+6sELWO
W12S++wdfqnEka0ps3XfuatrOJNKbm24cF3ECEYYvjHKHolZOOyUZPAVmzbiZqrif2dN5HGoqvm4
WYrtp5ayRX9+nGC9j8qon8soiSgO9EF0fnVSd/I+NOZE3Zx7bRg2NN1n3nrqnSVdsCNty0G/XgJ8
quIdyfOmBcJax9+RSVuKosc9q1KQKT5DiyX5Jy/FWUNWeLdsxZ6YS8wIk8Ago9C56vUCH6VY3jlo
QrxZ2vPO1CeHNyi/CU3pLrmRG8nFjC42OgxknvELXtTkkGtzQozVqR8ZG/LrCQhRaS3ewroAFeor
+VHMNM2DQh977fIQ+nB+RTJNF7ljigJaOhFRMiRPhK1fgEVf1nkTkkxX8G5MTBiWBhipfYjj3qg4
cLsV7tUdKKeTm9NozS4YfKYPWd/bqOOZwk/SsFv0JzwFKcwDtzXs2fA26f0zX6TqphWsrLUvwsgP
0+ppg9CjOsY1S4/pxAiHt2eIuks63bcEBnAPpkVcoP9RSs3/1ssLk8qavboFtwa5GKpg4LpirFjV
ZdQSfvLfgvtH0qWnUobhpyLrFTOjKKVQSS+i9SP2RS11kSDmPqTjGT8ii29tG7m/ltHv6pq3JpfB
rfyqfFtb10OPjw1xSH6SqvVLKxXmkrIFU6wb8EI9OdJY/F71oZbD0NJjOmvOazTvWwzsxv7eNZgn
3O84pi1mfeoxWQbpbjafq7M4toCf917yMkXdhT1mfruL1J3iA5NBmwXUYU8n3XGb8Wr4SOg4i2XN
8jTHGP2w8GH4t8HNEcuLUd98M35oauY3PTGUY0SHkspQ7b92K2oc3HWwf6eM/R+RS+87nFFdEfjB
d8SY7JdUhS/lOvl9su//EaId7O2JsL9tZENEXyK2VSs/6xxY9wb6TNL2o06KnOGS2cxHP11xYHZy
QoVp3DTBmiMooUyGyDK4sqFm75Qex/uTi/8lrPOeQJHt868T66HzHFsChKZXi5Ag8scmjgVRSH/R
3yLX2L5ZVorml5RwkqCLkSd+C2cEyjknUvXe4CAV6UQcL+U6d06XxEPUM+1Ly3RhG/yn8cPtInUC
nIq5gE2a2w8nuAKQSi/QX/BXiUrfQy5O26+BQHtN/CsjMxhA17VILGkGEIac2Cl/YlX/8fpRWTcc
p/B4l/0cf01BehkO4FSPEqeaj/uNMxQgBciko0s2nlJ1nivpk+8HCGs0Viv9pF0yb1amaHRhKlIX
xMouWF7weCxDu0XjBecAI8YpWVqUblRA5hA1TK5iWVZKnMMid6/S/Za40GWygORth5PKjTySH6/F
3pFr45RVD+3N+PcOfAWQoOPwbVVnnRboPQbV2jgVNxXK4BrPcncQ/7VNHgsCgl1Awg0f4NI8MQAX
R4tl7Jl8qmiyT3DearNB4GZpWoC7SxyfJcbFCHXR4dAGhuE53y3a5V6J/+kqtnou67XHj4Bvj1mo
ApwsNkqsyU4bU2bK/G/g+ib1S7tM0XJ2KVBP3xX5Iwvfev7blU/cLOqlEgO/bWEO7SeZ/m/v1OQg
E5LFhj07guxl/vBykE4U1nDpOKQjWcjMHpRyV+Cz/H7HYRtsU6IkAypfvdHzW8UV8uXpS2JhCoSy
pTwiKOEQWEwn39i0FV7Klv5D8Jp9wBrnmKFNvU8ny93HuWjrrFlyjDTIQuIHGkAF4oUH7eZW74I+
SJw18z3jkAqyrb2NhG7luIPyrqXIdWfmPeUgO33Tsl92dXKHBeMt7DEYyVPQgsRXi2sOwp/k2FdH
Xw8qmAs0JyzcPsIGSVVuxNnZ7Qs4jX7D8H8F7862E0sL7OSqI+N+9tc3Agtr8kAKFr6n5II5S1wR
HVcp8fDDXGkE6o1+P4+zKJlInJzBBD8j1N1uR92awfyhMAAwUL4PxghEHO5N2D4xrO+34hvIi1aO
NMrxhDdXqH8BWt7zBC7xVKUxT73RQrTwATwT994bJ3sWQd5x+3Gmg6glLBmHH1dF8Hz5L7P174cj
nadpUlW8zFtgN1PjrVkPV/QhEDiSqTxMtvWVR7Upo6N+OndOG59fxATVy0mcGzdrNPYiD/mOgJv5
NyTfF0tIP3HtRCY7bxgluTtery90sf8oLZHTxRjSM1W9RF4GgiIIp8sG0HCt3vo+XGWntVbz0srY
cO0iMHINm+qiL0Btu626XwE9mvyfryVXisD7i7Dn6JsFA+nrceRQ5dHuF/PAg1P1Z0qXHEXOqhvu
754tru4E2+dJp3qEpmSSE5hYesEk9QpmEGG1qevCk02uEG5ozBE1TuQdpv9ZJmj3wmeK8/tFB0KI
i/jyzt9wzvHQUnzZbIzazXJTdFRaZCtUPSN3kFB9xlRtwaFK9ZgIeWgXOjRNFtuhNA+RFJ9kVp3W
e9zub9pYiDqyQpPv/WdG04G2rZ0m01uF+PKhu3Z91cNRif56o6CjAL3RKKbb5zJzrOOLKAUuVKoZ
QvB9sJcygY/Vdk5nwMoGfKbc9/8ATO3PwfRWwhBqUO++xjWK+eidWwzXpFEf73J1xmv5zIUn/hpN
SlzuHVf48tTUlfeSMCYcTcpZNXPyTfVmhbLGI4Mr5EpIH7jUNkOI9/lNCIDq9xRWQBAEgpykqFDP
zZUMysMnwkqDJja/Sn+H+lEfBibi7iBP6xAA4rS1ZHTySSJ/0mSsKijSnfuE8jCW0XTehtb2uuv8
4ApBTxiMor9eNDpchd7j7wsHyIZN0ysTSHqPmXybl/Pn8W3s+SuWGOqgDL99DZdf/pk7eW5daca4
1LVpw9oIWfj/h3rVQzjHkETO3TrS9eoWBLhHhIRlLxvF3Uf9JxLjf+mDpxTrk6CEAZpMQgVF1Y1U
vzxd+R4YaUNsNGZLR0v9Pn4jTSbcWjgsmVzk/2VEKRvmM/o5yzaeTHXuaEXZMjBr7iwRm1ce+ujS
yBE1auYFlvDbdn/8PCcGfeXlQRzIz5vFVx5j2OEBuQrvMK5ZHB4BUS5mbTE29uCKhixZ5gfs1Bk9
6Ua01FRBMLCN//Ym7B4EtwBwHYllWmDZ2Bq7Mgqv/OBmH96cZkGPDgC0X4lvwRNp+6Ky0fFLFYjb
DvBKHRXLG7L1gXqxf+UlwxIjh4A4ArfI/Z2PJQx9kNMfkG/7jR0XqEtubOeHTww+ESTuCQmcz2rO
FBqhG3/o/rkDpLF6gXCrbcZ4+qJSt1bo4M+snjwZgeuiVjn/zTc1+pkp2GZmLv1rCyXQ7LPaAfyK
xfVSEb2KMSjrH73sQ5ueWCNl1mNSIVYZufCPzEBxMFYK3BTtrUI3Y2ARFX0Kji/uFBryHWOpdnrP
svBSI/Acknkjrv9qHgfF0TtDhnhzPUdY53Mtyfvh/Xm8NUor9gHHM8JG85EFwR9dnGl30SrsqpDV
nMX+d9p4R/jKdheOj/wX8l3BAMb3ByJK3EO78t+VrMVzbC4GFRa0lJaBqIQodFmKv3N79CgBp5+l
VW+ccNewtHJ3D+kwQWhdJw3Op1OCDLa8wFVsNaWX72jGc1IFEOWRkKaqnDVPSvcMO6TSs75Hit0o
9DCA5t7rnikg6VxRxdHHh/ds5zv0fvcsH1nAQRDIx1Opdkg8CEuMyEauBH8jMX783uSOjz1oSynw
qEe+5fbqHf4PxSMNinfEf0GCsYztY8pCvGh4mgOkRNOiB0IWNNdhHERsCdhx9IGnP3nP/hXwLpMS
YVGzucic2qI9aXcuo3A27Gxyi6k/obLVqD45IR5C46vAf8KjHI7+ed5NgfRKEPCxA1994gZQ7LOy
kTNK7iKyPmxPb+H6DTD+0HzuzIzuE5Zvlusp1U+g4o7w5ZID9AnLcO6zDo2VYaXFy5KyrJU442Aj
sieMtKXwHi0OXP1kvO7V/Xp3l/sbm0QG6Cho2uw0dSoX0AZYIRioDBssFBcLIE1mZgs7Fj23UFnn
KxO8OhZSQXKZC8iujwm7CDRZ6dr6XnV4Xb2gtvr1AKwtUBk5qW9++jHTwIj8c9wSLX9tVwvT9g3n
3qRbHdqy6YvhudoJX6Gvf0wQESqzE22/H1XiFRnYOa5BN1umE0TLzA4VOlilIus0HTUwTGv3Wm3N
wKtdUY8s91ZkmhukamXores7CZHnCSdr+J+qamq4wRTVfk11Ye8dLFIVgschhVYg4lsRAtZZPbtv
Q+QCnO70lRmJF5OxgKc4jJCtzu+PfCRoxn+CXyogVsLb4zVFFv9QR+22seN01HtHyHAW9UWo7CdA
yulxDrAnBgC+cKR2FNM9p4A3/PbudVAW2C+sXxSXYBYxBiBb0VIkRCSPNS9J6EldrnlFtC3y5wY8
BTgK6aUCLx9eCK5si5r95Pt55Dhu2Enc/oz1VgkdvYX//JP9v8o2rRN4Iw2n5EoJMpCcarVVsiyv
Q+i7VTbgQKCAztxIlo9G3jrxXqguBvEbtWUUGX3UIVvrcNFisZtl3qVsIY6R1dXIP0ET2VsnCyCL
RIFOSth3giF0LsbjvrCd4zjDwnaSBFU4zj3C4KaWWxiMPQktiv8R2teIctdA5FBxgaOuAD8YBX2f
vjpg6kW0NaOY0rmpClrZnKAIWxoIhD7N/KOQOl4wx9kjLeKex1eIqTDacM1qHVLJutcktzOoUZQ9
T19R3EEIigBOgI1ihEvOzN0XeQAa0jKyNu2E0TutynZhUZfQ0jcxVJaatsEzJM3ziIMG3f2fc8TJ
PXQYmd0Ea1v/DTawcKg1DccKWXL4/HIQijihHIuCHt6HsNOpN7AkuZtjB3oj9dYHj1NpF+bcsyms
5Rk5HnetzVEt4gqi+wF1q2cU3Ez3hlR5u3XcH8RVZi4HvOSpoU3riGNU00DvJfvm2E603nb6nJ0H
7szWdMoyuczsLAxIHglisTCHJ4j0hdY53yVqWEGuhGy1OJ3R31+ymdcRN5Z82IG6CKL/1o2Pu0EW
otb1IXPHcxdgR+Zz3eBLlT5FdPZAsDsu8yihr4mmhAMepGjYDujsZ+snwqcP/vEATH7T4KshI3WA
2FvqX4sx0DiVQZAAxecdLA6XYAotv6fn3J4tsMk7zfkkhY8O0twSmtVf3Wvu0UkSuY8H5IhTXXmG
u21JO4m96v/eYcbOKeBiXdknnx4UwSLMFB5IDtr6TcOOrn6874EkG7pt8U0Sx8lq85Sf95apQ4xR
HkE00rSaKsWpKbcqHzNLduDJmOu2tEcWA2ge8ZnYJrrBye7oYFFJdKYqTMUtt3Q2017NJUEoTHnt
JYXvPm0DiEoGFQL4C1UzqbLRvJ279OHpDz4R8z1MBrHJsf5WvnpgAhKML65AM1LzSSdovjRaj/7j
acuHHOyG+aUPKsfgNsIn/fP6YWFoBYHUjAA5k8MZAon02aaU8ygezkDbimhhcgGVVyKnMuXJfcge
rdPdcUilf2vXy6I77708yNjqHpdu6LTdhFazApMxZB6sIMyPoVIPxkDuoizqtMWc1HKEvUAv9hpY
tGc+II6bzLtfn8qJieIhmXI7ZWVk71EYB/b64mJHNzi2DE5spE9d71b9OaLR8FffGVvq38ezTreT
3/lEAYt52xEnZqOmCmzAZk0RrIY7Rhqt0tiI4Eptu+phpkC3j43/vBInXdx383GVkwQKIB3U/z3N
vSIbDHVb+8RHQrev+fmwozEU9vC+h/eu4yplGc1wyCN7kJAGhJQ/nXAy0T/ZEPbB8dY9WqEsLymf
aVAT/FTFgRwtzcAa1EfvqL1j7ixXqUHqdFj+t711w6PiijcIsJY1ZOBDar1C5LQU+DKUIE4qWAZ5
fWRnEupFJLl/iFM4B67LbQqtzqVjCuEFJbzABQ1ba6NsweWSPit1J+7/J2tGelwWDQoMeXSEyuWE
wj4E2+WfYQUg68fyyw7s3fy5JNMQ3MkZfxj3xyOnwOJ1nqzU+QkQsRBZ7VpVdHWHYUZxQmVysne2
oP1KiOTRs32nqVRJulhHILf8bcn2lFSvmqXwl1Wew0ycCrqkntxe7GRg4hmmkjwiGMOmh5BgC9fF
tHlmNb804ynvApsEi+vBMkUDr+uqSPCsVqgITSP2hXcrjsE3lVtD7I7Cr7XtTX3zXRYmA71szaoU
/eoimnbzknJFQD73lDoaitNua2Gk7LCr7hBLr2kc5sF6GmiHcj3mILvsi/KJselL3q+4ApR+A3NF
CtNY+PXSXOW7P9vZNNoEnKn9RQ83d+RhgORBbKWvnxxplr36BuPGaA4sFDtBW2CVDDKLFyCj7oaj
8FWlJ16HiNMYTZ3KCUk3iZbrdB0fOLKPqFCyFsn7UsABCpxifaxMYLEnpa74eiCNLLvKEIBcBFLS
S3EfpcdLNSEyiLCdYifWb62g4fYn+F3tOSVTYa8PgnhBZ7bMkmiURoBHlkzA4uuyXp0KWK4oYXEd
SSQ7l6vWfzsN49s1srqzauU50wkHKkigVN/a1OiLHIVaTDwtliI1fbMqE4G9atHMp7qdVHvPO0kV
ATVpGqy14W+l3xRO0PIwGGiv35DIJdoB4/Z7SR/4whIQjXyJNleZRJPbj6Dz2mAAZ4PnXwFgzlFw
ZtjcZedPn7CbpSj6TIu3JwmHp9BcTMOyS2Qr2uzAVdjhqOv671S048NwOES6gDE01VWIgpTu5R26
wVaqyObMdbpa84iMXe/BTMd8At3XWe1EorQraeUg8qKSrzYYmhkvxFo/H79SZVPa8tVmXl+btp5b
nP+6AnuyQ/D7tE0cLw66cIUJaDC16mCrTjtvwe5S533cUmWQwvd68mABJtWOvpmJdgB08Cuwq9LC
SWK+UpbRqfVmv3AkaVHyAvJyCy+kpVRl5J5gCL38G+zBO9C2Ii+YHIMIWLl4Eufn8p7X71Wxl1nb
hvGGHaidTkkuzhqj4dkTIrX+9Wl5puqIxd7mKe63liyUp+DAH+u6VYgvBDTbus3or9i/Vw2HE8Fj
jN7JjIuy0eXdy+FjsThRQdDcujt5hrk6C6XHcURZzmwjpPjpHOU+qsFuufYx3DCYZrx7uOUT5keV
v2EWm6o7UxMPrCXan95KNSc3LGeBSGo7l3s/QkTuRCm3JilelpiM8a4SAuFMT6aEddPoP7NEJ6Tf
DXBz7qc7h/1wM0V8Z3os72cw40Vx4wHvhpDmpDV2YOh4CtzUJoMNt0qrg5nsPAGJYBG3WazRb085
cxCMCIY6o38FBBM5NXaKhdY++Ej+ejr6UsOQobiKSX3OPLxgP8p8j5YD4Xa+Hz3FEnoiFTr/qqmg
/1o+YXtpk0iUSdjgZtmuaM9WoBICewgBTauVYCpEKNC9uG3pR7Aqr9f9vwDq09//EAX67CBlpoAD
HyFQWMNvB6IP+5oBe23+za6Vq9Xbb8kYlyqOaPNg7sVG9Gx2/rrerXCYOkAdIEysPzcoAMI3YZwo
O8Qj6YaZn9430cgxOfmOF8ACxAC130ZXIwUgq0PVBlKwvAD3aKpX3w3c4k9VLKKpHLbWpvjU5sj5
5BXFLS5/vnnQ298lDgLIqg1MkiIbZSxiffmP79PXcIZEcddAgqEDwglT6qXYaEMosSE+2FGxXj91
mWqlpSs434u64MjWLOVDQFYH1pVb28Z+0P1OGaCjfODDNE++Z9qRUZPifentzgYZvp0bblJ33/7y
6lKAkXRa/n4pnm5qJCpotDY/Jlycl8LY0Hy1GTHI4jL8I3/rN5pLUf2Ij2mBHTaAoYGhI4U5mjcQ
dD++ZW/oDC1xTXVNKgAy/jfM9hI7wKcw+o5IVZLW7FMj9iapKV2iGc/aUXuPx3W5uvEbflsltIJ1
JCXky1n3NMYt2Atk51RvTKLolrFZwh5yY8nFKn34pOrRnvFtqMDBemWY8rb0vmhqJeA0lhmEqxk/
XQPBSNtw8JIvAwNjhMmUGkzHhIWstlANIq+nC+19CNNqw3X22/bj7AurXjx8ak+gLKoQJFkC/q6I
HtPjrBgZxajnT0CjpXHZnp16RQ9CdfxpmiUvqu2hOouxQxbGc4aHEuPGrM6gUQydyZq3HwCWwmFD
OMpSSEUMnjPITA1YPOlqTy4/9QG/thV7KA8Q11F5eMQwVY0Xlm3Y6dnbKDjpMOSJxtAZFYP+udjh
rtShjfO329aAKW1y211MhUsUZPVaSKOwvCi6JHu7X2HjhAkUIPNtlPb6mhPbTMcxMqmVO5mFfs2N
sXmKI0w2E/xHedHzPRsXhXY2CTXxbYwxGDebQxnGCm4vmNo38SknyhP74DAHBG6JiGfm5/R9jZh4
ovSai0yEewyVN4zfCeOJAy4qHUTatw5oSjOlBUIfAKI7zZrlD3mEBdEUCyQUWsCESBydBVxOn1Z6
Ddog7RWyGnKysFOap8/kmLlr7aSe6xy/xqMucJ49k0LAWfiaF1Xz0+WLICESiB/uW2KyFg/9zHoI
50T5xFLWG9TmbOMMGLB1RwOwwNC64bbfBHEVi9zaBoF+FW1QOKSuUBwBF+1uwZgEql3jn1HfpfEH
I6NeFW4bZ4QWPyp2XxzZo1k3k+KY7Hg6zV+bTLMH7tLFjhYvLBRJMdah+3oJSX+lDzI83db7eC1/
KsXZzrc08vxdh+njUZ4lJLeBImue07KXrbCR8YARv2r5dgRh0cLHbltdzEa9fbJqiZl2YtkKePQw
kdoAlOIkfcjHIRdIfDd7+0LXf4MUucDxMUboaXfp0AgGowSJAskJMsWuDrzpbOYiPcjH2Qm/feri
pxab0whGjl8PYQtR45p3FVtWWt1pTJQPcPFCzN74/UdDohnJjG5nq29GHIkh7LuJwV3Sl262f8zD
WtuDQ4L7z9CoexB6U6VOIJIK7dwWb+YCpLW43RLRSR+G2Y+U52qls4cT5y6NPTnR1RSSapFfrIGl
KF97J4X3i/izY75yplNAee2KDanZcRl1Ngrmn/M9g7lFNDBiuZwBsuCT5W7R/2fRcxfEUZS1jrLC
SM9xLsIDA5uTb5tlqZYYKjfEdoZwyURT807n9AdYUN+8O0APUg35/wk6hgJ3MsUpvMw3eDx//BfU
7gN7Hy3P2FrAVXsDcZ/x8Q1nNbFyCY/uCf6XCzcEBQsQecA1F36sMnvRWQPSBKuHOV6ZIHryFd57
87ZrLm+yVwY1PA+bPpLX4VA4pwHKJngWN5ZUO/EMyifEhgIK+Md5TfCDxsnE27jTmc51jAp53ZLt
PZC1qLYsSJEzjkt/ed44WTN7KDgzMCaX2FgUpPJWZQdAl7iXz1euecxIR90J24DyHQ1LH5so1bXc
tOVNwxW3k0NHNiMzSQi9fYHSGGeatMRAzx/hdKBj5YEzoUrEADZHSLnJNW70Bedh+Dc9yuwKdVli
fNKHJ/+LWPeY204auvPiedLYYuDVmKnei+zzKc3AdFzBj/RtACcaAZ6Kv4noCL4KG+22Mw35MsfF
chCW1scXjw01X3kaCl7vEbUDqv+Kmey2zLle8GO3c0g5M5wZIJePIv3T2GqAfHKvsQkT/sYhMUMS
wTEWpF/hTelT3FekrsZqgNnVliK5/7emypGP37yDVwYF4N/ZZBxSoYYoZBwfIkRrISoymexkbW9C
zwvSbrEfcLQBh/gzzla/WhuRv0xy/kVVpw3dMqjEvW/PTlVUiLOCIH9uaBPEG/G2tETdJxhcif1i
e8wUcyd8jmqyXrTOH5a8AO/M0OScg6C8kcpWsU26ayYDLM+T9cQbPO5v1raGgAN7iWqFxuki5Dm6
1+qhAoey5up/3pGHdtEKR/wca1PIhzNkucpNGJPHG0JNqEk7YCXo3jpz1A8fDjCUoF4utVUGDGEM
2N35BlCNKDndH4Kz40xmVgz2W+K6QWiVEJLmmjNINl8iugU9T8HaF7peSRrg5aNpWz5jHJXOlYp+
tm8cyZvMoPw7/OgLA60dgzdrNwmmTNbfmi5wA6INMSMJVzYaoW7F6/MI5xHDPcIAebQkxFXhR1q3
zrpPi8JZS9W6FCkzW3wbDFcrlZRbuFLjakrMH9uJ+K0zn7rjVyJHV5ye9uGyRWL1KAG4W4Chl6nx
kHQc8uE+R+54w0PRJNsI9ODTINj+TCTALqyzlK69EfRbvhUoG5vxxQH573ea5OaPCfbIRUOSh+Y1
LoKXbm5UD6VUAuiYraNGMIejk1R6FrCRpK6FVJ8ww/dkZ2rtti3e0VKbmqgH/UCaN8ilAy/dI5v0
66TBRHBOyZi8CwLVjcvpkbnz0jKfAMV5nWW6gMtV/HVKgtT5IbgUDfVjhiUs276lMIYK7GqIjDJ3
5vbbgLYop2/eCHYnk4gl5NKe8cwjlelRGhcWmo9rKyqhO1pP+DbOHRz/TMIXbfV+6VYADfFP4oen
X854XBT39N3CgHXCvcZu3u/5CRxA3BYS8dDgc9zlZR845BJT3yYNUY2DBuy4bED0EV1qx09YryIT
CqSHeEi+bCs79A/yM9NmVNVJFTaNLiWHOhZ9n8SqSGlol4+iHpaMMnu8FU+HwmeK5l+bgadpw2ea
2CjqjN2cNONzi1h04dlkrbLioILa4LNFQeopLgqHY3vXGYqQXNY7dDo3iDIKIG4sYYUIQ19qKiir
cv35hhn+zbQhLZd8obeDmuDjOhCZJT6GuovbU62DIcQAiOA+PQMrvCSBK92Mb936EnwiUL3pFwNF
9mst9Ao8Svk7qHV86oDhD9vB/h2va2xR/NCas0wpPK1Dzz4WybQ4V/oBVRSicZETsDnKpH+IHV6u
rsvhxX8h4FdE4NrSgyFbtiXI+NgSCn5alFRONohWBmOipNtltXbPGdmZ1Gxwl/t3i1TpfOTwoy2i
45s0a9boUmxhjtEEi+NaFEzj1Up5ZmkzQoDRuOXk5f96Fm44gVuSOnnf+G0rN3DjNgWBqmKk4J+V
NjSViB15ocTEpiWvltn1owfO6+S7QTnr3yWiauCWr/3eY7jU7OiOpcPv7mEAaIkP4GY8NFnm5aWC
giOZTQonKcVK3EP8ByLObYWzDfBvuxHbeeBrI61t0rON1WKFFN+gKOndetntQMdR3+qLnHJaj9Xb
ZqGSVHRZpEceflR0+YTjQoXy1onsbD6ANFgUXO/NH18dUFCcIS4z01Ia4pcXC4fs4wbArTGpxJVV
eQxIXEfnPcPw/Rifc0vqcIS1BGNN6nq6wvDibqIlEytez4Tn/plkF/tp3Br+CuDcvXv3/eAKXpcJ
xsNKkoYZsqHQydKTG8y3NeqIKT2VeSzd+6VYPKRgUcMXUz1RhFzjd4XGv7n6oj4u+m2VUvGyQ4/k
2VzxHGy+kZfXLCS/5Qp0lLsZ23TM6QL/JeNTfVR/CI95UHrxaeKUgoyPGUAb+cvIAMlEz0IXNLvT
WY6h9nAz9BtNNsLoMTRXx21HtYyM/ktvk+qfKCl6zbSE+BVYRDXSTOEjDbnXtD30RQH600qVC0Vc
xOJbXWEPszI7Gpqrpa1dnE5y6lSgu8HbG/MJQtqFtxV0BM3j58BXkJwnnLGKDLeyOnoz6Fxuhhbd
1MqXcF4I3zApZTie7YB5GYznYoQhrDgTD9cO0os/A80hmKvkyIp3eOmKVFuG0ixSYlu65yXMAMVg
qPv0QWzPcNWbhT0mpgYhT/htRV2AkU6GFL1y29XpXfAqawzwKH5MROo3QIQwtqoVtgeUeio/uqIK
4tV6YPAswR7SA9v/NfAluoS7yQDH4JKP7MBGfMqAEexXtz0woYlKOSWmCve7gT0Oyd9tmAI1zATe
3A+JzQD+WeRyKqPLf95aErNlUuVrO4qPMY80ZnkCCPoyGzbTajriHucBMkiMCjwjF53/jWy/2QDX
/YIouiPNqrGrRC2aS8QiN6OTzUUtqbsxw8eZtVNcmBFrkP0QZi8NbxiSEWWIKlcwulbo4wPX/MaE
2qZGprbo7QsIQf170j2fIz9Kydmue05N/aRk9USNPN9DLxarVO8b/SJy2jRfE8SRZ/HgeO1/zHT+
g4a5+iF8bAbO9vAwzT402vTee9MCIUodhvGa7kw1hHK1yB50yk3nhDSmoMUhSEiWBUNpkbndGhe8
J8zFCuTAq5QR3SCyRIWqSV/zQoJXxZJxAWgOJs5kkfd7KT/9fCNz8VvynGFIYk2Bq9AP7liGlKti
eVBbcTJxQovonoJ4H4/BTirxN7qlKDa4tXEVQTQSxZqt08vkQ84Ylq9CFx4vU0xfEgxpFAxjOjyg
UE9RnKStcvQY8ZLad73HobBsjjxGtDiji5k90Hs64pw1Q6lw9YP+KIP2sd86jvazOrQfjkAznsKQ
pkgdM8P9x6HexJa8otF3/jFZ3lIR/zrmik7hWa+99fHuPi9EJwjfaQyBerR4CvB1uych/ZSrZMg9
S2UwxD6ew1SpcZD2OO19MTkruzzNOjPY7EB8gMq4nzQdhb8J5gJvLVTNEO39+mUcwPtAM6jyDBum
snBJd+xIEMdXyrIY57fgRFUCNUbK1kXAi9nf6hQ2xOB9cJ673yx6DwfOzNtueTCm3+dUl9BCNJfd
G3Mub9Xj6q+WWgDE7OcaPevjqHNMfQC3yomEN4A2vpZs2FC7yPXA5qpbi66WBQwCPZDvaoFPMGDm
rDvVeZbqc6NKXEXrLnz7PVbPyBa47es3BcW1RveMXVO1Ajlz6hNpR12iOmMe6lag/PlUgMEs20M4
iLKjL4BjfRiarchFRidAfsZmy7Yf8lzjV/RIOt8ivk/7uWxfbH9jHSxPeyZ0FMQvUTGkTW+SMNei
AsAwGXvRQuUgCxqwEGKofuXAwIRJhn9UA5bwDzGP8bDOoH0sDh5UqKDTjbh56srXdJhn08CzFslJ
Nq7Y+fj8BX9lURVqMCSLUTuigmAFCwgs+HCMiXc5/e4+yl1Hf+d45+0vQ1P1j4vPvQFIMXrt5aGc
qA9PbG+v9edkTCHrI0MPjzbcYZ+6WE5NCa1XPJbgTN/ggTTUGGCwapsG6clDSNRlV1YSc8CsTsE+
yAWB7HicMVumPpOoA4Yuk9xMSyoQnnTQNBpSeHW4M5Hsss/7DGRc+BHlYHGb7x1p3R8+TK7uuE8k
7yXm7v3LBOby+HjVaiGC+Sz0TVcyR6IRraTZREDhTqKmfVWLO5wik79XDAe/W3J+I5pOOZb2/eck
P4FJ4gydGFVpiRbOz6tgJvZysaOQilBdASjHuwuaEGQ1SwIAhcf3WWRaPFXAp8xj6yqpN7asTo5n
ljRiYudF2jMvxbFLuvaHoKLsJkXkJbT30ZoYkmueyD+TnjbRIVfXk+DyMraomt9W5iOLgLSC5sRH
xXKBTFaprvyj3vJuJCoiD+kXno/GLEBnP8obbRetNwTDegJ5N0Mfo5x3CaW6rkFXiGCGyZbnA3vy
jb48sxhRs8U9JqtcWEfFi+Ggsn1wRpdrVErXMDdP2ejgLvwPUNfP2rloniZycoiFnzVEoi39f8NK
zJwtly4lUaYRDAUnSI22bpo9rC5ZC3BpCGkHG/knNRGnz55GPd0Mdb/AEx1r90eM5w6p4n5ziMQv
8LYfVzeZT62lEyVhMvMdRKjjFcuGZy7Udxwep92hWL3xU8KpbsC6Z8V/te86t+AChoKDjfXJzCTf
7Jsme7xH1umm//4r8ORD3TSrfNRvvGNJ+iMI3QIJaY3oGkRhCJ3P7ztOiMiUmq/+CScTD+Gg4kpv
QHuDz8jgB3RdlqNOnKdM5YPyRZDpggZmsH0Nhzma1hoz9AkFirb7pp3mnM7SvYwgUVydKew78gnQ
IjaHlEnSojdV9GO45aAnFYq2gH0emK9F2SWajNGE5oW4Tp96Lk1CsATDcwtxW8EKIKJ0lMBfqMwL
MxuaidFyJy+x2dNoofWKCf9lLF7lGvBZ9rh7CTomjCcWXCGHF85W1IPBN5ySBh3gtJHpy1aOHPFh
bpPn6rOjcPAANYRhkAHNq9dpVYMVAHuvX0gsyEcq8wl55OSJj/OCzV3WZ0yD3qEvOX62Rtgv/bgt
DQ/R8lfxogfi1dbqisEvvnUhKVPXrTAS/eJ+FYS3gZb+JWh2ALrKHspMwU/cJ3Sx1PUPuiZOb0U0
9wKhflon6J71cvMQjWoCFuCN+cqfZsEhfWwmATGiurWg3EpPzXq/WtysgzEb+d4+/i4djyYKppup
MO0bm8SS3fYZUz8V0NjTUvX0+CExszJOu7T+0FpvGFyB3Vca/qbj8ichXWmqdU9Y/bf8yn5O0RHH
5GsKzwf6YcqXferxwOe9AtFyYLhD/H8eCDaAIVbmLJUqNGP7UhWVkIFu6Ejy+UOf2zYkdtUmXkLB
lM9r4yA3GOdmwowisw1JZFW1VwmAAjBGnWr/EDT+e5nnEOIPryiRQQcyv9/VtlqbEJxo3K9nwPDd
8EPa0qdE3ep0KOIk+BmzgM3SbnkUmvxiqaumIq2VfeCm8/oMDOW10QHu8Yi4RytdzadNq7eaKC9x
MMDsNodzfgIhcptUS7yn2PASSPujLEK0FY9Ls2VlZVt7qHQfiJ0YxeWeySikGDx3oG4y+yXDMSRo
7kjiOoy9mLyBPz/06bBqZRfkiEX4zvcqUesleo7Yi2rZesd37TL/mgUMRu+umHxgcECPR3fMfjuZ
4JRDeuskWxsPOI9cSYfe29h42508BMWFK6M0Lbgu3H+u7oZ8sWdrCrk62P3Dy6dELZGcCGTDeYT5
XC3l2HKrq/CCG8h4nRuEEmuugL1RD6Pfw65ZdvYhelA/BOmZq/jQp6DUFH/JkQ4GvZEV+qChApn4
3CcGPGySsDfJ4zRJK0XrDLezEL1Xyhz/6T9tBmtNAR+bzCAphQUw8SlW570j2iVQH4Gu9MdWH0PW
OKHGoSwMITwsFjs1TJuBH15ybJGCxBApuID2ewM6VvQVzAfuq8Dfb5vFRFUnWej4ObSZaVBL72E/
pdKJpk+u8QSfPdtalHdQJPY5HRYcv8zdQI03Z2CMyK+MhL9pLPvVqZ2kimP40vCqLldquEJlJZ4N
typhAc6F6OO52JMEtJYUAE0fJ/j3PiFFTedUjxw4qnEnrmnguVKQ2kDq4AEmZGWYhkppWVSShQ0l
yoH0rddNpO3m/sW9e34fi6xA1rA+czX0dvpyFLEGcYYLRYepWOOJbVjURNVG9m/XWJ3ROfv+tvms
kB5XCxc7kIU1mg8055ZhpZUn1M97Ae0B/0QmaBB/sJKxPKUsPZmEtLzQSKyTdUqbP2h3/cMeNLZB
coEDGsh4YVVR8DWhuW4qD9N4Kdk56hgHydHpkprr2WBXgcspWTyPVaq2+iy2EgAYjPsa8zZrkFuz
qHHIwElhE3NOlaynBbj05yqgfjVUvPDlo6PxwyPyoAzCPtjaGbN/jaYuOyuTMFYSNk8DduxBrbrE
zyI6BuM2ECuFI36F2+thcnMGZx3rR05nkM4DYxSmL1nF6isZ7rIOlLwHg80A8xpDxl9MK572gBaR
DA/NGdgmWaC+SZDjLdhEuTB+pyR57o5YvxxLYwFkmuigeyFLurVfbhWddfp0OoJld8FkPQNDoa2E
mV3coAfev9I7Isioqbu02R1KHiV4psuIaCLWcnmBAIjgg9HaG8WynoZbb8YnB1OTPurPzpKEiQN2
kO3Ky49CmoKGXoV5cyRkrV9qAjFodSvLAADVPoOOlMJpvdzPHQs9NGz1JyCgORjROusb4Kerwcf/
ZaFc6LpdZZ3uuzOgPQP7lRfjz0JWY7KXNqQsWLjeO/w1C0cbIaEjNGj/MfkOPnueuss89vpebwC0
5jzphyQVQhDWLJbwmnXIa9u4jl3GPFfxFCN3UI9XeIsp4QbZYYl+C82vyn/GBxqpxFNEa59SC9Zb
682saYqD65sRH+7MzFDVc/rviK7ycfluqgTqid8de2kHbcrvubV+HECyQ9raukg0P/QtjGzVeEyv
nPqea7fXjMUas1LKwt55K7myMihgHvaXrb9Flp73yxkR56UC5LrCv3jjkM5PBJJcvuV6IDlnNp3i
liY4ntb/iBCG0dqs8DdM78x4WnzPQpvGxWkZEvJr+0GueweymXXykdcN3e4KXHb1SQJD/byk4LUP
V19ADy6j6faejkhXnqllCr+K8Rqk6EdvYHbYa7/oo5gFRRTb/eocRVo36nCEgl6Id3eAAxIH5TmY
ZhwYcRUoQj1jlCwQj6pwyEp1iy3hLTt3WxgZW6YR/S/B9E2HqStwgqDTh+UcKdz11F6sk/g7tBhP
7irIZ4WUvK8/uoYFE8cAvfCSq3Sfy1p+zkw20NK4ADjWxfBGO5gvB8JbqL8h5TWRyAJTJDtlyydn
KHlvaOu3QplLFWuUxMZJe1rGAEzDvxU/0+Q/u7SyRwn2nt47K7K+sQIr6D5cKatBRwBn0MIhC5Ty
Jg6eTilR98GmKr/LUaj+8o0Y87PlUAgVlcbcCgmMMNr6RWWS78YTVPJBQcPl+ZByfoQiTlrFf21F
WdaY4cBTFJmFqNEnZwBJR+rUnW2CwHxviX2aEnJpCBRhi8aiVr9MQPyE8BuL2NmIh0zeQ1qtF1k8
SHVm+YI68xc+pBNX7YFfxj8cEoM+U+Nbho5ptEPAzcPtgoCKx5yHmb6MUG3AXOtmaI+ENpEAXrtO
akwfNt79yVU6/WoWN1Z42NqpuTuSLFIh57uHIzcyc+Upm6EsvBe+p7IqoUHkOeRQuHdncpScnynl
A3KSxAjLHz86GPkcxYx81uWP53fXqXT+1LLP4R4XqCmZ1E+MbUaN2q/0f6LZsSEl29Y9QJZMHSoC
fDLL5rTTyvLx/hnrD+x0gmid1XXN1c5M3EP5oDNlC3Ge9dl0F2CNOx2EnLEUpteonn8WyfMpWPlY
MDMpcKpHLJklw83t3M4nZvAXfieUYyypCF7vRIZxJTVpn2Wcbz+N/bfefOlunLVqu+QEpaBq6lOJ
4AUHkPIuCbPABjFx9Cr6C3QlUYBzC0m+jqssUEnzwTP2ZST7he/rpypuGQUVCQHuAEdr7zTvLVys
6vkyi6KywMt/iNMXWbxz8PVhekfjX6wXHq5EA+TWeFsaDpktiQBaUp99GUcitKDatjXR+DaMdAS1
eWRGnndGiOujmMQOGH4QZstYJy3a8e6f1AJQsUWaMT5ML0WrPvdnest3a7KVEIC3+CeLgJfSFKm8
tp9zh5heZrXBYSTbnf+7jBY/QRQkrvi9XJIGPRZ54GzPEN/lQGsJH2eB8O8IDGYMV+xMVcS05/DM
LdnYknsYjdWWEkGi8lbRaBj8Yi+g8QVqaQeuReXhZh0zGzwJ6MDlvrNe6AokEQ4VYn2mYqlw2enD
13eG7GKk+XIhNdEbe0ZduaSXTWt1ifKDKl4eG6g8DwnL4NAaPNzOHqIYIYwOw+Dm5n5+hNDe/eFi
mecmj6U0jybdNvcohly0DvOXVQHt35V7O2Y3tUAEWNqd9WtMi+hxd0PnurJevDGaak4aPXrwSC/N
60xN5GUvgQO2RZ4mxNI2fDFtLrbQHkMndSl2E00xbMkCxpsKgGK9u8TCVs7EDQuhA/F7geYktwuC
WiAPJYucpurW+w4Pp4wVxDHeFc/4OGVacNzZ7moQg+5iVaC9Ea5AERI5FHXWp2luKBk0ZBfNRvz5
xOm085uQHK/2JBoTyhZVLkm8Jun4Dedic6wdEGJs4Kb6sMaxqQ6b8Q4cwVhbaHtqWx2Ug63iprbe
p6g/YBW52ZtWaIYub3RZJesT4a+AwhrNKgGru+w1wC71RPDGt62UlF9iI6FUC5P272nXQGlbJAWj
6DMG4zA7vicFOXLfhhYC0dO/XkejzFp5+MgzIt6Anb5GcEpAbsccFL2h6zsB9W0gO3mzPi6uLJBX
B7X2XUgOHwIp33fN2p60j+vtoOED0Bi264b6jeLDnW44JAzlZFZiUVo0U+lgyFRtoMh6+CkVGhn7
GzxQLYy0yTegqcAGSG+rpM5gyyMNg50/Roeew2OOXDMTbPz1Cn3XWCfoEBPLi7O86iMjxI5IajGD
xyVBPfd/NA9mtF7JvWifxCY+u/QQjl+RYwp7CJNrqjWn9l5MwpHsfPAJSStZM+81/R+XOCz02umG
qrjmBjLqfFcSGMt2kleP3gH1PtKHIx6ZmP/yvJCJUfHD/zNCldF0idgg2DIW3NBfYO/ctDfwOg+H
DUzrf0UqChG5sjdUiiHLQwqUCFo/Z0HVyvDFXJakB7YiWbXL/s7E1Qt28dnIzHbe6hSQ7HVl2d+q
niJlFjh6jGv10EKxr2WyMUqwW3sicUFZnpVtbzJJLKNTvUE15Jhd0nj1IxpEA8bD88O2TOrOUWAD
9HopAlC2EKDPOonLfuhqQclRxO/toXeh/r9la7NOM0Pv/uPCzB/2fgnqRs4/7S/e9kh3tN8y39PO
h9ZVWd/1C/6Vq0iGNVsIL7aLxEKWSn/wxn8oXAD74JXMyW9DUpKNGaux2ZKEfTwwDOxmDbX9Tp+D
neYYoxpztu7lJhaac52xav0eLXlMd5VPs55jPRU+p98X2HH10ifR9NWJvyEn5axr7DVn44vBuTBV
MAy/9CBglNL3cVVhgtIWT21PNn+yGcvIJQpEonrd+OeNcv4kHcceCPJFpKlU7Kwi6+/yJ3964JeV
L2Tv4dWod+yy41ZjDybUQJKwnL47z+ZNQQmR67fU52TabT24i7byRHIDBQYYQ7kPX2072kWiokxJ
CY9LVv8d3otE+l+Vb/xc03/S3mEufUEx63hnRz2MpynNXI/yghVQHQAuYLvMgFDYIZeua8k5gjmf
I23BE2fToQgb9XEMOfTWZ3l+GXNDZuIjIgWBsz9Vb/jnO4c+kPvYNuOMgy7DYtpuPHsu5xW0DMoT
+qCSDWn2rCmsUztmvX9bgdBrW8lhPPGBSYW1W9AX2D9sC85F4+TOS68/A+1+AJd76wgXyBjLI1PT
S3eyE+wrmft5ICw/XxIQT68cojNWtZZkhMbi0k5r6faimlOIV607fKmv3CqR/rc2pVQMhaY1uH1f
i5iT6qrVZlLrPcyRR2Wb2Eu/1JVB1rCPDnjmNtN1qYqwv6u3uzyDPthKTW69nvRmfhl1ZQYMT9Sq
Bp2Iuk1Gw2Pl7vTVbiwfxwjkjKhO9GH0SWU//Mj1+XB/sZH2XAXbHFMj39H17bN4nmkJtSmsUbz7
NgEjDFiBLV25/fG1zmTKHhc4GGgfnUGMAVCQp3+Wi2YumV64Ljmwh767nxe6fIUecrZR7m9KlC7j
t0hWWv89+uJ8Yf/20VXh8gGv7oEEu8YmA4VG27pUsrhVT+OxdvbjQwXb0//cEbaWX2pm746z2KHd
XffkQS2NXiUF4xnrBj9aC5+s0dP1/a0aaVYpSdRvhB3fAMP9AGLUMHmLFiTLS8vqIM23sg4pIp3+
8+icf6RKheYY3D6+18nopdofx/N6599+mEeAzQoZq4R+GtnjKEbEwhALsujeyBmtkmykzrh98Xm+
uxl6zAmZScDvZxP761QmpSe6cIj3iQtBsqx4jOBXPDDfaMnXKP3CSr9HQG/42ZLqFSVcNmozaOXH
RvNQqT649t8ad4/nSrjfy6s+QvCoDfmd0IRafBlKyBkrQUwdCSdJ0xUlLIZ2zTO0bozx0104l8e+
tWbvuHsuoFAdYiVXihOjWAPhhqurF/spJctKuzwPwg0jRRI9abc+WHCdq2QqVruhzLS5WUi2/tsI
bO/iar8yG36pAojGaecywqYOI1oFeU/ixz7HO6Y8xjimlMobw5sdu20QVKXSaCL9aXo8SVztmUjm
ATDTHFv2qmKgYTs/KVOtHTvVBzr3jm3Mb+6hqVQU48J/3IMXulSp+mYSP6z2XpuXDPjqVy8Fk+Fr
hvGztyYXAUDStkn2mver57Mop/7QN86tuO4XQsPdWNK9ZjAmateMcu/nPDByb1CSKZKClVXC4gqu
swNsLfHZJQtVYSAI59au1E0+CK8ZLTWeI7ZYMXLqw843yMOiGJeF8K2bgt62t66WxC0TTVrs+PS+
09RF3sazXLrXZMomwV2x7E8a/DSS1KfYXAzQfmkfuV71evpdrFg9duFvE9JCdF3LIhjZHKk3NZhq
PvnesQwhjVjicsyA6hZAyfhxcmnTJJnl1vhIfa9o1kmcn1xX2wz/GCx6eb0t59we0+tI7ckJfAor
MV0deDZ8f1Lmwdyrm/yxx2M3zJ6SBcyOBWdyRcZjGiQTWrbHXl3Wa8IfIT2k1hJNAXqUQtuHVvTa
BRnfQbq4oQMDVJlZCS6SERzV4xPUmhNNf40icUwpDSx4iwNcOkgrwbDvgr5gVdDQgOEyWEpf3yUH
+EhVh4zR5V9eSJKQaGZ8ku+2UAkoVsWFmwe0WWev07cEiNjAqE4GzFnRSxgPtmw7htjH2N4bGUIc
sYaNYo3nJMc6T5GQ4OIRI4gwyZt1f+OkUvW1KNCspAYNF/gPdu63GFga7Dgk2wa5UjZhSiF3oGOI
n1zowF56RtsvNs7YdeyhXzWslvXBD4IoEmR1GL0R8VSuKHHqYxhTytSEeZfXdTE0Ee7FgCNjXBdn
jzPljT2Xeg1joptjIYHv6kJLMPtzu1b5Ns5oYzuKJv/bo/mMfbjkWxpq2vR4WxD+z7K0uiCOBASX
s6/X/Kb0mbD9TWsY4RqXp/Vv8kKfBxJYOxSjuMlDtZOvdiX8Gqh/vSJONy7pzS88JMvhKbZt36Am
7giBeTF0kDNLo9egTCaYTS/vJ4DuefKJVG8zcXrd7s50/UDFExuGyENy7FAJLLzh8mOHEBxRCQ93
3vVgqteAw+7Q1xFgQnblcUd5IZxnBT34VLDxJ80b9Sh9EjEcnzhvQnVbVev2bwj6wwt+GmSBMZ5V
hKbkm1AgP8/Ii8StDQj5u/+eLNcKMt2sQoOUezTnX5lDmFHg/PIwd77SlA799ITaxZehH+ApEyMl
TpPfHIBzaYnXqijWR6P9/PyYFpgm3scqSI17BoGESoTAEIej63VdZnxn7/bFUjWEM+9HQHZAYO8F
ygkKAPoMNsdcAvSDs956UVahqoXYuiSk1pH6Sbg26e6GhvOgVb7n2s02Innrno1nlJo0F/c3wXPq
dht7TUplcLbDKDzJ2+6pgTcsEEXDDgHC0XQPgbxm+eR8+3ihPVr9cYES0aAP8OZEg9qR59J6Y1M2
Efq65w+q5eUgnyB/Fw02ykMOzbsS3l84iqC6Gbkw7BleXfPVO4QdL/IWsNMXdYHa+VHeQJOndKfQ
RnytCyDHXsfbRWlAvlwwnTfuHxlhBGRK1p58yTmweTHGnCkjwW3BhBU9qt6U20qe2Lr/j7IFBVtp
ITq9KyllNuejZJS3I0Jir36OGKC3oO0OWHKINdbfv2zofVIFWIDySHnHtQ/0vR+39me89zE0W6KQ
RY0rgDpceIqo1YrD/r0iPqZaRGQpB2tbFxTz0d2iXeFPant3sitjAh176Ds1xSXMmzQPkoDctfyJ
w/WoXQOCWo0i8R/gzv9v3kgfWDBBgwKz/yKF8tO7EhMj4H3yDZOrBVs7iPlTziEmxpTGR3DEmrGP
ZCrsWSuUPmuujWQstsoxg4YnZeaCwGl691Z80ZKXy0OiAuWmLTG+IDxHvc6KNZHAsNMvcBJ3gZlU
Ruv3XyBJ1RhyI5sYOwX/1Vkv336FteFBYi2ym1IZe4JuQeI2sffe3+6aLsZDmP8mX9DRn7HxhZSi
bFKpXr+GPMQRT2yOWubJIkekZLbMfGVKdjzrllUt5STRZPcjPS6kgChqoaOlQQXodAaAR0dxj3Dk
xxvGNhpZPutvVz1Rg+Iog3y87+nUoDueXE/W16Kx+DuLFBTCnP7f2GFneZmI8oA6+GSBgNMrYXrO
vTs6KzNBuRX9G8tGq6gdAWf790TSI7369jMeAxhsU3e/OdSN4deenMJA/5HPjEHVRR0c6+csNQX0
DfIGqyAbA6BIcIxoXAUkySmHy8RsMtVRaGHsKWpK1EKKmpKqbhEPc/wvzq6Br+gGm7khYwQbrp1m
p0ZVR2Z0Ub+cmqz+zsy0XQwoPbYRTQdWYr4xLUwg2PK15Q0RYJfy4nJ1yycX2ku8hsZl+EhPYDv8
mWb6r+BjCMKld5GnYDl/L/DwAkMh/EixN0fB5F408GJ7/13aFjRmxDOAez69DtV0WAtAxXUdP5aa
m3JbdpjRUf2rlYLRbC9KpZ0iF3411lkUfE43jDE2jHg63CSHqiUdMAufzLwhsjZWugxVljFxCSR1
kILaoulMknlYPM3LiMtzOi+fXlmP4WBrtrPDlN06Ewr7OB3hX4CjR36iNZJlmk3wHEd60Puhp18+
caVgfBlC4ZzW/GojzAwSBlrwxwoKzt5hC943Bc6W14bs7P6mWse/qvXh/VjXMdy+qU3jDX84E2u5
S+Wi1B4cQD0lMessF1FZBiA3IWkD4YzOzVRYWV8pCf/EQwRyfy/2FNiRcIU12vq/p/uOLeJTLWy6
VVrOsGCw4Qv6VULOm8t+I5zsYkXhZ7CwOWdjFl6UJ8qskDE8z+UIpwpwyE0c7KaIQSi4JN5CHRkY
LpYKlaNVU7HRiMSB9ENnixaGEl1+plxR0eYjLIs+qED7107yF2+yoXt/1L8NdMGNrG8I2SuGyUd1
Xqp+69usE7mfQbLajvyM4Ypn1vjci0hszjBPRCXxwKCiIOsNhB/wCi6fx4zp9/kTsz0W0DBJVnmO
AZeQGKY9HzJAO3jPCCAofR39VTiDXLlDTYs0WsDR1MO5wrRvhH6QTgRx7dorHRn0PczGiZYecl0O
6O0tWudr1Bsf6pYJlVrSNheWislajpzAY36eQsz3jlCNKyBGfHS/Ts9cLYwhw7ilT2ouZUMX87lX
GTx7Nkglh2ZkE2VFymbOoLcy66wjWf6J6FJTOdVsGvJXVvNVR9BkmUta5fit1jG0TMx98GGTVVRi
4XAB7/uNhZHYXi0ypnsiw4T+yNugYBWoA9edgdUy5bmg8eD5PglQcz46OzY6qIXQKX3aG3JmdEoA
m/A4MBcDIE3g0SE/5W+zdq9/AusYX9Jv1qmKJ1beeFkse/ukvI8D288XoqYQ6Qnq6jGUeU9CwsUk
nvazou/OvpvuS88+tq94qzNjRLa4jso4Iza+hlFzhjvsFsZVCRm2WRi/M0EnGD+2ow8AZC2of/T4
6FDTcPiQDAUA0Eo1sE5MX2zlvZaxR9x4HYKOXX06DXMVesIeyQXr6N5v6/OJzQcYBYEXSSlyRBW3
upepP+e9KFwXPS0H6T7N0XEeMaYOoT/4W/iuJdZ8oCqytid9hIQGfLN8ZFcIZsJqsbCqNaWByY2B
xdMTC8u9Yl2AHP8Z+nMFsMm4sgUWnrEiots+R4iu9IzfgFdvbOYr2KE6r88d1jdXcKdljfFZUYbM
w+BqwGzUYMy0QM3gVeVXBnTDmSllRg0b1lJcZHhjGjI7O0O4+JMeR20nHe7EczOHyWJpbBrmitBE
AwzBXeUI2JNG0e2pvoRJQJPh4Qjq+nlqRRqA0tS+B/YxRut2Z8ItGdBhM3VrL5kgV6kC6eWCDFVw
t1XomZRMp59AgQKtUvR0agH9kOy1nXK0vMJQ6eL99prIRu9Lr6eX96zv8Elff+/EWbvLoZrPgqvw
6z95B6KR+eQDqdbD2VvWcwuvdT/gSAjLR+JJpObY2kqGfW9XFfVNsPg5/BjzYzNijRd1dcSDk6A7
DxFhSQQrwBfgkJSqwgxHXb3gDpToXl6uY+4V/9jt7ZSCvWt4eoMaiJ4zcjrcXXllUTQrp38cGvH1
a31rs8kxYmQvmEhiv0K4HQRJ07imdHoBuELYhga8VDFG8vnviNabsULjE5i3yidtXcIAscpXrpnb
8J4iGXbJaITd/XIvvM2QHc2dxxjxl7xq7xFKJlxrYwPBxKpAS8fcUjpYPctG5ZWnSRu5QY78twLC
aJuJelrPUm+ZR5CA3Cfk3lX4S7vRXFS+ybWC9WN1aP0nYRsKLaetrJJxRbl3+q8GeevooTlyT45H
PImqr1PJKbG2LCLpsfdxN063uI0FUwz3C/tI35STZJUJaZmQ6P169ttG8ZflEA4AmRXfxdrDiqIp
0LdemKGsuGEH8Q74Bzxc0geUENQq7phXR7xdSDRv34rIWQ9Vw1CHIrBN0XH/v7ceVb47K4Dr4sUI
OfduHBRYc9gypFh9+Gf+ZT+Sksljkx25O/IyMHILFXzu1wS9WTSTwXqJVMqlUvVrqdD60cOq4jM4
6VuW1jIyatmI0wC4WwnRgD+knmagyKyBhANtQQpYLMp2yBowhZ1cbRIBYNtjAM3bVctaOc4LO+wu
bwi9twidoZ9fYqkn5AOLLqov++2UnHout6EcaIv8dhavqYsbnA0cwmM/FvWau011vdLaMGFAeO7X
cjUuJUm30FYJi/tl3bV5iBqrshyNsfhvOLvdS9C4/VVLJx9rHa4dAMqAIOdCUGRueTRwyodcBnPP
2LqM9+bD/XjY4n1bfEzWT2HH+FBlM6vr29y/HPLIRSaWX4zhaUjqGiu8NNy6h5sey0+MtO1rnW2T
IOoINL9tuS4MvslHXLHJMTkEEvi0DNeKRQ/9X2IrYxcKDdVTDjXzzWS9jpUOq8hSZsvgSOxqTjoB
r4k+643AVhKUpOgeQembTnje1OWcJTS02oKYtbP3EXMXivqfY9FgYWcvdi9OZCLgIfDKU5AaB7WU
NlT81ir02NH8xw2z4SIx6hAwadZeyTVpfHcu1B31LVRCZz35U/yyjxY218kjdPXy335mCb0hgETn
r+uqt7a4OZxdup750d8JfkEOJ8BhRyiQbc/z69jAtcApxs1OCEfWY36MsbSN3COPyMdK2cF1OHsp
YkZGE7xC8t05VxwzVoS1wEAnWzyFSNgBDZ5o0gpuyYxfSxDCuKgvCW2EuY8zKnCTy8xXuNv9FawI
3MAi1ms2J5kthu9HdjnZMAwcwokM+99OWH4w6sx6hLkNadK5+JlugQRL164qoaGu2O9qu+EbntCR
hnHcJyD6O8OdbLvMo0RgHe7rpHiUEkdFAX47d/jry6MbdwZkjDFCZ06ZkybPdiMowclD1oyq/Zn7
2imxOWAIKZ6/jyxUiFlyNvkKvC/cImiFoN0a11O2hWBpKqP3cUQTfIBcUtgfkB1HX52jJsVnUtv9
kWHjZSGdDfjW6/Vd84BEh7bf/qT9E8QS0LFV2ZdOyZIO/ul62gxOo+W2DiZH14kU1+0SdtgRMKeP
TPilT2aQOuqF742LdILZTeVerDEXEVfn8SHtR5WouHEMC//KJpRBcI9aDuPfvlSAYxqr2/fWlgH5
ff6DjwrpaVL5GwY7hZNrK467xBED6mRlQA9E+mKVBsl4SjclV41NQspZ8mR3t0yN8lwLPdKP1hgY
3XZ5nnP+DdfBMrOKB4Ys+BADAKfM4j2Nt3xOCQCLGZ0kxO39pnATHqomQgQFgWDOCmgVqMGp94as
N6IU1Wtbg47guXYGc9iqHiD4n0r4pdNCV5H0xX4FVrqGUlu0Nq3LB1NqAc4CpGQaX5H9XLjoFED1
HvpunfMp05/k3ehkZKb5uaysWavAnUFl2i+/R6WJluhHGWVyi/lcBEoTb7v/ri6duTccw7S4bm6c
Koq1KSigcse+kppQTkCfv2QBCzNyOEfaOh/p+itAJxRGDGmXsVgRlPIw3CCl/gDhqTj6p9onM3ri
Ttnmrdp1pAqPfDb+16NQx6pqsw4NhP6JRuwRS9Rizt1Lbgy7PfbgGImlmtaKu/UX7BDbmZDV+Hda
y1S4UPw+QhY7kHRZ2V4FYM4/4/pA5xc3fY4sxDE8b9wwOSuC6aqrdVwOxhXS3sdVBuLTfIH6OT1E
8ZkVJenb2JGYYaAJTz43Wleb2u36KCDTjyIGlDKOMUs0VsNNPc4PxjpO46tZg9dfUSJGZGvpB8MA
kdqJEMbc+BXA6Y/oExkw8wrqx9INYwNPkTAPh0EL6fVePsC1qMUKx1EIaLRwa+o3SHCnegeiZlG0
vo2Mey2EqQ9G/lN4x6aTwP+0Rv9hCqvZpha0b9y/hIoTRFuNE7RCWbg7wCaKtzA2tjmugv2W0Kng
0C92mAkVjOfy41sJdE2FSh3TIK+JmVX8TQAQ3xh2QIpIsK504TThFeyX6YuZPx4mW1qjMIbJY0xo
vtCSxnstcbsIvXKOvM0EDBB9E7JccR7ScQ4kZI1VCn5reMuRISq08EU2W1N6+Tsr1SRcI5yeSChC
8TI6gX0up7OAJYloYTjsAk+LswOWKCgI2EEZERcTwUUAoguWUYutAv56VdtIwgocB8qY4716iirj
Pd1nfZ0mWF/WosyY9hR/A2fhLdDydeAP4PXPVmAN/5RII1vbWYd9d0xZaPG3cvqkxIgQIVNFpgW+
IPu502izWYaKdu5vXHfNBHfCrMDTODRDtAg3Azowmn6Ex6cK43Z9HTBJ5xtfg7aU64z/g82wSJha
rUUZ1jxOax+yITk4+2racG0lPA5fZiHBvTPcS1WppCZ/kMpIbDbs9tO+DRp3AtSaGNjIJJ2o+Sei
6GjObplrJYOLBWtYKzWKadat6B4ZlSL0+9/sLtS56X5t7LDOAzWHn5rvynpYmyOumiDUVfE1otLu
xq0DsV3lvlyD2izYcrhkpOR6QV2mSTEwyJ1kISxmL/VXU9gtysphxFV3UCuAkRYwwWjCNT9IlRCo
UK5MS2lPuklo3lx6zyCTOMA9Fz6mB4x4ptpWKRmnppZqjVp/O+I9KpfZwlSa6T9PJ9Pdp4t5BarN
3USYTr9D83mIAk3DQrJpdEvfDmVv037FNk/WG4sFGq9AyHmNaJ6vTQSBep2KRyjcXcBifp/l9p0K
0YPF6ZWWNW97tpGzYyVeJg7Iyi0lHZtGR2PGu6Xl0GkjYUJdm+ZW/a1liQTQBa7sF9iQpIdadH5h
bhGNB5+sRsCfwJkVX3G525moWTFgK2oSjHLn7woaW68ncfbhlRWG2bWZjs/lFe/YiOZ66b8zuAnZ
EHKHIYVmp+3jgZytNn7GwLiaXvUi7N3NDqCmkXwr0WModTVQfkysaYVqslJc6rDOqi/ZhII9/ssY
Uo8SGfv0RxXO0+TOb6orsGXcFLezDAqGhF/w5wVwc382utoxQ2bSU/PoXGDGbCxjO/Vw1uvT702l
slGkpRDy/b/5s96hS49qQSY8UqMfEHKft6qFPISq82mdYh/rFMkbDiFF+fpRi7mNtN7hoNcLS2mP
vQ0mG4GJM4fH+hQAu9TRNhtnqTso8damd/NIPygUBxfnCDK9zsXsc+iV3ZfQbR4XB73sq17ojS4X
WZMU89gf9EW/G7oGz2j6Cyc4JmwhB7RfL4X5314355saTkWgf9+KkFEYDruh++AYAdNY7z9uNxYn
NIaq/ReW7rFJE5o4j76Un4oy6t3dBZPkJU3nnK+rIa4ezEIzP/UZ0fNEdaQmB+/wJHT6dV2qkCAy
cKGwRyRgMY6RE0P6cs2DV2+5Ua9feND4ZL1IFaafp3B8hdS0lrTc4zNFbCw3BibbqBAAUHqH1ZuV
l+BnT4fn6Zxp09XulZx5/ZZNhNcRvEUz2I/uALRRQGfC7SeA/Jr0cKD5eVbxfAYdEFfDEIAnUnKB
9AHlVJ9WpXgKa3dqAgVa0iKeV18XqI9KtOr/8toQ8aIZF3UTRHHLYzuJfeCuJygLSUgdgenyK2Hu
vPoH/cq9hUetVEChb89wX8uk1ZRVrcGur5Ywl1wM4RFMwvA1iO6rbjiw3NVM9seZbwxv2lWbSieZ
VgE6uilbvjuQUJiDLLFiseYs13trJkcoy0F9hDbsuUCJmTD9QQ+7TDUJmEqYpMGydfaw2IVHdizQ
gIZD0tqH5EbHVHTuIDaa+lXvQWBsVyLS7JvgX/uTxrOImW8XzgCYdSUjxpFlWvX9PbY5SKvjfwK5
k7dID5Wc18zX21DIx+Ww2jP9xjWZJ6MmeG3JWymn7eJ3qbMS308aC2bCfpvIEV9wdh5uBZl56FNO
GEbEQdOKHNWBLzcCsDXJwdPosqh/15t0iXZ3rLeNeKfxwPVJGc28pht2IgXctG6HftUA1Tlw5Uxw
qy8kto6TU/bmel84MBm1vF0r4eZnyekEr1NOLf8+Ipp+LPZCDhHP3o1GP5uL5oy+DUBut5mtSlxl
kd6sxRd7nK27v3HuBSK3oP7Wr4giWsEHHEW0pzx5BlmHUsS6h/2QQY45tNYmBm262wqR6X22S0a8
SYi1a3I5f6dTtUJSPBzK0/PlVFATwLCi63pATan9eQJj3FmGhcLm0WAN61I0PaV3RD1dvJ2BspLN
ibAuOk8CVhEBKG0AqpinP+J+YZfCr0pPVvMo9Etzdv9/nYFhwzQITAmOR9WPJJFTtPv5Rffu7geh
lc/R0PAsHKK48kD68tUjrUXLDe+fTDdvxKZN6MRPFKaTOeP5sJcHjeSgr8DK9pf+AVr5YHpIefC4
IvwT9Vv4VQqjL7DGtA/4XmfCy+wrp6JLH1ih3XlEI9v1WxT53jf+7YOcoy3Z6KVSNDEGLdKG7qez
Nx0iyVG4Qe8gszhZk3mUELwwlOoVK4nWSn3jN+y2lD8LtxdmVYDYxseVUFm15OpXwCELzR4nmAUH
IQMhNYnf8AWoaK6Q0D3V5w5ehC7GMiKyQ4A/7tn+YWfN+nwuaYb9Vqbsb7DQinXrIxtbMpiQjLi2
B8S3VZw03ZtVXD/2h37VqCt5QXhG0PPysG5G/f9wscUBPMrpki6MMGvmP55VyCH8fhSkZxRiUNrC
/2LhrmwQAYYqXETse/Ud4a1aoBtNmFf6+a4ppVWSoesrA1TFc8bR8BiTpADwjnhK9QWmS/169S02
kz7KSOSmV9Csj0u1qsug9nCgFa/BZFhIytAeKP1KFVbmn1SUfFDJkuX5la4szBQAJj7BSV2C48kt
rgBmzcAF3w+/f5gy3qPRhpF8hwUkK/mZ7TSJSFyT65i/1nzTJ/8vBqowo4FAzJlvrHBgJXKZV4ff
G05TDMa/nwJ1FEO6npD8mHuNq9Cbm8S/tzyVqAK/bSL5rKWpAA401423ytqQFqcM9YOUHyxXfkSK
1YzsoE/JsqtJNeL202sxqR5OJ/jV2YCsOEoFZHRHEkeMe7U70ZX+AEJ+KeFBJRT4Quqec/hI2uGX
b2O/HIK5M1Bzr2i6hNq8lpZqJytPooSj/7YohFaBrz2erQzrNOSTNk8FhVbwQ2LmcOcW7kAM7YQF
MzDewOdZ06ndbqqXOpTLN/geVWPeKLiwQOF6yAzvOaN7paXugoHjaKtqIdyW8BgRXM6Q88TFSkcv
4689twGVd9dJ3PWUMnBatAqOujA5KKOr0umYncE4XoPSFwhr3KScjdvLqq9PgFeZP94niwtUJMns
qhOCjjOLHghC5eqOMzxHY26UorpXJ3+H/0q46dzmA4U7fGSMcPGhLWuzOZGN6iM/ftY14v++MjHl
uJOVOtNojt+bTaenu7hx3dgT7m5NlufBVrbDWdy3gCmYU78/JgyklyTWa+8CH4okEVJlFIO9lDV/
YvwAr+5uck0CfZcooZkW/cH7NIJ4aRCVjV3bH7kZzwU6HTthZnZ3elTh7AwHD47cOeU2rR0I/ThM
53YqVtP85ttqYttvyn8KZhWyy9fGZa/hgtEeOarbIAUvIx4WGqJhmROPjfmlqFjxjb30jeL9asG1
w0+CqP83KJPBCuW4rSR9wSBZsvDn1++lUO+QjDdBQGvCRTvdq1PvqPC3y6uB0m2gSda/Z5bzRbpG
8vsduK5E0M3ZXfF4k8CR4Mb2SXg1NaGY8L3eD1CZYxwc+PGY8cRro8ARjwn2O+vbty38tX9nWXlb
lsxG4lVoMPUze4aiZjHyw76RszP/IqUwULHhhDoCPOzSSlBnK7QGumnQej6EerKTlmWuyXjTiP26
RtX/o6jzSgakYuew1ovk791hX87NMh+yFK9gPAbkTW4gfWcPJgbumA3xFq6f97HxMOIKxzUil3yY
igsm6UXYZtl7M1SkRzRs5d2JSpl6bpbuQjRHMbdoLHWQpE8HV+xspmBD10c7Zhm/5oGQJ+39dNRw
WsXpNtK3L/hluydWMsolDRPdX6uc8FXtVUU6NqwPErW0tTSP/VDStAVlN6d2D4BVBjrkTMrFezlG
eoVV2geGIopHaZmVXQi5SVF2OjQnl63n6o2TcYusxnaSkmCfO14QW8mjbOBE7cTFWkEEmjhA890J
FYIBLGVn4v3z/iMDeABmm153T6ZSKbni2LVhDkgi2B75vGumlF/DGoTlpCo3Xt2KfG+zL/xpaxUm
4SXVXwgsCMkIVqUxafTKyUzy2cfjbTMRzyflnKoG03V6sGCQzEXbawfQ6UAg0teUaJwBdHTW151l
IdGxDFAAbLtqRKkgUIC3ezZF6M/sGUViRD9Z35OqkrTYqWyfPFxGkkuklrw4hcC2/qW005CqVJGH
uCrT44AYVIVRigJfqU9wbm6snw5J661xycgqGNSJM+dQusnQiZ8dnF/vkAw6gSREzpA5RYhfzipv
USkIdxGsknvXRtGzfUPvqsKOHjGahK/Y0q+wL336KJhTZVX503mMRNkGIEigiB+VvwxII6ABVHEs
v4l2SDHAJyQ+xLpI3beahhZ4V0ELqDC5gvBjPOuZkXMP78HAoT8hlGpNA/Su5DR7/rK02vyVf5z6
z/gOE04GeQc6UI6vD4PPNofjPR3QFsq0wMSKJqJK9OXm+YQ43eLf3wG9EGud0iyoDD+i4r4Sok3D
XRVul+cE6bAVvgL59f1NNSp5kPZEtuoi53uFJqWmx7o34d82pxHF+qmPxrZaI0e5AaRRoEVp1XoG
8dGii1G+Oc+Xji8QdD75ud4y0pRnQ7h/EUlNtGCuzKTy6pMfwZAPavVCltJvM9EaeXCr6X/sX5TZ
QIRAuhk1f0QH7cCvx4UrEmPsYKhIYiFfDkrVE2AhJPVyJpKCketDiUkgFlG48KMDoinJ9JU8q1gX
JzAqRPsIgYo60NN3fh6ZGkfZvrBNzb1pcn0vsuDIr7NLQHLa+EJLD6Ps5QlYd00VctwBEhL+ekVQ
6zXJPojyCGlcQ0GFAKerENbRtEjwunL1i/btqmMzkyPMaQvcIpm5/KeCwj8Q/NfMyDmuQAsbtggO
5aZbgy/Za/qvYNGdjhhkimHY9GD6TcapwDn4AlbmJQ0je1ClwditFyl7uZXoDpSbuDozQTEmFJLm
4dUmn3RBvIUl8YfUC3aEAQDZYpB3ztiIDropM5F984azM4iXZXexLtVy/fij2KNcyya+7eBh2zb9
0/tQqMqEq2FHMaRB7H+iAtt3/1LTccv8z30dilPNvN9s00d37L0Jrh0h6msPwB2wTq0ZtXuvpwPO
OhphEKeD/8x949CFQQC9ZDuxVFL8TQPB56SYV2IXtXgT+K2mjNSijHThVFM1KwSc+NcXRqLfPOCh
hstkvwm6HqchM5XsWtuI7M6acCuH2jI80EjmGfD4g96qKcmt9RvI/7yT/AtPSs5eb89xSD3/jMSC
194i+aCu6dU7oEqlks8NYlDbToRGMy7AiyJQp1XQab+QZeYCfE9IS2eJQEa31Xf4YCxVGK5RJpod
pC1k8R+pC3lChE2l7CQhpR5w514i2RV5p1BhkZnFGOZRNbC0j2gjHVi3sK5hbkCnEDX1lvEUPwLC
0mhGK4UMPQKx36gShjF8Jl4Pvg21cr+xSt33jiRVSPOniCO9Vkhch6XnasfuSVBSq/Ck9I1SH6DC
ievazkJukNSC/IOgfddxMn0XaOKRDE3dC5HZjmbsn3CfcZKSa/rCV3ThiCnc/q1Zelzu6KnMUuh8
8FIw3kEapksAVFpupX44Z3ZxWJbnqjf7h4L0WeGfmlpKXj1BWwb0Wf3xQlVcTxWJnnRaONmgmFyq
8S3blIBU2LgWFbP8TLS9QnX1PqYdhnSn7WO3uARLqkCo1CaaX5MVEm61m0G1OF3mS2gSNK8+nRyb
fZn5fbe06z7X2U9v54Wdl5F2PjgTQQqa1iOYv+3M8pbrR/fXD7ZP8km/W0zJfnn8Ugg/j9VGF1Mt
qhqCMKaP+rfSRLtpzwCc+dM9JEez2YmPkVJHtPH6bM3SvGWEcKOMPNaAkJgFtKwoyutlGMPVQQ0g
2nYc9hDyJvw4QNG50RV9qUtNmCnhyag6rfdYDGrJy0Ew/Z9zWeayn++MtaWB2GzwCd889oqQIrih
rtyeXStTkgb3I8PryMHnrRIHcAq8Nx4ddG90uqc8qo+aP9+rAdMZdRpsX2l5vTx66UNxxgcFrLSd
DavsKbdrzMUu+fKuIkB6wqx8iOEULyOYyyoNJiN+HvahH9lcpT19joOLtPSR1fzcGXRvVOSQ3knz
xEwespD6moaZxMBO2Tt4NQupllW24LVOTWNAC4/wC5vl0LvHNkes41NhQNJUNnXeh7rUOYWyaIR+
U0U7S1wn2nj/w41J41TNl3FsHQEz0Gbs0KFZ7Jw+6LcqXddbn146Wm+vuEd3MPjDo7xqc5D/64kk
6I9xTO0Gi/y/4Zf6NJeL7GdeDSlCcQslzQnkWHRTFwQ2xj23ZXIwfW+NQcff43Twu+HLRVlWxPz6
8xaDppnpAExi0upVGwlssesxOKKmmO8dz7bZ5AZyWycL8xKTf5yUq8o7y7xJ8SD4eSPVCXCqvlNX
y2Y1MD6b2GRfzTlUicfkZ1LhkB7gTZ30xIi2UDUB6GyY42qk1ZB6SuYOVt5CiBepA5tAPtqPT8cQ
LFLqyTjTNIHlwYgnrDlkwopQhjz5ZnKZAH9lV5rDeEenhUo4PYMi3ccxNHLqZ+qePwSX7qobyBTF
suEwFY9QAeQg2cnP27GQl690bVF6bGoXwvtXiFi99Os9ySFA01JOwHM5+c+IyRk/W2bIZCUdAwY+
k2sFY1dbzmtRlIV7zGi62zI36jQaYloI0cRxUIKAEJquopQ+ngWcrYyXKvjI8SUU98t41zi+LfT8
tdBY+XH3UlSZhZf7FXJsqbGIq4pAoFyFWyRfTHY62v63+/bErLx9Od3e6K1GcIRVLUUCxOyXaBjN
THri4llkdkLk+AAh2J79L1K5aZw6fQNzcoQVg5kfRV/fSnjHIZTDVCS1dA5Ehm+FdmpTuibc2/i7
Iu7qJgGtGhZCJfssDSIOD90jPxC8rqbUi4NOvgc+Izu8omHHi0Q4yZ2T2kh55JxPA3UhDmzEnpfr
qVuqFxlUUV/SRbL3iJ4ih87JIR1cpCCIEZemV6KJSNXjIqqqmZNhBdO4kFfx2vkBlPBVDW6UptQx
NowDUVPQbSbI2+JNI+17MxlLiwX6prPji25HI4A2AS3UBIWHCDWollQoeYgRnsBJwWNccGDUGSvN
SfkWDLWk2RvC/B5zfmc/7PTgGggLxLeV8f7O0iMC8TTBpLtxImcMVtI39nMhRYAQTcdKcHifyKlz
Af1XUdVmHL9CVazvjZbdFgzObumGCO7TepaCgD7Bg+NjZIgVe+UjZXKoH8Kh0Yu88IuyIdZ7E+H3
bF7SNpqsbakhrN749bHjLo3ZzATD0ElbvyoPAQLUS+X8rgWoAyYUVVHWTlezMCQWIwKX9uFgr5oz
+O/kIPNBiR7rLcKSHYXjX9RXnJN65wBxyauKgafnv4NHbiTc5xHveEb0HD3ds+/co+jSpd0IU+gH
laI0QSCPAfZ4eCWjFqvA5yC2vP31B+mwmrsQuKrLqF+ZDomoirUl9S67fRXO677j9IWhYPBY41zX
N22w9cZUMPgGJBjwFhQekxlUtxFCkPtnVe7C0s+ei+4lZq1DYg9av1QgFMHYGK44Kp6xGTnFLhQg
HFJiLbTGYLxox+tURQT3KFNjk3vned5lTuTXjQ7PLscjZHS1IBM2xGVlcSMQR7PKn6ezc9gQ3rWf
JK7TI8o2nsM70Ftm9ctGlExPbjF0C/yEM2dGveOESkHe0ItQsOiwHPJXcHkk6zGCoBo70i8Yr4Ab
DkyiYexysodjoN+JWqIJKoHRE8QVvOMEix7nw/kA2rdPhXOYYKF7QAcODBhYSTil9JI5fgsjqHc3
uqUKpn2jYa4ftZrmcYRjryn2dY09/BquCHBCxfnQzbEi38lQWZI01NpDl47/4w4+mXfNtBms7HM8
se842AcYtl5WUvvdsVsbkmgpzCqP9UswmDtuMw4tALOfasxlBZRUWue8vjPebYR9WHT/jAP5+EvO
6wCfRMx4U4AofZuUAzrJd6STQ01bXq3Imosp5tsWoha4Y1Cxzmyxr1ziJslsyBZVtJNUXwiOVShu
Y+GaX3+lCwAxFkDVlh+9us4c/LsiA0P6lTn/bS6I+lC3d/6gdWvHjCeRvrU9wvtUVEHocClM9mBQ
/oro0cwPGrw8GGjk9W81T4KpVGMh3lLd7nz3jOWQXo7a0sw9xBZQXL8lc8zsIcYszBW8kulja26O
3SHmomYxGZcSJ/Ph8riUrZZvqlb4AEDLXyjeh8ZWj2r2GkgK0R5y8iB0ksSTguIGIxr9/hoAFKIp
cPZNBc6dAjxRjncY9DeZz31/iMqBQ1ltQfXuqfUs70agLUxgO9bAnz+IHyEevaMaf2dE7mdJJ8tD
lECAntf6+HdSgIPWpoq6ai5Q7U7nOPb2ql8c4/et1nCVKp3tTDvLIcK4BhfN3q0bO5YeVzH7E2nx
qIcoq1a4JdyhBtHJL7/CxjcmvN4Ml5Gi4y+Ip1zf7tAvrwwEZ7gmG6Rn/FWxqTO8wjTphxUtCj3B
jVb9RO7UoWymSuraI4ChUU2L2brEzjW8xcL0J3oRBw+4j3j5wpejLM0ZWw5k0JrTeJfoNIASH9K5
tA+n4cK1kFfF9s9iiDryovUl3t144/+ir6ggT6lpzTi/jq4z8qaBBw0PV6oc4V7igqnOFn1nHzw0
yr/NMdcC3wx1rA/swwPWxPzrbOUCDCUyHuyiTp/H9saOa3xj6XBjOX33YG7vWQuw0J6/DqZMeDyQ
/pWUaXlG+XkWNcL6VYWYQNKCt9/KjvOT08QxodxcukyFx5vLtbYjMjxIWdcECiylYabGYuI/L108
mmB10ecAS0o3KGM0VwPitcdOJFausi3iYMt3NxpTqdJR0F6T1P93CkBnFNpu0jvwlKBuPdZ+Bjzc
C3p2rafnp2jjaDIIajxLbSv8UjxDY77ZqS/tezmYHncjGrJXhiIocVLw2HqxqbMOA414Z6XCQHGj
zrCdPBBBUmia/gu30VZY6j5I0+4IH262nIAo19gyqHzMvd36A1op5zUKzMupKaMrHY9Ukahc9unl
3nvDuz90RFvW+Ibohoh+0ra5mG5w/IyW5Yutr4rPdDiHE611paQGVH5xrNjBjQgBb2ZQTNEtZ4eo
TdJT66RtnRVMQ1jzkFpGYOYhD6T1sR/D8TVJDhp9nbrwRUaYKS0FKV3xj+pszPT/eJ9EU5Q2I5Z6
yL9HUMV7ZJ97pTfJEFtdCuJslcRIqq2vqkBVWuVC86rcK6NdTxlEIVWISf0Dfhg49K93+37JM6Ar
Dp6zmEHan5Pz04LEr/EOik+DchatWhoAP4ukuzsSK33LYzTOFIyuaKsHQCyOaKnUVgSkF/rxhCk1
DPnJAYWmlhRfIenNNpDYzyTVporhjNnTGCUe4xyY3gUkHQ7I9AQUMnUNEx2tF7+DV8GSn4eN8zTC
ltlcAjjCWkomkUaW+J1Aw1FecqqnJKN33gUfQ4fYqtmWKxHZVUYVtU0ixt/6xkaalClT/bOCxvtz
uwaaB196VchNDEgSEk256boOwsWiH6ycRP+oGSe74QobpZNu5uOM3ACu5SiBZOO27uRfTnaeXSKl
zeqetfq95uAUf97hwnahoMIEe7JbXHHcM38KMHJtqeU62x7czj7/7iNEu7jSqCzW0bx/viocgIw7
C61va+2sfUkFH/L4FJjG8jS2ld9bsVrF61zXlLJwGWsrVIskWGqLomWo/V9VQT3z/yhor8jdXmgK
mmDgxg7dt9CwR9ujWIFeygZUuc9TsJrNZxpFpG5PKR0KXnxBBwrIkkca2z5CpMSU++vTMhnF4+e6
MYlzridMj1IzYWALj9PuScgd9ppfLgiIWLxb9qtJKD4Ng7p7BjJSfs9m0aWe2LGqufP/C66jp6vu
Evs96Egt0iLDx17biB1djt7edS5zyJEVMHUIopDZPPDGSOLCBPkm2z8TDqRyQnzHd+7AvtcAhsO9
NImAvbaDWa1ATdTU9D/p4Nc/64zRi3i91tcTkAE89e9kMTVtXttiobTs5Ev8YMq490JZzIMLYtrI
dBWOsigKGuke6HiI84c1fVgJgBrujj8EqP+OvFrIYaia74eEVu42b6qVGLFLBlDj2kqxL6+mJrHF
okmMfCfTdfnhmxiD/TeNY7RjuGHC60+vw6CobQFCecCQ/Ka/E8frnxIyiTozi7nfCfotuyCgktAP
J2HdilkBHeVARUMQ06wJ5Gccq/ef4GfOSO5fJGEkKbbi6GOKtnqiON4Ah3nILnZP1qMylqoYI2HI
BDR/5Gkco5nIIY/iY/N8y/fG2agUHadXtZUeLSavmoHba72zIc8iE8tqrO6LDbvF3J4+j2nOjnGd
O0qBu7BwZ7Ha1cocqoQHmKcxnlrrBbqoTCZEzJWhiOaS1IuUoBrvZ/LsQOaulGcxFBgogg7Viy4D
l5zVCkzKLe78Vp8qodni9O0acoYfRnM23vdjCHGkG1LQ2/7DvEY1aruek3idazZ1h1bPeTti4KKp
7W6dXrZBm+uJjH4MDCWgPARtkAElArDcfsKVr0AfJstuuZ5O+YVWkbY6H/H09pF3r8+zCz3Gq7b1
QtWDWr8jnqfN206U0wj384arF9i2xk+G9DWM+K1zikJrDegc9dtqTc1eFufJzh+cD8j3NgD/Gn+a
IygGCKmaTQn4xTkUmlBUc8yuzHqIRzj8riF1UHPcfj2D3nZ/obxbgdXaPRahv0A8ZnPQMfzH9c7A
B3J+2FUoMi8X8kwd3hipJVub0Z6ELmySl6L4Ande//Z6gSdv94fEfmtkx6aRCHCc2O54UWhtcCIX
SX7PSeeZ505HFj+T48IVuDlH2lOCOZhDuiqcj7PRsAZczRqRja5IOClPN9gXbc6/IPWviSd6stbZ
NINAD64LH6ANfcH3JFJgq+cYmH1Xw+bI8tZE7obOO8dhk69X0n4x4xULY214RUgvLpZmn+dAEL/o
qpQ4dZc/0qnpUgNxyrGMke+kLkkfpyQ6rjvOq9xnDxz9pH3zufeRPZUc9iTNwjOZWmk56XUJv2g8
gf7TcWdM+MFeOUk5/j0C1mHQ2Uh8nhaNpJrTj8fwhBTcglFZ+QG9MLmF8Lp3Nu65s8A95p2tXKL5
nUawBQKoxqeOJfs4rXL0DXdLA/MY57QtdGzuk03N6udwTSSO+UCIfpKSa0Vzizf1Oi7DBEpEV2Vb
1CDBbEmCd38t5DsrfOHhq2Tk3MDDWbtEPtUn97IB9WvCD5hl5HCyFk6H6XdfWqdBbQimitr7Kdl1
NJ9nn/1inwsHERwHUvHrLS23LMzoCcb80BoWeSujyRgGLxeu/Q57/NtHYH+A8Hl7fotUiWk1fmj/
9eHOGx8nJb7US8Cm5hDaBtA9gJILF935NI4k0nF7beYgeyxQKzTj0hIc7bWfh5CAZqY2kbeWXW8f
PHHAB6ZaaSfjo1kns2dNIwQYj+MF15mh2wPXHz6lBbaSCg1u+gXYcmXKKlTDHnMNh3Q37mJkWlth
nlP05OSh2MgSQxoYhWPj5JIEVFl3wmHVCtvaupE0tzlAUkTXZuyy/rsf8jKiW28PJCTW8XsB/i+a
1Ewa25nojxxKknJFLiySz0N2wDHIOsVwWUncorof1EniYcv079jldHs+sLamblJRI1/DB5YEx/yd
gWjblTOFoOSNDME1xFPYCAeK1963Oq10TLm3LuXcqeQDb+47Zr/e3DRBuTUdRvg9XT/vT3TB+qlu
hnx3uOV65lN4E2a5+QQ5PeUvM8FnTaAOzjSzgl9fuUMs6o8zHRVKE88wo7RKzaK2sae5Ivl4r5Ts
J/k3i/ZczG8ijqrxY2ti4IC3qcdYDw56e6DH31XIqxi7/tGLdVVHGAy0vl2cVXnrV/AIKtir+YHp
fj42UPAnPOapPrnGTmzELY1f4sWiI6XxTGl/lpJjRA0d9tXpQsucJ5lf9TWK1A7iYsK3Yasz+pKM
etUE5sBh0WKF6AK8+U0pHfbZB9CbDM8eX9P7HZ8JsNOUO/EjkBADc694qiMUa7fZU3GwDo6ht8bm
FQU1AuN/9aRhF/cp7ZFs3Fb2Yf8mw/vS6379v5SE1sCvXMYkagVGZMRSQtvk5+Y+SKcmZx2hloEb
EecavWQyJ4IGU4jEynvb9s8A4eFentSDVb6cqBA3rf/g5VkwVItH4tjJbqDvxgXLOpbaqZcFSXzQ
NmzMcLcT1ghaDYnQhkQUKwMULf1bGg3KCNS09VweX6g72BY6CUVjVcJBKsdRtWcBKJUnbGnuOVeD
Ei5g+6ANAyZUXeoTydqCziZ7v8GLCBbuW0BBk5D7/ysKvPk2o9egr0ET/wl5TLwD+sEHErwwjOJw
T2sSwU7631+XjIKYa9koco50wResvUCsvWiSeSu6wv5tplblQfa1wBvOOK+74uo/76I6k3tVWLZa
8E6bex6PfVosHBEpbgSpao1gs0TOeIOPPrGY3ufMlPwFlNzUMaligd7OF23ky82WID2x/T0zRBcX
JN+Qk9KZFPkVS0balZEHmZaz0BEKTAjsbltZaWW4QXH5C+9w/Y+tcPdymArzQX17GixPq+UIbg57
FENG43aQ/Bc7+f3GpUwMuDHdn3JqQkaQlJy8ypa7/53A0OT4Qar1BZNGma2tijRYtG2Y65bMP3z1
dckK6thhxNMExh6NqI/5sNuuOCvoJYfqo+T+v9lKhLQbn7hBVJGsbzzdjj+oBVRxp6JBQ+rZVtJv
66pHAmlmeb9wZVfUNu3fXZeAa0NgKqFkMK9g5pG5LVeUe9K2MVpr0CjE5+HaKDdlbORKjjVSb0ML
nxsjfJ9Fm+yeJev0NqIU+AN12HguNkLHhgHv+kBtSNB9Uq9xCB1MaPkpn1WAgL8gSFDxiydB26HZ
CG09TZLmergTlcSa72lk4S4RcjaJVRr92Ebma9+EiJ7tuMEvPASJs7o+JF/2Pvnjjr1Cs2Z3v07I
x1GXoPfD59sPkMlPWqq+XCzIFS8W8XP7T8JGaQj9guKRD1WQ1m6c7V0cv2LIS43v+7NkZU9PmbX/
rd4h3qN1q3pbEe3yJycB+4ZB+E2vWuSCo8eocQxKH9OY7xT7ZBIQPIyW/UD7Rpr6LyICeDwBeGwC
aFsdGH7w11gBufsTwLNEmE2XnNzO0VlFO/u2zV61deRZSF2P2Vo2AagrviLdltTtUIRkX72X5+Be
I5Hob6NA0n6o9MMs3Y0tyULSH3dfVvs0Ck8mxxTOpIMnYQpiGYwfU4O3i57ppYDF71mBcYO12+Xy
vzXYlCpJ5PgcvGqKdEegkaqux5Rwewz8D9jl1kNMXhajulZGp78HasLBssoC2TE3jjjermqmXBB1
x6r8/ha/UBVNef1sLF73Dd6/IewUFVJY/9E8ADoxEnGLNywBcfT3dP9IxEVa4SRI443JX94xpxNS
OeCbXGBJm7lZj9CsohFkKReoZEQpN6or3SOYWolYwTOdQfkHEnUKMxUPfSNkZ0LuqW6rE4vC5vkn
P0gFFH7Id+1UrllNt16/UWA8Sf11SLweTrwDRJx3tK5aHvilK1BtBoYxonW9lE3dF5FO4L5YwYiv
+nPil9DcfPU7IBPHJyF6VD8Ep9VbGAr3pwPSwEG1iQpC40UNs/lDXomR8Yp52tkNJi+SP0RWNjv6
lkZ+0On884sr3H630iFboIm3ekvYrewe3LqwIVkCqaVR9cbuva/mD0/0HhSHaR5aSzIpuBDWyRWr
wadFBr47XRS8RKVVr+hN/OHBIGrcZaWlhtaTchr21seaEv3LffLdXlYlWlryXu1a9ZsM6Ek3kZQG
D8VpH9+7pD9eSfB8nS/RXjpxRQRDK8+Q2IoWSaQNafqzS/xsF1JJUW9wefSgkJoq0Uthw4pxXWyq
+hWqdVGH1fGfY6bfw3ZjAdh1nAQMbo7WWkYPsaMs71hEuWTmdje1OEijhkT2uOC93A6xpHV8QMMh
cvZwlnB7vAW1AMPNFpII/PHVGt1jri9JdiUOsAJJccZHamAeu1zhs7IzupeOcbcXV/bOU4OxQ3zM
3gNGRTZaUHWT4Q7KT7CCgNzJeDYN05xPL/N2s857uy3eCoyLIYeX4YPKLyr5/IFguY+8HUeXyG4x
FDKXAVD1UFj76EG0Rmppe71w392Z2MlmjRI99IR1e1QscBmnelDIPLfMGbT9xs2MGPM3BsAEWpfS
vxBwqdG78/ALMgLwXSpiKNw2zEYh+4IhGoSvJFmhY6pP8z3SunENUs0Obkeb0xWN6gGzMdTRqfrg
kDSNCx6AC7QAdgm0mYMXssJFNRQ14j07LMF2BDeYNoYgNScfpHxmLrc2PHjTOmxchcS3iltD11Vd
vTlxp/i68hQfRYhkftIWUrIHs7qy4CJxFzxEXom9ifg2/DsKG0ZPrz7iSEWY2ljAapoO4yMD+T4V
QXHjmFfOwArCwWd0RlNaTD1cVs3q4gR4xGBnf6T02pxKHLKB24jABoOHul6V01V2bz2PYqhbU6fG
9lsMFVF9Gk3LBVzKQ0MQ+p/pHh/DeS7KCMJU1TXR1VLya6dqgniZZzLqFDlkxmX8hvQi9IBoynWs
tCqWtOrsQmf+iGlWF2/5BCwNlV5MXBb66eG1h+9k6Fx03LL8Zmv80eeJbBw4FQq0fI93bgaEji17
+NkUKZsUvT2HMvECvPwrqE7RoA65Y0KDM86RoHTi0jwyVLBbrWzQ7BsoG+yJNBdvzGGTJcGCaIXD
Fp8igsiakEVeRVGRkGgOMYkOe0NtkE06s2nW0Ocf5aEYZwzPM7jgR0AWwdgLSJPgZHLqALsZUYl2
E4LcuNTdCOOp5gRUTQLMooruHSJfAKvUL/yTIp5vCyx+Gm1uIwHDPVw1U4kcoQo6z4cRzdIiZuz6
QFMy+22XhSZ6/jUApjJ7F1uy9SkizEgjSuCqR6wTzf5Atb74YK3YymOfLoTqLFWcuBIZaz2QwrKT
D84iLKacYT/EN2AmIF6FQA06sNQoElGZwdelVK9GNJZpX4kGTc4Yy29r0C12lfIPioqbhYTnyE9T
EsAOzcYPzJoMP9htH+GsWQNLwtDBZDtOaib3jBdjc5ANGLxK7/zUgd/tOBrJNtiNUklAEPa+zWzz
DCZlSdFFhJ01ziJkQBmvfSvV54OhK3U8KeVUPmww3m3J2azdaQh8XMpPmGCglFgI1X3EYnrFK5q4
Tb5/00sJwOs2e8WYDlTh+x1QXqFSIF2ajO8gtLs6x+XN/ND2vXxd5ppu923LtnT+mYgYIuj1YFNg
uBjWHVINPrFz8+zNvO5PoCf9FNSohm8hDy7lp/uYCgZ3jpEc+ckjsHyvHlRJIpwe7pvQFK8MkpOD
zW8awvqW3Tnjzk1UJJibNNqLFn2JxKC6k5DWIgV4nYLAlvtQ2NdgwjRw+096NZTtUfyy99WnM6Zx
n4WxV3EtrTvYPY6MZCN3Q9ABz1GkxEa+wi9npwOF3aufKMa0xHWknpWWMmqSjbs7wWsFydb9AjvW
ikmNmOqRLN92lyULkVEtIiyfLg9jg2Mpl8JxJA/koycvkbI+MITh90g6+ljkbo/yC8zbE/vSrZxx
j+a3jFk8IfipDIg8TEcRCMJjFP0Gy8QPw13XGgLyoDgVK+Q4A0zbxkxogcN6/IRjXBfEpkPr9Z4h
r/TzM6uYM1XGl2o3QX/Ms3hWsMLDSBSyj0v8QongU65zf/A1QfBHqAGvYA4B3BaMLC+sT2vxPT9c
fZcALJCTISuHD8zUufQRW40Vdz9Vw4YYONJvtXTw5RTLuSobfkbnvYfmGERrM7lVn3RAS6fAP8yw
bTr+NgCZtL9uYgFaR/oT67M8lc0IdIPi7kfEXjgTNgNjN+gWGRSeVuel4fu4Oa94ehfnFZexKaa3
VPYVHz4pMBLvFeb7aavZAcVEiJvElCo053/njw/wSTcCSzARA52O+AHh71onqsXRzNMm/gf64ReH
h74/HuJOZlFOhvgRGSq+ESKk+e7fdPsP+OuWoERyfRa0QMM6UW/H1Z6nGFt5tnn0M4+1ZYF/z7Qx
bdCEJaVlQ7waRwlx69dh2glPGCo4dQpLouXB6h+TdLt/VaHxxNu7jaPrIsaukcDCRaA6RfCNwhXI
qgd3L7dfrOeI5JCCKomD9nA52Kl5Qd63QVGCLVkA8LiXBdJzTDcbGcc1g8vjdeMUeDoko6ejMhfS
Yyho+1k6EyfCIL+W72z2It/FwQmGBdGTAFqQQlVR/6oLa16A7DF7wWylsRRQlmft8c3bonJz/Gg5
u/2XtSNcFnkacIN21/ynCHxwfe7yb9PLKRk17FM/WkLJJ/mjm+0nrpiZZWTzhiCGnGlns43PnPxv
vqht0g4eSutgWBpqe+7kvvqcckFeJezk+3JLDVmh42zU0W13DnhN4tftj0SY6sGNuum6/vLhcApe
bkZczMxVzDODx4zatvzRBJ71AHAnjHGWPxiAfaL4WXDq0sqS2ygEMeFYpQTQKL/BXdAgSl3gHOKc
LDLspbGPBzBYagsuUp3LFdm78VhI4JEUGBEzAE4agD6dlVP6NI7b9ZRnWjr2X2zUqWn99TuBqv4w
siTmc2kJaXoUuemWXAilFgw2Pr9fTooox+k93OzL8q+pZa1j7fiFe2DdwhCFt+ZPSKF0zos0ASNv
+G0mS9vEpSFcSjb36qsZY4z54+zAyG/k+efBAHrLNv3gB5ecmGHSijx7vG5S3jtF3vOb+RsUKFh3
TKYQcJ8cRwhsBUx+ek3g5jEMEVjR7nVUO/ypi3DXsxLpckPhru9WTerdPdjyMWyKDDekIPSgkFrn
1LYA+JDCDZfkVHc/yWNQRFO1g5AWV2KG3FIxGp379fNTxXDxTrrg3GSgoYfXI3cxL+39bf/VSi+Z
BQbFt65jjw7wS7TCniZDzVT4DqOLePuseR4YcumdfDxCy2Bj4Shp3bqExd0SMObPRA4bfUDM0zxj
dOabzSIbGm0TJ1Shp6fHJG12oHhKjIll3t01gvakFJgSVzPzGd/+qCM+3L+rnXKtORWHP25bWxRL
FpkbnQop4QAYJoDR0fHicOuBgqFrNEIAdd+YimmNURZuv6Ahb+EkAmbbHzP21phtlp00Kc+mIg/z
36esLlXd5AHDF7lBaRu3+RWTcDyPf9wSQcAdZulxH2zhkTjDkR3BV71yKIkJd5jqBizR3z5AaVfU
d+JUKYh8ll5DJ5rI3LCuSDxr6OtTcrCUkXWFZM/5DlvZZbJ6wRAJGdiqMzpzIwNQQpYGUEneD99O
ghOK4RpjpUWMr7SUmv3jv0Xeu9/wKZ3/YxHCpmjseZu7O2ZpkJPPMtCqygsWgj6o1LTD+t/95p/u
LOGq+fFf9sMYnwOn4mArrCdYIDgUkjckxgr8ZbMXntHxDS1r2ghXs+rjx0F7/II/+peQX8XOlMM2
mRBQtgLD5Tqyl0ssZ3Z76U1cGcttr7M4x+URqaU4bydgH44DBzPk5aSlXo9CsLaUCClz/cZ3BOx4
Hr2HzmngarGhinrDFkB+3znGFxXZiG69I7URkieXQebzIMeqdJedY0ZWObV2BSNaJWa0oR1YowC9
1DLr3bwBG9XdMT1iIUZerW+anEc0ERgs4KitOzKNtZ+fVnI1NC/DQSmqomZ1/XVY3Mw/bndzRDiy
xVg2l+upLxLTFj0wy3mPyhtvEjil+gfnPfD1qIY1saXIuyL3nTNgNnugFam+im7ufuRQbbDRkLX4
KDMnnZ7EmAOo3VEijok5omVuh9BoUl5/2xwqwoyP+cJkmSOV7umRL91R0UBmJ45yeFn+Km6otLTo
iN+q4F81yVkEKo7qXGdlbEevpincZ1qF6Qn2F+XMmg/7dzkgIhogZXgpEJNkRqPZQkh/gVfjMOk0
vwacqJHvyi9jc922WoByHzqizuaclkM9cbwb8H/1KgwsuRCWGBGk5m8ISM6SES+HpLyeN9RwBNu/
08thNtV/Rp+HSrXLjYEz0JFxh6MAg4VjVrXZcLk/IvMPV7JgIhJZGbf2zKtAG421hSndRxNE813I
QQ4jq4X4lq1ItoJ0NF6MNGcWGBrFfODLv+/xQTgBkeG9vpnLCPsYj7aBv/j9ZGy6JHZ8fIr63phu
RiDfeBeTN2E31L8Gee1xeVUyQXTjON8KQs/tItnxn22hp1KOM8e6cpCLevAVaUsITLBCB4KfbHQB
KLUlpanpkBGsnhj9fV16oHXrN3wfdlVP2L1xqW7CatGYe9Shmwh+uylgEq1mXqSYr4tWd6uBWXjy
hefViFcpKAFS2Le5MH0pKpRyrLbsRPS20iUTN6X08yG/X5Fr3KlHlWWVB/HtKriOSWCZCc0P3v8K
1o4qCyBhaNb6KzPmnfb0R0Yvz7QfGDq0vzfgd41IwhYXM9me9NpS+/K4cSju8RSb7WcSUMp8//6p
Pn25IheFHOXVxKoH4N4x8BbmFaubhck7knyFAk7Bx8TiLIaGh2nLZVXNq1k/zQq+8Yevo1MdXZp4
q/8O/BWowQM1oGl5TlgMSnsSI877qweFXV1mA3B926VRdXJsbS7t24gGQ0nl9Sb/eXJTA5+xje96
Wqd8Vzlgkx1ExhtZT0S/o8nPK3PnMZkrjeAZLc/wzRzvfV7cKkaB5DogTLgcs1hkZdZJNu6v2JxZ
EPKkb1FrrYYpFHUXdfdqkfzxaKw/5wSzdjYwGKMd6YLsnLTgmE5RBiFqA/Bmro83YQDPGzLf92hQ
ghB69qqx5Iv9UGo9sH7pU1p/FBRkUH3rBpfvy8PcQGoY04MJy1N58h4AMQpXBO2Onj1+xD+dZrhe
dxmEoNSWt91w6YP77u+OsvY4tL/4FGG3z+jW9MCsKtBNIzso/cs4vL3kya3eBCfNIc0m78D4tnZ1
59Ue6ir3xIEmdHOvPRVDtTAmyzk4RLgpvPl3XBUkizfJxUEnAjT4/wrd11UjVrr1W7TUlmGHIFrs
qs8BtQKe9hdgEWDFdXu6TenwX32dL+il4YyJFV/+9PYuPiuTvxfdw3H17hZIBTA3RWxW+N+2bZNO
L60E9V4d6lmhWppUPSSzpcxtUEQVam3yFRCIoUnJwTl8kdwptFbp/2hWd3UnHCxJOOozU/9Xdt5P
WcvAoBixQbc2bqW+sUkQGN1CZDBQml6eS3T9jDJFObLOK4iV1YPO4H/R+0pHeVcNga950704F0wR
5wym4hl33FnVP9aaAUrhfRuf4bngy0C11ZrCd/bFk2IXBstYASYUmkEVSM+tv4dEcWyyDlpR6IoH
j34QeoJokusBQPmJWLc2z/faefeR5GtUTlYfO8mP7qs6795fTpQ1RvVvuIlxjtZgz+VSsNTX3nXm
PuaYSuFeZ48hZkr/87c34HpEnbuteo0311uNdT9uPDlP1XuRwwJrjrsPKQcTt+xKujt58+SRGkkT
drsousI1hVYIx38PrnHkyclbItq0/x7WZL3wK+oWC4uDmRhVZGX5QKTGAfOl1ctmtE7RKZOshl/U
SkOMh4wH8J+9YwaOHSf9Zrd3qik5hUvZBU9tLnR/SVSJyN2zV7MoANyhbfXZgOeLr5MCeQ+jdET3
VuJthG3eh3fftBhk5KtViVjORLfVJqI+P+IP8VX82Mrn/xJAD4h27E4NSnGQoyZ0MJVp28VwooZA
2axek9ceHXswEX5973giRWX5A7bDXN+H+MM/IMc2tdKYBCf7rx/byHcUmKlISRbf5FuMvy4cizBJ
NOYrd7Q1A5oES3D/oivAB0J1Ki2dutGiRt/MaPZIrY2YSwvn49/10hYv1Iod315U+rDKwDKdcA32
vKMriXTYXVh1i+3CFnsUddkDhfQfeuJbkZv/9c6QNnhTIYncOfbL16hilNk11uHV3BFWW4xP3jXT
IX64mpNa6C71Fks53ymt3sDjFMa4ph/jRHsKWIA8yKhsntvJ+3cmVpVHsdvflPlLan4m5X0LDYFg
QEJbpWz5y/C/MDI1shjdOAqcspsGQrfebI+ekAzni6M45MdhvUAoueR1ZjLnXEHLLW9OzjJTlGEw
TPAMMqMGkyxtSiio6TyZPvDGnteGdyNq3DGtcX100LKw+Ayra6yh82+tuY7XGAOeFNVMw01s9tRM
1LhmsmZtUNgtvHdU7qObU+PHICxPKZIbeXW9lUdB6bJViQRoJBIFY27Oo0VG7QuEcmlJ68dTJSmQ
QZVnWdMgo67qac+JiOWAm8L4fbLbW+ZyWn50tcgYegvage3zfkEzt5WZFeIHlmlQqZpkBh5uvlWA
t04NgidYAqUnu+3h6MMS34Qz73arvu9eTe7MqoXZm/73rMzm6IKEnjZdlS9cckTEF9x/uRnLLtB0
ZPenM9AN9/P77bfmkIdqOYm0Fog9bZs3HYAyVrJiPi51KKr6M8kl/W0gmv1RRfrCKo+beqTjio/d
ArG0oabz5xKZPcO93WIRPX9QIFq54FKlswKV0Jdyen/MXgfWDWcLosYeSpYF5V344zSrQGTBcSj6
6xY7bYMmgRI3fSVAzqFrvItjM/VayNMHA1TOm2ORLQZ0gWsnEJzBMkyAxWNapk14UjE7wcVkMaEw
YI4mqJnZ0exh1sBdXsuP5GotxUryDHaU5z6kf158JAFaLDKx75xVDqYYr/QeP270dMoUpvqMVAIK
RmjlrXq8JSqUNtBo3ZS66h+mpv25JXXwoSDmh3W1Ff6x6cT1UNm3SWL1ib8MWZfYempeutowx1r4
r6IN0sItof+9hebiQTHXxM7xaqJmMZFNjsH/TVqCBGZJi67izAFpQwcBx5qBfJCfIlMrPcnZ+m5A
W1hKBKw/NItEMR+yoeu1/RwChRIg6oxnNmA6LhYvP8drL39fit7v+VT/mM54KqzejUYbWCL6/xhb
mjTUpqHe1s+t1drk0BXNhfGOQLi+cTkUtyJgYoW9vqi2V+T5Af5jLLDYvqfLw+WtP70EiV9LVuZc
BmBiq57fU5vreRdGM5/O/FUR33nxzeVn5b/9I49UUVPwaZB7fMbitm8fX29/3crBFdLMde5WoGJ8
Bca2nZrJ7CosyHK305IZBI/d4w4kzSUay8ga4eOiIkP8XPbCcj1+5IUNss9pmnCGU6G14hMzxkQA
+JpdFrM02moClAN6DGWk1ZKPrUbBSdurpWr/9/R2ufCATjYF/86wp2SWPYa95+NMjuREJHkdaFyP
wAsfBNLNgKvJ/QHilfIQyqIuSO+8Flcxbk+lbMuRmw3TeSTmokDpmYOsMvKzjoHH2VjRJArtJNJS
l50Ro4xYNZmMA3LsfrQxFs8xAt5ZGpdGqVr+L2JKmDjIHDLVXDGr504BwQYjAJFESuXOagr0jMgD
nbv9qfom572KRpCoMI7yUXsOr9YqAIV+tUMB6vb09oW2xVrb3/Rs2r8+JRzFd24nK9TudgUD9CH5
eBqem4wgoqBeA+9v1vu0Fe5bW/vTMplZtaBkcpPNKZiJaQ+VE+EEAJMMANNJGtvDtS4Cb3juoRkM
Hca0q3g+6+5PQ9rr0o74u4UrkPIp1t4ET6wCpLOrSSpqQWm9JvfEoAX7oLGbF0JwNDaALBTCNi3T
3eYxU9EoCavy4vq9CCns6wl2g41ureSq67v3wM4kHOv8fmp0fRyfSmJAMlT0SGV2RINh7UhQdTou
idcFMGbcnfPnyFcYvyPQpuBVxqLg7MWq2NxjMYT0QO/wL7deUBWs6mI2XreWQ6nq0kcN04quAJ0m
OdPWe2MST5eQYh/KvSXabpuqnBEX+V0yjRBdWzlp6+yfm8WbjhFne3SX5Xy8TQr7Gwm07mzq63Uq
nBznbnwFi6bSAAo0b+dCuvgNQGVqC1skvRI8X5HyH/iOqRxdJijDngziro1K/HQhctwVqoI1nfkY
vONkvGWEymDtL09Y0wtFPiewUqtsxx24xQSek6rWQOnygkgfS6WLTgCcfiNbRaBJ69uea7KpJfU9
zGA9KYjVhWkQIX7C4cPguEldAGVjc24FoN4shqXeql+PBQdjPxpHhBq33jcZAuX5MctQaJVoOUMp
xJNq5J9eN3hR0VkNxRv9xnTTK+G0JiD2MeA4AcRVqpULLrsw/62PTbhHl72zOaIqGYsNjyRVoKnJ
9LNFUARcQYzo3wt72E83ZUY588Drtgl9aaOAQEhAEWeP9o2RU5/UxXzVixtHUCleFgZfgyzLabYl
jbUvN++wrj1CABSsyDpO5W3W07v1KiGALmmTmr1d9T4AFqDE8qkC/QyQxWMmVfiSkUHA8kziEcZK
uFT8v++DVFqh+A82JSbBzIHd7jkuP6crD1k5GsuePDN5YddZvDFHjyfhkv0CtBmun+8AiBbfvMFz
xRc/qkz/jiMODUp3Ej64nzR6AZS+XqvouuvMKnYbwCUUA0r1EmyFO+zLkdsd7rT/Uh1oJdtkA/QK
Vp23ZwRCADXpOzvYvmk+Vy8UvadWidAoh3Rl0n4fv40bhcOOdzESe5u9/Nxw45uG6IIZm8O0SI26
vRXX5Kij1oJ5T1oaBiEo4oCoMvFD8xFNABGvbWTXIcKS0JgZ+0c+q/exwqXdVgpacIqT6DJ2PXkd
m+R7jlTLXeccCrPrlW5SIVo95g5vN241uB0HfL91YGOEGNEg4gfK9OjW8ERNgMUnFHJtYbrJ08XK
p920yP+kj0cVENoppf2QEC+hn3zIIzApVTEY3huzRTmuGtXA4fL70T5+SlMVAYN9Q3CbTGO1h/Eb
3CSP2Ab3uo7eHnQh6trOzgWRPg4YYwV5/H9u6fyBp0ftoK5CJYODQLXGJhBHEmFNLaK7v3WNeE+a
g8HVo1SYRQjqzTuLh3OyMt9nj9Sm19vNY5jfkzTlYJ1ExHlAaDqTqqOLRcD8z+TzFXuzh5AV+lvs
mtsUJ56rbRUYOje2rqyv/AZbsCadkOnOzm7hfmSN7OsFfDO364MVk7vSR2nJz05Va6l/TWqIJlKN
DhXBVevXxTzk7CXcM5vtSP1CWEa1nxrXznZ2S3S+2uZFS7FqdWGTzNH026gK7xxmzQsV7sIhyVHJ
vCo5xEBErgDQTVIXN/WbRV2mIglPga1y6kF9PFCfyDLEvJPzOAZF6TGIzugSI10sVBg8WxfpGEMB
aq27TJMZaXwPqciBuJePyXo6Ss5Dy8VBYDJZ3XYlHqObPTXWst5T83VL/a3J6Dd8X8HW7tE23+rJ
YEEGZMECNf5EYOM3dTfIViAZ3ykFf4CueP27boF7NghT7H6tZvJYkwdIBFqxxkYZwwzSgYhmtsCf
TUdHgKP9bPkB1hoVOgqC13TtPFNF3K+CIY/6WOE5kvbsveI8h6PYs2itcXHz8Z3VuUZqVVCuBy38
AvqI3USFpPCqJ+HU7zEQM88VM6SK4wnxCaxV+Xsha7ZkYjsETKxS/KjlTHwt4w6psESEOnPdKu8f
MxWgXpJ/I3J/cwXBewgPHpQPA+MSXH4oBfQ0LeD+6H7MSRP4aP4y51kQivzImxddJevovjbBBlX1
fuM1aCQlIUORcaNlijQWPddWAp6Qi4a5HAvXshCPRnUUXPKthwznakI3VfLK2tyYo256e5243snk
uM4jhim1QIZM/E5Q575tLPRH3yab1CdTSaSHgShXwbcBCcNWmJK6+/tl2JqtqZOEudNBvmkqPeDK
oI30Zet7uMQpR/ZVXUWSClN2VX8Qnnz5B3Z85AjyF5aH96+f0yobnA82XE/VO8i0LmcgAQohSEIW
Q0J/naIGjADg/CjHqd2+WNXyKXBr/+C/V2SxZGA1dmbVRzlxxV9KlFzf/u7nkS/OfKF6odH3LMHn
xkewLAYxu4EcK0OonxAx5HMBT867aIE8/LJniRl2uE/TVpXeqS8qC/CDzv7YfVZVKoNNWeVlJZtO
ZULTbuyY3sklhxE8eTKmL+vCsomIl1gomeRUiCCEbUtcDVBUI/OooxjWxeCtLfUQC+KpTz0S0XPC
i2fg799zXCNSRHNdetQs9Pz9dPJtE/XkV/RMnWS12aeZjYzTPK+99z04JJo1tpwWramCStK/CGDV
tEwDl4ec2ArdcLQ0iZ3qJqU2duQ4cbiacLoLlTtS2kIEbbGiIKq7rOLh6CONM7iOXFjBoc8aPhjE
9a+mViuT+NDjf2E9g8mtHwXjHOne8E/aOR+uA5A9KHZRyJ0exC14PxVs/80rzPeVv4CLT9Jy2VMb
HRORdKWL6XbLpdZROVV7cXDv6QrfHC9fdYLiiOxnbzBURLTg3uINQH20nfK+3w8cr/S4PI+kasyW
PB0G3CLS6rn9XnUtAq/mD/Byrj65C44mbb9HYwTAPqeuooJbfdQMqItIN7QpbPYRGqMfOTGnQVtD
VopezrMLrHTl8HRDyUL4OkbcumpxVKzzNXl3x26caDG6FeOwKSklyMIIOypWwDyGmHU6D3LBFfbv
vclTytdEyFdDH7Q32866t1/FGLJacV+d800Zyq8WqzvjDhbQ0FM92ipXiqQHy1LOLw+1Wp1Klsn2
TGoGlvG2KeFKhWnmlHhS51LWQoqxAomvNU3lm4l4tiVgfJnVecuZe9R0bW2dPfDNNvZ2YbhrELrC
UovF7949iYW1KlLrmbJxctIvtjneWVJig5UFov1iiBxL+bvEx9FCRPaw+0Ay9mCjCJAjuRtHMP6G
fpHM6bFzTBXZ5ib285kbE5DmRIFkMfw9g2XE6sUT3S7bps6uTDcUZjcbc4xpF/f5SCvifQhOwAEp
T0plh0EiBkZv5+tZSgrDcZ9iNMDOyOSTB8cG9wysCtNWUcOZvb2z+7vNpI+rjjCbMuDb+0Etsrgt
oV0l97RSZ97za88wArh6fymAKA4jbCiftaHwXtnq/96PfOHgRU+MMVK/itETnic8rZcq8DSoHEdM
Prx5B8WGXh9HPwSBftD7pC6cbSy9c3Vi1hpBmkmw066hvldUghGdm0DNnYzP7dZVzEJ8ulW0ljpM
ug1jOxAmTsswtKAUExxKMcmAznV0cxr/+IF1xrZoB4L1WdCqwbDKeJEGNgkuDC59xCS6toMm67ZJ
aefdJBI/fB3iYsZSiHKezDiz0Riv5DJNyigs6skBmFUkbFdfvu0FWpKif6CEQ2YaZWRpwLqmO/2i
CWORFLCqtwfN24E8exdlfjZiSYL4/Yim5wdSixCSib0c7x/EC+RX7iW9O2B4r8xmGXCHjYeTztuI
Sm1p/6Yzj4ZUBfAGg15ZL87OqBdvxSYoUng+ydW1ZJYKZ8UrokGj21l/4RhTHUYOOZCWVCoazpVs
J05WCikVPoyWw9JGMhSwtvuhQJdwdranVPT5A3xiCi2EZBzVl/40poNc/f91Cb8xBiVe6XteEMeP
FqMAeqlOrbkkPy/UXEhc+1UeAJh6T+HrnUKi/Roci52WpBWzPU9KAasUJOoytAU6ynF405GcxRb9
IXzIV4fWGRQd9ApgkPKIDtkjmJ6Q1y+y3IuQ+8LmRnPffdVyU2KUw8eculF55ZcOtHjWF4DNYUsI
SeUP5dW3QbShqONufPvVg+EAZ6wkFZwV5EMKbffTtHAjbHFMiXL+AwSlBDL1wWrdSnQnOQlthJTb
nQjH3WjtBgMicADOSgqtM3QYy7Nw5+iNfmAOp5YEslQwVJdcYQyzIpgIVO7fuxOMfhUaesm5Xt4S
ro0BywoFT85rOKot8QDtZyAj/flPFeuMrZjPh7H8V7A4F92ulJ2t2iZrK9kIsqAlncX7qtvmkmXz
d5Nc/7vbOWhlohxm5VAXKSmaAQozrSoflZQ6Zy5CVli56b50oUs6o5IYE3MuWAqA/Syz2nHXBoHM
9ntV2q49OqQTrPZE7IUSDEkjWkz2JW63dCxPPc5BbXhY3tWDH0iEjQ2YCFtnMi+tn4n3g5KwW0+k
pXLnjmhhIBFKL/+LzPXBT5uItmtaWX2djhtQgjw4cuylYxFULZveJoMKCpJ2WPWnloqcbaePo2Vj
lEY5yh+8T+8k3Cpu1CpBYLpcAibxTUV3f02ttSQEOwhuYPaa3Uuy2l5DgvC99W789wk2hyMBO86o
sKoUrkB6Tvpyfw6D6O/RxcAtbRIyTU8iw2xFCHF6MOtm5XcQNGuvcuoIbCYgh2noV09FFg1kD6qm
1gfD8qMsCKFgirF6z2rrQo2PN5s3Jmy1kbF1kaCCmVow5dAT7zBVQBHyOvm94uomdNLRx50pxc1G
uwZhPuOaN0cDcmqft2w/E4DZzQURHUDwvUXdiRx4TfYFm+pf3geB9XOhbDqtBhDVdcClvNYRbHq1
yFoyUKEjqczikNVZ2WV3NaD7fiyOUJNa/RoYSZiFMyD66jPzjLvCVC9aXUbzlFELwCnYNDtclhaM
s6bYujjd6udVSIHBf9q86wKiZIQdzNVh9wOKXJSE3/WZFXtGlzyTHpZfEIRSeT7nZgSC6+s7+PDQ
d3wxyxFICxfg8CFZXWFazGug3JzEV4KSCLfuB1TyGYS1PUyj2dwiu748mbSR5GLNlGUDQynS+85Q
YJnxOLdWTIeKOJKRkGkME+wqsEI+OiGE9te2gOtw2Dc0moEX80yebAEhevtfhsXdaOqSSFSzxsCn
Imk1SvZJTdeQsIOiwJOMD1M2zccSXA+fzvxNzZnyJCrjBPbvPf0jg5zCLlPtTEi3qGa+nl+8IvHI
9ValbFx3QsNe/gC18xSQTtmX4c1hZiBhKOGyicjItEF8LcWuSyznEKYDCVCX9KV72vh5sfeYgqDs
ejRrDLqzKsTq22rh7hpAdg04ibZmfIURKSS/FJvufybC3GvGXSGcsfjss6QVeI2lkBlA6V8EhTwd
w8M3aVTlZadL4h6G2nNXSfuUvF+of9Oed0KjuLy2ClIFqv1MotapQ7Rd9/T6FPnH1hOc74GlaR+u
rsx7ZUn596L36G47P1eu7QPxi7NT2FfqFk9uE2qesLZwIXJe0sEGzB75x9pcvaMixzyNKLGutlvV
hFPfr2mbeT11k+e5Zwy26SdW8Fp138yUe3PUsD6n2uZAM9Avd+iIOM69+e+Rf8tjaV6RFheiO7lE
K1NmPNQj2zgo4JyAHhE6I9Nn76yysA5Jepcv2G1VWcQ78jBi4vEcTbEfhFkp6/WFeBqllZGyr3Wr
9zh+0ajvfIlVlrHHwv+mHgX7Ec0h2JKTKMZnOFJ8IikFRvLAC/KoFdsqv3NaWqY+JEi5z00HdDnh
PEyNIh9ttw2WKY1RlEPvfdJSuuS8ld0aEDIXFS54AxDtxiIEhV4oxt04ijphM2BfBGFVZtaQcJGN
+r7ICtKM9DGefBwEMcKWrCOrW0wVZ9i4rVXkS7sSVUXGAFoqcpoZKGxH92YUkGW19CRKU2VYbf27
GEJ0RRK41IkmLdBJ/q0ryjD9bGJXEbGweQOV3wVNp/X+yHodSU7dGO1ycTSC+4u+D9SauovPZnqW
aZIoaRE5Y8jw1soNeBL/XWQuzj+UejXBaUIDPKDaw4tS9fzqIc93tgcw3esApPfzZkvXx31EiY7W
tQZo669cyeVWl9Zs5R3b5EnF1zTghgfWJBgEFHt70SdlMy1TDlY7z0mzpy2kllLT9pkrOLmaU2px
j+AgJOoQxrivfLgINN1n+6JTt4R6huOGHfEB9vXmJvTL3Soy9k8LHI8YJvDBh3mW90gsoXgQZgvm
IL+pBSPb2LQIF34pnDmpN7iUi9wc3gOkqYhamoQe8TLhuTQ6i+R1t58qNbU80req3PRUhWG6SG70
Pr1rYgy8aLhc9ItyVBrp1GZpoaM6j1IvQmGkcpa1FOSVxH570brv2A1BGph+xK4XCg8k1/oTK1n4
nB98e5A+KOU5wZ0UnVNAgVvapjEKSXxGJ7sFuB5g124Gys4PMu3Rq5DumEO/st3/TDGrMBcyiv0r
9pRcdQgFaDEJQGFpYq5ugF/alEsn5ISKJFV5oSCYvbd7HuiL5Vdu5Pszp59cZovx8Kwr7/PzNWZR
dzX8JSZvDYcg5hfImLwJJ4K+0bJaXd9Jw2axZ0QiC3HSEZr1+rMXGB9h6f50UIGv2RrMhdENDrbF
f/kjq1XR6TUeRIpCKVlKXPZRfTX611e7FMkedIP3uOdD67Z/+6oE3obW8k8bJoZeq8AW0Cip8gWu
ZbB/H6JVyuYFa/T9ZTcnwZnhhm3itBrnwFR7x+aPHI6k54V/kW+s3s02uaWsYo0gtCb2Tk4JoArp
h+O9HWhUKQ8QcizRtfmVF9VldhDfWU6bJIOSaQOrLswh54zHdRutslI7TLabCISPfUUPhyEp2HiC
DAYrdYDnPtsNCujxWU3TNSGOTXSf/snl7SjAAMNVwbq5pgoFcpacEwrlJQ6Nvkyzvvxz0Y8K4E5Z
4m0XAgvNpOZvPUTj02vGuowjT+H714kjbeXIxTOEDYoRdBtIp+ocv1z0him8mbFKdcUlRSMYM5Z6
ytz4kpxfBBo8jWOwjcT3Rm6wG00a9MJYTAGlkS908Vx8BvUc+vXqB6puoLVZ1ul8H8vzWOpD2yl4
LnCIu+01FzOCmn4mH1AyckYe5hnjj/NHG9fV+TUp0B1XtFoSAHKM9RkiZXEzX9rObIdut6zWWNGf
6zFOGZy/hVx5YXCg/3uNprJEAJvdtklkFkwbfwRm3ollHrdnCej6FoFQNWHr8WszwktwCKXwLrTL
MKm6a6g7l4X9BhwlKGi/yNt76wxoMmjxoPja+hcAOy4E3M3Hk2RbFW//rUB1NaegxvzOo/kp7fB/
jjrc/fMSauGARge6a5owWHaLgS8ylCF5oKmtVq4166GJZkGEZprOy17SF1kVoQ5mp4v8btWuF5/q
2qBCg/Q68PLxYvzROD64J0IwZf1kSzjqj2eJmzY7wvmaJnAFR1Hxsw+zM/NJwSWvxQr2l/dk2JZv
TOZd0wRQi2rfYoyJG0Y+lEXxfoQXfYNXrBExQLpSUK8wMuX/zGFEvD13+Zh0iIka37bxWCXfmRlk
gf4o6uKyHU04QYt+ZCH/sbKWL4/tCSrmBKepqiLw3wlHCuhr9D8fYfjZkbVFABtfhnI8h7yJbNGV
6JvH5fzA4KFH9WTHdqUKq+6SrEyb2mkMgfxfAmwsYru5zStKKXJg6e69N4d6tiQasWsjImhdKZqP
deqEgt6l9OIux7NWxm1GXZgxIfWDlz0WigZDOqscuXv9zJInxB3e2r3wuE8G9jQ4k+TPmU5r6ugZ
ektRNS+5xn2+w8jxnQacfXY9UBjzZ0kGr4SwEeBjdlLbHfFkfFC1R/dSkFImrjS9avnLGNuEgFCD
EVKgtd84lLwbyneG/tzMMstPPl+1IghhB7NubAqOcajAMkjjfx3afpVZ7ZQgI1jaAdAcgT0ZLTpP
7r2X8D4IuU28jATd18MVo6boN+0NFOiVSynBPjsONkN2CYADEXN7n783m3MLbxbRjhy7EXpNyAXC
q29L50cUH6YHvPgigCKvN5gITdK235afiKxuWxRjiPSVMA+bAGeQoFnM3kX9BOjYbsbifC5MpsR3
tQ1MF89ZmPyOAAflWVFDVoVK46Gky0zVwYUc0S3qyaOdDehdUm3X0HenZrlcDTRDU0HyRsuJ2UcL
6Fni3dsGNoi9K2G6cCGho/Zumy2EXF/qjMjU4De2aGXAI3ovWQKcWBMqjS1EDFHLa/DIac0qINvL
RDB4uK+XQMAkPKBxlsX572wCOIVjWFg9NtdXUHh9XXfldBqavb/B4+u8yUKkvs6bp98vaOddhMXI
bERzHiFGCPYhIWTJE+RQ/rrnaBaywPZyEYPgZG02NuUcf2DLOvnp6luuGDFtIvNBzqy97dIMEAuy
f1hpp8NEdST/908oR56NCPHAOacDZTtNEzQlv99EV062l09fLoZmwlTxDQw3qT7HzSW/yjhf/YRM
/SNJSLGmv4CpPC/yMvXPsWI9TqIhmqo/QNF2RoNP/emsti0u0+Yj3FRQQ7ix2Yc0FQSBrRyOEW7j
MGR+r9GpaeE8zky0hoG9pujGyxeOabkIjOfy258VwdGOMkGRVkoJbm6xj3hNYmrNTzEiHMKvcgIg
+QPc1zETqPrOj8rRennaq2LCOIC9eoJlKZJqS8qOVIeC+OqmWulgq1cFvqXNFD74ZKe7uMQ+Z74T
OX/BkO9pujzkaNlQRfqludO0/F94yu5AnjFg1R84+5Uo2O66ir8VvnXTDBizJ/ZUNYz09JIGhR85
H/HTsZF0kkb4UwQIFX/mHqcZTrZQ5a6lf4U+sxE1uXILHuLxwsjJey1Ya+qPiHP9VlnXLbeLBSTN
fod984SMW2ZBhIU0qYY8LPaOlwcfD971aqCEKH5j6R9OleJGBldqpKtBmaz9eZoR6oJiiX1z9Nir
GJoQ1OnqwYrG+T7x2ikuho12wKYQBrPrgUz32OImTH244hUjXZVBqZJRHtO54QHSR+B+4TkX623P
4k61I2imjxvtxTDaJmctwosoRW5qSlx18wn7tTJeul3jAOor4oo3ruloc5G+rAGMz6di0SBXajB2
MAQeNUSTA4Ny6Znf+i5J3+J4RA6AAlWrVSi5/wWR8tM3B4Y2shW6aMG0jVFK6I8q0VZYmIN9OnFS
bycU3K7LUX4oBw9T3B6sz72DBourCdMTwlNRdFL6KxuZR/QiV5NWUVaV20Cu9g3P2ZGVLYkVm/SL
zkqCK8+9ZidI2WP0cd4tlYZRlU4qcPVjRkaIOVQRoyDTFYXSnokM2GeepG8bfjh2PsGfzGfgyb4v
errN0JvZF30/1tEFjshqK9xnq0A3RQQahN435pU7lUlLsTXRkZTAmEyMCXkCS8abU3NWrvMm4VRe
fMudpRxtLzURO08jQ7XAm6ul1gcrdL1l9izn0amusEJrtytYW+xDeIutHQR/tXUZ4rjx/IYQmtET
WbwaD4kYIzY+qs94hwx6DZmzD2h2OOIIdb069cAuIwTYBv5g1M77QvG7EyY2dNuv4ukz6oUKHRZG
jUlXBnLmVBDI7gy2/aCD2z7yReqKng7Ic5+iZ2dw2MPN7znTKEGqQsimiiCk/rLmxGJCim2zzFIM
YTy3FyEWZb+4Gb0U542jtfOzR8PqXVy2IUJDwEb2VfURkyF9fmzGcbxW0MgNrf24dTKIRHK8kJtZ
OtrU/4GQ58sOJPCkGDc9yK5RP898/8PkAr/kkGUrdwrQqZZZBageiqaAgAiKF58ZFx89XehQUabL
BoogsTapq/YBcOVYlApbHvH1MRqy6fqCryV82L0r+bg7Gw8tAg89JFqlwP4uE5bnwhvGzfFxxhWn
DxbrWiZ+w5DeyBa4PKvCDgInY17UhNrH7wSlYVaC6bDIcNxRGZvrn9wi9LxQW9yw1wbV1uWKUi5c
hWkDL2OOChG6EuC38ui+9LnouxJ17j6vTDIKiBuFiUBtBYN9uylpkNiNj7J6D0wlWi2Dwxm6Pbaj
DjuTfCvOn3tdu+vqdU0MdbE8ToZzxyIUIm8YTPPkMx98YI2MncJlV/H5HqLGDGL7jszHkrsPwz2P
i9MXSr1uIo8pQXQ09lJiLrZswQ5A6j7C383sXFxJBKbgP7R2HmdDKOr4Ci+tCfep139UJLxf6ETo
52ekVxGwz1Yh0UDx/GcIKcliuufCyhw9Zs82oejQ3pklx6g0QwPUmYHQNgL2OkZ43465Xg7jCsML
VPH1A6IQ3SSl5sivEVTuSWylfTfYSSbcqCowFNa1HtotPjxBo5l1jxE5gmaKCSdxOTocBAGkUw+Q
yGg0vIgtuaixCwXf8mvdw4PaPoooswju/cwestA8j+HBIycOFZ67lrjz1FKR4mLcrEshKPGMlkHQ
ya4N9/19bCVSmLEXRfZRzNOaPPEenannKm1Fob5/S8B2zFjC493L2TyMzCHfv7OEqz8X/RPgFdBb
BLIdyUl4Xg28Bu7mob3ZdRYF/x6R3RrS47AwupqXhQTiimqzrqnfjsrWjt+X2xAz1pNnGa5/38+o
5xrgd0gn8r+eoDEDhkaRhQkJvkzka646fFtOZVsa03SFTgMKexJE1qfhmr0EYlFm3XbyTGjExnnV
Wt2vVkNGu2ldSKfkm7j/iDfmS1a7KutYt06wm0dE1v7G11r79Oyvke/0bmq2lRKIK2KRXWlNyfgr
sQjyZ5OKM6PFDrCRFY2mDfyqHv9hKkP+OEe3+CaOctUATU9rSEUvLYh+abizROmxGWo+Top1bItg
qnlwLwPeC0DpMpxmmEdTZ3oET+CbE6nD9HAwKugqrYiwzkafZwq5SuapkOOisIjahbaVIDYFDbo0
zxAbUSxAkqHdIfr+YAx/BYEHJBCDzmh4LH+rFR9aV784mjISUumCTro8c7Ks0a7LdrFxvm6qarK1
v7//RZoiJq0chFKg3ym9qMIGBlUbzG/e/XO5JN8CxPzmAHqMTHePSpzmpZ6oNtwHtHOkrplD8lmg
xyPp7xmp0m69jaVb+m5eO4GT3JA46p/+pGl+a0Z6vGIvTucOG/Xk5q+/Dh83Pwil/1swZFNrhu3r
qyJmuodfBgH7/QAjSlfKdz3Ub718DCx01SEBkWzZg2jksFmE6vm3mjL0JyyTSPNcY9pp0oLEO8IA
j/KS+1xcoZRpvSCc+CjQHAi27EPnQMMY55ilROVZ+ejM4STDEcs+6F8lSDgma4MJCi6dRlw01P3v
0fnI8L18Bb4DD+y47/QlmKF1ZLqrz/ttsMdZ5ihjpEsD6EzPSqbu/kT/bIOpUb5AAlEgUeKdS3Xi
KyrJ5rYig/HF22m01wso6Uh1+MoInsNY3Xx5fGrF/wkIJNTYq9EutUPv9NMbvkSmeP20vXTC0P2C
1L41RyUqsZwSSJi9M+egHUKQ3DE3kIYZMzQrxaajUd0SkZkb/BaCpk61JPDWvajbBesAqq9fypXz
OuhmYsLEKVy8YDJamzu6GjpItJswSSpB2+9U1GvQuuuwuNLzcf2XyohQ+sLC0Piap2OpOwQ1pzr6
N0wj239gimOE7oIvpLDZENwnRp34bAybCjcdZhsRkNr6ZfHVDAU8SX9z9SR9ZTATv5cq4REBMxTh
1LSOW7kV67dDEI4bC3NJxuFQznvnHTBkCJ9uutcwBqhZvcx5Xdoq6+ABRRLCbvFfEq8xU2z8N79V
WMEg73b2ec4mz+TbZZOPm937Su2DKqwGgIxvriNqQFP9FWwRDkupPF7DAHb3PEwX+JfdOIbueIFX
OfV7QoBUNUFqZYKC0Oi77U5M52Mh7n/2OBVt4LZDiWqfC4j6Rr+LybXsA6f/FW077PYy8Qm5U5Il
Ca+/WUsu6D0RnOX4nUUrjYG4c4tDrNrEIKcqFS66C3vOSx+0oPrjbfQoFeIt6VsCQFjTi7OGQTF5
+dgfnw2soUv/eAiUUZ5Cu/rWHgMKlGDuPKAwPLtDEno7nJdoGgyjGzqXFuAMBhpXaxyNIovP4Xfa
sCpCjJq7eLF5kAYd9YBK2k2KR9kgrGMTnm1AsXypNq4dp0mkQgUnGfLJwRIi1qBPLUi88mk1iuyN
oPYiYS4/6c4ZVEN7cUhngPuYI4ps0GOQjG+YumaDaUYGO601fp5DHVirn29blZEwbjOJ5R3XBdRn
tRsyUr8vPk+7sNwBD5UIq2riDlkkqv8lIyDth+O4uZuqbH2LSs5LOtwUpbgchV+MAaHD25X4aV1Y
4WNaGtjiRh1q+QMt18LLT8SSAUWEnBncnZYhqZvuLwfKAvlQwWfae+mOgu5dlwD2OdOUQHZMKFsD
bm4uD6TdXOr6DSFGGiurRz9CuBvaySJDwfNj0TROwwH8nI+s2dUd1ZoaQXftr+fUGvnwWb1ZTcBC
bkIZnSs2InCaNjU9Yi8H+7YV0SBzxvfz5pUODW8f5SEZdkGhPZ4VqDiZctGNP3MtmS/9chbV/P+o
7zDUK/imnFzam3kqjRSMLyjc/i5+XA4PUiX+eE6h3MDsV1S8GW+NJwVhJOJ93bQ7iNapgR3Oa0Ee
X0ETXNb+CHvdSJEQoLL/qMkJHMYF0a2rOUsfrUoAEzkhCKjMhcdYVY+44CzdbgmquXoLIu6cHq5z
8YdVqLn2ZywjpL751RV2hyOwDoVfSZgb21Pok0c8clMxSvbqXyZsYsaht02hjw8mjtkFYw6M7n3B
U6mDC9Ut662j26cReMkpU/Ij5av9EY09ys6BRHupnhJ5BXzx7HAIPNjwKLI8rlHHjbobB9SeZhAo
g1FNt4ottb5XsZVjENLQUjkSDwI6mIQiENViE9z939KgxyVjooNEQ549oAd8O58CqnJaO1frFwuJ
hix1KvLGAiLVAqLrUni+6oFLhx7vHSV4ZeX1se1lmWgWjZKba1Rp2IJlszSEqW+abkvIytuLcV2A
kioGmD+RUNmIT6CVMoxrVzO1qRnvWu5J3LJd+RWPXXeGDcmMpuyMwGTjg7MLWanXD1LgwedeWi8l
50P+s+6Bc6p7/jKS3XjnawK9K/suAEL3j0WH7hRE4SpSPViuxpETvuVrapr4HSay7UmeYnRonxZo
uZXeDnPSdQIg7obTv1xJFRtfwOJ5cZytBifAxbmNhFPLA0AXDzDPA4YACbR87cOKVCHKt97j4hyz
PhrS6HMvbSLCtV4Xs+EuIBHEdWRgu4xSr/LFcjrlacXcPC/fUtRatx18X7PqOLQjcayST9X/I47K
kPp9Mi7xLDAtsGA46wT2ru/mtUu4MKsJPDbTVR5K4ZLTnXvwzx3eK+hTpNtAgPLCQuezrO8hqt1t
R/OlhCgj0DReEKzjTsKVUx5TqOMh1gD7VwdOGFxUlgYW3uoss9yTiaBTqmOeSoIUkuQE6Xb0MiTN
6i3hFot5p2f6Nyt5mSJFmS/+OlU8d7UX/zfeTowNQ8VjpsNQEO+YVDyRDI4dkvHdMX8r/Yjs6A4p
r2ImaOQUJgkf15emar1z3fRisQVXmMxb81DD+iu1mbZHDqGien4KrSErVb/lr8wlm8QAiTvOs1KT
2QHyxfLEM+198WrYVs1V2TLh6g2tG8+4x27PGxQ96dxMsBbTsED/JK69x5tvAYNhbXi6vP+qccN0
8zhLIuh8N+Wh8f98K4NDo2R/67OVfr9AFXrebHfmFQsy/QekdqozZLXuUR2tyDeqHDxMv3OCn1He
ZPcD5zzIsejEP27FrH8nxr2X/LC7lAllDa7sVmNlFHZhBUzrcYudg6c//5loYzsDK0EuRts1JDlR
mtce/LN8psK+y5gz+Xwzvmr9t4AG0KJOnW3fFzVDt0OT4zN1FdnvJtktCQdY87S7dzG7c+3mJQrS
MN03JYPsHCaz52QtO9m9GenS6PyNhnmvaNNoYne6qdOuvIAbpTZZsyTBliV3QI5tjqye83TlRjKl
k2IIjDBpV2MbK8uZWR+jYw3kuUCiD4D19MT0f0QrcRkXRyhkx2NbwSjcSGMJbwKGt0u+JnWkJR4q
mai+0ArzAupOfaYtAUi7TGz8uTFZSIiDF48P8lmv93Lysw5oxcIdFqWOyCOZcrPXZYclkns/Ls+a
niYsdwmh9U+4ZEv+kIIuCFM5ju3QdzJSIIZzdjmgawhr73m77WBpmsHDU2Dppi8/jiDvu4Uc5srK
Bpi0B0kq1fPEoU5Lk3QmCnHcPCX6t0acwJXlQ+3lR+819E05vkoCqac/O3v26eCJtwkvZMTF40Ws
8wPxyUIUV9oM1wHBsAUXrvcEMOATB6r1bY9Hw1wFCtGbJzBkYB4Zz4JqXCB4OSM2H68jf0d2y6ys
qGWtnqVS30As+YV2sWL2W/0m21rL1WTaZksi9aRp7qWWdBMNJZq3LGGf4JNE6ZAIyTBrg47ME5FY
tTZ/plwAP8bsQKkIZPRl5tOs8sGls3ubKvN2vNnN3ylHTWP5AMOapGt3EeveFqrXXZDkTfbmnTml
jbT2WKIWTHrGwMm9QQZIy2LEOqdPdnUuHos2cx5UuC4C0s4Og0dLrjjSUtuWH771xfOfjK9eyrcg
XCbbtD+idYiVqPGvjLAWHWFpBpY6ExL5vNSD7uDs9MbrsOW2v/bK5dVDAMV12KtO1paBWKmS+w8t
QQQq6oaAsu1y542QFTzcumLrGRyByOCvG66UobfWGoanagrvtiFgyxo8FPaNtlOYuu0NNVj4A0oL
1NOSY4jUifPu/Cs2YB2xFsTGC7To1MaI+KAFpSqlNCVjOUZIjCY+EF+31scFiZQzyM4HtA+G5Rlk
mZAFP7BHs4IMGsSZ8/Xw3PO0dS+r5z08I7f1zzoha/pOEVDtVFi0Kaw9prmiBemBm603V4iP7+et
CzgIy2eU6mwuEwU9ePwKTV9kMmyel3246dt2xRG9rVQBYIeQvHHgc58iLBx90+2U5kDVm534KWit
G+eca8HFZL79LZcBC33YTzwbXbTENQ2wOBlben//UlMicXris+yqZn+mjgNoT5BqQpqrnzFc/IaP
DTCtGcI4SOXBQJRGbD3KfzrqbbYpmAW/PyAsOeB1ya+Sh8gcm8dtKXOxbKWivWlg1ST0hIDW1K5g
JpWSJvNnGPxaHOxfFDZQG9kZXU1IjEhQUg1qYoIdXW7EIBC443UdxjlIRzXLxD3NDhk/xDZdGFXH
GpzhZIswCbnexCd/eirjSBOF1nMk66uVFfq0ak9jxRm04j+Uo4280+0K9cLF6g6G1iUK3M/2bgTA
Mk2tJf8+/vvf7JZ1sQ69addoD7FOwRsxz6wBFWezT3AQZ6lY0YktMeNBMBtueZ+7HO52pNNtbH0F
OECpEnk+9am0RUEYM2KBqI6kDnkS0F+LlZXydl5V7eKCVAdBXkcAcNSxfco507ii305hEA+PKw4S
IrcKjIv0S2ofS0fws4pzUoNG1KvEzM67ZFD/NRZNBAQNhBZ6SnunwKSN7gIKG2oPc31RjmhHfXIK
rbwxoRdT3BCcuJR7yQ+SEhEVGXjmbISQP6W+xpcxAZXx8phh6DQMwuU18wPYsuoV4fG7o8KH+15N
kAf8ok4o4Sc8wUtTRaxVa0Ak4o8rb+Y4jhlxq4KIX3/IcvtMOu9LmPFu8knKi/nr7dmKN2DrUv2x
GqvfvTg4Cd3nSiSr1iPHIO//SdgXx0TmX3WnQ6yftpGLd68/d64kDn8IHQ0DHSfKiodc9knVLypq
evsM3+Nn5pa4rRF7ASwnxeC8EU9lZcVsrgxW2mvk0DrOW8q+ypWspPI0SCVYFzz+V0+INMXhco05
RVwhSFYRyJMHI7Me9e5xioJorlFDXgJ1A8xyFVCKPvCmpt+KZ08RGhBMLQ0L+dbfUWT+QbbSjG6d
7d+KHSZZw/AStuTzko1xht+FelUnL3R4j+nDD0IN6+27jXzL+ljJ9D7VwVB/vrcpxtL+KEdiIluK
Qq1bUCFfZy36OZdoZnhjMWqFZTzkfehmLRYenQehnCHoMtn8EfygPRXkzlf01szQ2LLcsUVGsKs0
b13VK3v02GVB30hWkgJbND3Ggj8oTShWocAIlMqXXVHOIGb8kdaXqlqHx7rrSonXaB+N30v064xh
6VTnmilqDvYOUSBiXQgGpRiFQm56uAXVAQQN31heq8g9mAi1GfYTWAuVl0lPmowZaxhdyCmon9nL
J8PGdvPulhWtIri/S/7gKSE+YRzydJ1xzPnb9upwFxKlz0vl9+idO/ZP7yaOT7z21gKDnbcpX3me
AR87h/GK7WZKcxtGp6HZZ9fTB4ZC0nC7BcHaQr6BG+z8Od20NOT+ALmcHDs6k70A5AjA2X6U4x0p
1hJJ0Q0flJOznuNadTKIxkl5yhkskXV2fBADUXESVMn0k/cQULin8Xo6NGXTmrAkpDGDbb226Shp
lVM29nDoGZI+YNG/TQ0qePGcazYtc79ZtkWtEnvZJSSdKjdeXJ3Gt70Aoh3kLk9uE+4Sa+qWquh+
FQngVbiI/dpgfiXe5kVpC9peNC7mUQ/zpsBo0TCIbrmUyt3wNNfGQ7kEyTsFIjiHfvUBnuAGxbQ7
I0zg1c79RvSI+qK17GdsUCnZo7rskGwbrGQj3NHfV6dEYG3mawS4TSY+qFtQXpH5HsC/UlJktS3G
nsEhfrv+n6I00gfnkt1noAbYpdWIsR3TstNvJyLPAYumTp8XJdR9SEl2MinnFwDHRPn5oNghjLID
pyt1DreAkCGFU5JoLFZujvHBJUGqjdtRsn7OjcdYJIwYGSsDQVewpgBjuXLebYZNhxswE+W5iooT
7nJRB+gHPxNC5OvokDMO0E0tyOjKE+isy4X8Q8IvwK7rtmWziLxLS1qTSl4Bkrp0W4VH4PtqXZND
TFobLMjT4LbUwPrjkcU57f+3AXhM0rpPwKAQkx+upmP+If7vEvL3RnuyhcLU6IEXjch/1kBPiuJg
yCPFeIUdSFtVp5wD0M15oNqJgg2KAUwOJyhGEB0DDil6+gjdivenTNRbOgVUgQhtvYDuRAka5dre
/2ZQRd+714dzleXIqt0afKMKA4B4YmEi+7LUqzzGTbPyxAi6tgmcAf6rDKozrIxnmDCvnEmGiBpu
QPAl19d2eEHor0GcxTYBZ7zjs9r3FS6IqmyXX13FDkm7ugr7MmSQ7560+efX5ioRYwBNeEOYhdqY
qUkgCLnLBkm43Ie+X7eV0tSk8EdGUrR/3gLA5dmwvqUQ/LPUjJo7/aWzfCoVNFbgjESbFNrnEofk
ldtCvVQN5iyUxKBcHSf1e8tXB08Gko14E2Ykk1pQjzOgT4kVkL0gKE0YQhEIWMp+/qdt+pwQP7BK
V1vCCdBT6pbgZHlF6VtOEZJyxd0h0HkhEmSwsHYYAmtf/AkT4xjAz4yboNRj+IZkoC27f64kFqLG
NSy03YjifxwSvVct4AzGahEDts1MEGDTMHYNn66Hi9x5XumNOcoeWLsnq5Ei8kEf9+keVN1vNTXK
aUcdt8Ktz0J9Vgqc7dp9nDCHgCKB82VHX6oKuGe3IagJLdMrisoiHunhGOI1oxmsjhlpYRvjWTSk
qK0OD4HCTMnnQVV9SEJ3J2nDJV0EmvWtkfwOSqFmgg7FDa3o59JoNZlUAyRAtARIOMo4dtro7vp5
8C8DjR+POcHC7mJivYjNMMzx0aPIoY0QYy2g5Myzp5cL+076InGdp8fvo74CLI6XLoINRT062vvn
yZrFxZKFREmmgmszHxCB1MGJ66yrTzmeXNxOtIsR22EW66EHIfzSAtE6GXpC1vDZx0BynJPgdUF6
f24BfdXstwlws9FJq0nc00FeDhcFhyARsSDAfWuJbSDVR4nJ4vccgcCacGNmK4HGlf07T3oZFc2z
n5GD2f1p0eLuMkBCnkE6NSRmXG6+j+tP6fW6MOGbkASlErSKdoqP9GOy3Z9enowRmImNaFz8bAGx
rbyEU+z8MMG3iM5TG6zhSmS5btCxpTAA+t6cmZXfJifu6/kigRBH3o8sQ22iUOEr3SCJT4dmZeRe
U1RY6yVNStrZ+5dxVJFBqvUg/D8bygSrb52z+JVplLSbPzBKNF+f4kGt1iV1PN265wHzyQxTBmh5
tVSK7UxLdHCSe3XCf48VzbaoZXFnjUIGLftjFm8GR1gQhty0P3BMfJnuMp2CsYwV//emsVSGSpVz
aaNRVi2c3SRwUQf7I8ndMGCXTDoTrIiZyo4Kf+gJ0IZWx7Eu10AGXkjElCXC8p+WpD9nufQ64qvj
QUPNypMKCP3R2UxTjqV0yz/3Buty+n2Y2R0VIWq0GcvcESVv7Smb+7JfHiW0ZRDIkHFWldhfaE65
PSfJwrovTkDcHk7zPmrDHfHLcc1LbU7lqjyKtOSMENCgFmFVwK0LIYAG5M6J00d5gFURf2su1oTA
xhwBak175TkvnfpIGWI77VODdbcU/c5j/vxVDQwq3vlOVKl3nCsKCDq7uNahNeOK58vcU1p3+N6r
mdLgD98bbi7LzpNJz9HS+QZ6hftfI7iR3CCaXMCfK8RK8hjXWf/qH6/wbBftfHjN5XZi1sfq8YaF
ImVlpK/eNv5rH3yKAcuIrUfZmxAyLu8dPC7cCAotgUum5RY8KL7yo8WuV5JdhN8d5U9Iw1UsZ9Xq
RlDPTRbG9ea5SuQVNXj+zBWGU/R75jFIbBkNWtoOQ5ceZelJOwjr+MgB1O1cSo8i8i3l22KgvXbA
TM1eUZJvuDrghtsWT1hPQ/Yoi1Rt1Th4q2ZDFh8kDj7Cy1M8YFBujz4U7zlf5V4sCqflrug4yrnq
qKtFpZvyoNIfmrV695xC0dzAQBR6X8TzeQ4158a+58cm/R6tORDXPBCVgimM9Ue6cRc1emgRb+4H
K/yEbB5dTdvX3Xf18SHIz2WP3/dnvCNPCb67n/8biyOGys2UFDjtUd2qXO/f+AIH1B+zU0Qdosy3
dSppp7i0zBYCYgFO5Y5ZfXUKcY+LkY4hJ9av1RtyNqiUBa7lDsGtu1dV53W5RcLwcb0usj3/dUds
4RR6v2qiIZmV734Q9VK4+3WX4eG8mfLYuw3oCa7cqlEMXcjmIPTBTFBNt6pqrAFiGJqXDlRBzyvb
4G8nRKsGutPSBpe8WU54pF08EAFX9ku1jHlT2wk4Ko+OYoJlL48kGY3E3dXCvpvAt8HIkDdBmupD
CGabbAz1mhGt5nEBedGkdESbHFkDyMEUhfiHqy8HrT7g5FSoyfV6udh8YtNy8RvI5EspUsw0dMyH
2Sk5dFgTvk0dq/wq1csI4ev7neTUqIXbUsUKitFUqm/VWcdhkbAKd1FMl5OLbZt117z2e+8uXRhI
kf8P3f71P2c9lq9RfpafYxmSlOGHCFfVKzZ0Fr4MXRMcNYPHwgylKVfvzBVchMrrJKAn9yxufook
7NrZn30vkqwd9EWXwygk9MF6Lgv8Qrt9749zr7guk+S7J+lNQFGFy3csNlBU/Jn/bdjqoi4PDqYr
73x+B8gf+Wn5vQ21K2rQJkc1W81lw5TXwfPye39Oz2YqFZOjQp4vlxBiXC7uWOm5r5Dv+kduWFUa
rca0yxViAz6/vhlC4+3XalOgHPcUhAORyszOcxYYt7xa/M+/HtW8dMGmIcVYBSFQCpLqwEKy7F0Q
hG1c4NPKUvxYR9uOwBuZNO85ZWJwxfaZceQosib4iR2dTwrqmtfiTLmM+Ma3MlvCIfp47CCr+An6
AxdpSF/+1R4LqVYLLHN0nvGQS9NhKtIUxdtCczGMlALTNJBIzlzAOfufM92+60Gf5OuWGaKoR195
qgyjxWKnB0RbuLqgD+ut4KjeQSh8ZPj+8Qss46UZ+EFlgTV63gY5/9O3yCmekyqG/U+5c586ukz/
ectGSizwF/63QosCkIwLuwY8Yc0TOFYLsWlt5WUUZPSUcfYW8alJky0d3GQ2B51NCmVJmyc02Pyj
2Epgfmhma126hUrwpglqtGnOsn1jezd9Fe1ndBgyePhVnpKp2DAW1aJOhoZZJvQqwLzXa5UTWAOz
MZw+ZYgr5JQ5xUjoFL3V2qCais+OfdE6J5nLgI5uUq9X9khCqEd4qsEOz4t2MckbEVh2ALa2IeTM
td3Zx8AavHLc4hmB+xZbr+UPai/hLRvz/cApMDrpRqvBvSmifCgSy+ypMEo27d5czsOx1dcgyaOF
HOMTiCkcKvevgW4va6gbahZLNttoxRu2yIECMZLhFU5IGwHz2xC1Vt2p07JolIR4rFfeoTxZvzEl
jKGgmyLDjsTE4yVFFYGbPtzEJKOhJvyP7A8cLdi4qCj/Etz/JC/bjS4s1WHBQUUh1QQH5BUgys4e
CbEQAzbML59mLfEWoKJgwY8B9ws8K24Cpicqsl+u2AeSpaA3WECPzGZZwt8QDy6+pjIgSQYFt589
3lMf7ETAMGRUsabmH/LYeBsN19flBXLY4xw4aOamkupS7ceqTRFK28EydqKToBwZrXCSbZc2DWq0
tqXdp8jM0/stC1lDSNoAnvrb5y20iwa7Tck/0SFWn3fFwnKM62Mdtlzh4IGAuXEKFDljY8mAyufn
1KqYVSHAAPVsYbtNhwd4nzt5xKNSpGRc0rt6Rwfjey+aF9xRdz10nEGlYJhQJJV/ohahpI6AgtcZ
BwXeK7OEEmep1mmw6TTygMntk+qfmz1gKCV7n74RHQkqQzTZ8lx4GXMmqTRBG+MdoOCzL5/5rj/s
iOIm6c5uUp//YI9K0Zo4s/mGZsjlwPP45daZ+7dElLraxozj4+G2KktrxlXatEuocfZZbzByeCFG
GBESrr27GJiPKOUG6R8W7cadcRsSEmhiTfqqAcdFuriww4fDPHlVJxnYknyQBir+xQOGxVJBcUoS
WM34FtsNQfnw3LSnKyo5QwslxoPkZWPQD+1kYosu4RWJrc959aysYrc5JcCsAecLCS9i8XPQiVPP
ug9BAYMD5Kpzbp6ApV+SNrjeL91/IFUq/y1xlQ8mL0DbdXbEZhGAowB6SKpz3bnoE1I0PL8z/ri4
K4ltbx8xTaFyst/y0alYAYu76Z/gSepAbwSnAN6RmhdQalBP0T7N+MY3kO81iIc/hIbn4ruZrmfq
RmBEPSOWCmjsC7Fktd7Cwm5v8IxsJl9tmdQJZyPda96eUGaS/BUT/vE2Zq/bzhDDAZyHy9J3PEEp
p5zRbSHMmTVt2g9KAvXDSlbKYs0EmBEvnjSjl63BKOrGwhMu66OdIYpoJXziO1GY3YSQCi3QGdRB
qe7DkBjUIxm8dJD/QsLkhr8Dcp1+jn91A463ehZAqaas/XJfe5K670snS4zKvhQSU1fi7/pG9W2F
0FGO/rFpnpPjJPMELfjW/vtG1ffIqV32+FLIUtoh+OnewdXhAz/Ifa/fv9tLe7NOABQjODmDMuH9
PPdc8i3sm/zMWtmwr1q2MvkQ3Etxy/2royVDn6BUGXSathMmvRH8z6HM0srp4VmL6pS3EK7dRk1O
NmF+JBZVwSkAwMoDg8ogh8FxMajPAZWcrF4CQb0pq8WFXpyUapjrrkepVzNwhcCih9N5AHU1fmxo
NXv9QQWl/Tx8fLfnTPCYOoSpHVLst82WbM8y3a4LJScfsbuYYaBmSNq91dXgP6smhh9eQRhVEsFe
PESDjbpQ+p2b7SBHkNetY+6AgfKc+XM3fdOGHTDVbuFhKNR7IAuNOhcQmiyTv6ea8OsxLFfTB6xR
1myxhTz/cBkkZYaqCb/fGwWonmCMwJtVn01zixxT0uBlyhe5avIzvrNkFyriNrqnJMxFhewTYTUY
yzMxiF82FXb6I3ZCI3UaAQniyXUFTWoebmlMuwFmjjFPZDWJJVRVmy5GAXVx7/Glg7yDzl+h9n8k
Qc2qoazHaUhBv/YJycMzXisBDfZmJw1rKgfkQCVx7BhqxHlBJns0254w0kanZ0AwV/09dlUlddcm
MCIZNQ6qfncUf6TspVhQ4UYdw6kFI/gS+aiSm4AUt0N6BojH0VDpKRSJI87sndajb98p/eSEC+Z/
kY0G4Ifu0gsTmLJ/bSWxqrnJOvzwZYb/K5QT+3XYcz3qSgN8GxnlmZYyP83n9rfGfZ7KjlZAYY6P
38+yxo4tblX8xq0wRSwjYnUoMlAVzMHfygUIq4rEVR3N0JA5pSkoSDfEv8AfIiEG+RW611uilnNC
q7/dTxM1keBoLLwrkBeTpW5hFWqrQLlMxlTGQztW9Q8hQY9OihWMv88h/V0l2DWX8fyV8jToCVrm
XxG2i0pi0ZkGI380LUj18Y42F3SmDnuoJtRq1IWx0KJS2WdqENd1MgtAIp3Y1YdMNSkvAAiAqrXy
HslG+4YXlffdz7PIi9atBxq0rS+4DiYWx7hszChKdHCtDIE33q2g+Is/Mrc2sT3hPSIoCibUKR1i
SBdA420i5puQdaWTO6B1ZSNRbGmI2sydnSD/ULdT43fESIvCJzmPpbQ4y/MQ8FupYDp/o26HOgKR
E8jpnJCr1+t41aVd0e1LUR+8HnnTC6L6V/D0SPztd0zilRORnoVKMecNcujYCvTfWG0mdUu1LCMW
VtCGuP5ELkLMJvjY9KRijsNkO5dOeHzandzoPxSSb0rG08lSlGY58bFQwnIiIlodrt3hp6x7xcJ7
nv1X0Dx2kzu++FyHwj40/oGkk9nMRshWe0ZO6nL/USmICQAAzgk19XFCxb1CQsg6C1tbuh9L7ZiD
g7GsCcLuKx304s9nLLW3cayXjanZ9x4oCBuoLzUW81pbWOtFm/U+wnrMG5o3BduggRr+TRxED379
+qx/LEV5aZWP+FMk2r0Gc4EXVumT3FQ3VFM6HQ4vy0RAbqOCW2Xl3HYhjtLVNs8Er4CzTkxbr1aY
lGhxN/jGriFhoFbG+ivdgzdfLdCmVXEIyiKHhk5vgrj36Xfq2R6yGmF3/gXo8Mb+xg799I6su757
5XiGbiW/uSZmoXAOu5e4mQSzntuTMzCNNTpqzS4S7erYZfeRj7bcfe25P+1wSa7+yUY5S/b3e7oQ
zP57XaOS3cmF6xkQfPkx5n+2z9Sx2vlsuhpbMWcqRqJAs/PnSm5TI73BvueMq66ezkHYikeYjDsp
xC4Vg0w4oydSwjI8ktKWjX+U6qD6y15Azn7Unzmil6lRD1+q0ny+3gOw495jPkUts0RpppalcHJw
/uq4WuOeDIPFcYHywS4rQluWcZDTdUE+ag9Gdz7OeToPYaUlknR9nphnwMITjWbT5/vqS81BUpFD
6n3e5slg3lagIawcEmJ9KjRLe7LXj+T+QBAfGosy6yNjZnYaPbE+PjVBsTlG3IRAEvTmghbD8o+Z
JDgAlhETxHQSLLKKoWYveaWxZe5JgOtYhC3hKq3oNywAC7gfC0i8ms4j1fkOsqr7Q+Y2qwbiaNP3
Hj/4Bo1IHFLZMcdtma7Ag7djJqq9Lngoa01EnvV525U+04ssuRjhd0JyqYcpKkhFLjwUmGYf4jIz
lq/AtWReFW+8nI3jV2VkLqw2LpkFaIOyyLk3XBP+hPatKN+JTW+WDo1an4JhbA+kp7TfR1zoAJMH
5VsDCKKlgjP1usOYz5/dfcVr6hsu04f60ZLhnMFUrtpjT9lf9BUpZqEq6CZtjQd96ISJoqWVYXlx
FWfYF6X0F3zPevErDFTR24XWocKNdc7vNX42U221xiNI6ykNgWGPElateVmafcPe1S8STPtpykBn
nwgKY+ru4I/JYz/ZB7BLBXCc5VUWaWaVGBDwLQ+BiPijLuBN7VEgjvNuImoA+ZlCiZKTs81J21w1
bt+MfkqWJ4VDUKde7ziTxtRf1aa8noTuGuB7P1ZGG+rOwxpQQE1NhF8TXFAqtvt4xSgPFQx4XWri
hIAT03TBmFSfb/rlyUhMMLeyd/OPHouP5h9xLHbSDr0PjgVM8xtueW/oM1BAky8PmbZS4eLyn1ua
ApMA1sPvAxPRXnW7j+7p2w0NcMPO9tdbMVLCmHeWGfuXKIC5J/CzxAWrEfQWAwzOMQWCJ/pgP/pV
jwpZELB/azhVl5Wee9noeqRnodXJoZG+or7lbm3eoMDDwGarPi9TD8OIFzTrdDxGn5WQnfVR1UqH
FAI5q4MKUAH78iEoTreK/A3SWbz1cDMazJveBd/Lqv5zARho+zWAnst1qejbh/+L14Y4KWnvhGM/
dbA/EI/vmV2olBX+EMzbkVrMaUZKeNqhc7CGNX69kMQaeMEMbDKp8THaJaSOafC6FoV5DC1WZeuG
laXHqbRFtT5aVx6ai9f3Zz9LKqYWotiVqTguT7usRZuibLxfxw5z4GIQ3Cu2XHFoW+cFmxmn7pGi
3SsPSFx+pyRWf4cT+yBdNlxbQ/OsVj40zNgFqKGW9QMbxhU1NrqQuoqUIbD1Rb0S7Jvc+YdjPk1r
JYFSLa6S7E5mR1+RB+eshwAanN+jl7/GrrD0GMaocSpFrujVw35U+gu7H1UKBqdvrx5Apy424uy2
dZ1PSJrSH3a0q6RSAC4q60pWzSLIfLz6LQQgLjJdvgQYzq7b798CJnoHo8bqPgpL2bqUhrYTfP5a
Nk10lyhUDoE9aoddMFX3gt8Nvbx8Q8wfuiG2DdB6vKJhG1PcNEtJhiTiEXiq7ySFIDEvk8kR9qZe
6XNxoLUze7SIEFl8YqrsVQ7aKh6nELDep7gYT7ma2RhiaWBVtR/fP53IMyLk+Ee4zxWlHiSoJyb/
x8GTuqMdqKNK64v0VdlK1kWHsERVe2JL6SJn5AeSCb4kV0tFetnrB+DxKCkOsu48SpSDVeqo6Rdp
5llHPwd9Pjs/KWVVGl2zaFLaw3bp9jkMAhbevps532nKguV4Xp8XbFgRWA5tiKXj1pY7YRh7CDZ3
deMQYiB/7FgK3N9BxgvxYW97qzYyWi1O+TsofZOjQbPTNsctM1jT1o4qTHYT4NuDxIXCZhepT+xa
/8JR1ADaUyFItdwo5jpJt+aDif2ZHGPzGUVky1KOVcTH2JKqsrOdw3x97nSnYCexqekNrDdEakDE
XZmnjN6uXwFo9XtHy+dFyr2fZNTCyg248izOe6FzgfgY+RI4DBZxosu6YOO59KBVOROCG6mYfdCO
KwMEX7bmYr+1sXY0HmMbkqruruFE6HalwvdGJHAppU1u8bf3qP65LOWNyro8GYD0rkmaPXkpRz9W
FXw7RAFiAKbFOFfOn/ucMQHl7PfNlwK2/LDMIffbvMvUYYd5e3hIoXxBLcHL95PxwW9jLd6a2MyM
KMPlNSHyKa9+d1tOfoL8sW/TA6a442Y92RYEZTgdsAJi/UKm5M4NcqVKFaVxxsLFbAMLHlRhGB8s
mN72bQ5kWT28wId0gILXAAwDjrndfVI89Z6CxkkTBDDUpXAB/tmmjBYg8YZQcCi1t4j2BRXSEyHc
ftNyVnSZ9734jbuLQBGWfglvfYyukvE2kBHZkJBqANLPIuWCGUccmz7ubERNXy9Hli0Hu/KT9ANh
LVxtYb4grwkWrebTtMe+0DJgGKzoJ1gydB1MLOGejRTFTbO+xnYW8tuS+58y2AgVDuWwYdE+N6rY
Y0at1HRI2k7gbm48G0Wp+oj2TP/vljhJVQDILncppZc53wmH4DvhsudoNoA7lwJrJd7RZEJaLEOJ
ICWSv1NaUtgBSkAeexfO37cHCe+hPGo4a+AZT3RMLin1+WfoV+UEpWNUGAN9VQgedNcLh67YVtH5
BE/cjC+ts0BEDaREhBw6KbjYKPb9eYjOPyDyUeYv34k896dFkj+vqfLv9vUtXouW4XvygX/gxH7N
RAT3ID2kQ4zs3gKOY6kcRQXql/nGsjKA918QJKXaDxH6YnyYGV7cYK3sC9ukZLmEA86SVuWiZ592
GI+NdC0itDmvrQBJYF4R0RgJpSSf+wYBE12XzttQLweH9Y2x4UjgXdyBUNeSfKMOk4lEF+uQ3bfq
geDvWVFPYwK1Abe1TEgt9zz4v9t5k35e5G0akLmzVKKuiKqx894SNdJkDxNQAoTeo3E6mYI/AyxL
RWt2GCZI9WWgAVnnuxToj7Q7kPLZu+pVUF2NYX10S36NCe9trWcBfGQA9WpbOzKrxRtrz3vJ68oH
RM7/es4ibBC3OGZKlrYthnAL3piFEQlrOOI5IDm9HmHW1a9eyBbskNiUHjZs0EIttfXZGI8DPAT5
80+nQ2QezQeXcvFeD8iRfurrcyUSw1U9C5RY5wMy348Hh6OGwz8u8lcptlBQ0gQRUsp4yeqmdIi9
51DN5i13Zdjc+Ksrk4aCEVj+kqnKaSQvq+KHbBhntnwzlTPLT2VqiBc3+TwGNVciD9Rkr8iUIvDX
o7m28FHwgvbespPn0nCqtGMfcjvmSj4uhNHalIGaqCZcAyt7GsvmsRbO4l9eDw4xJnSvfw9mapfi
ew4T1Xcomn7cCJTLfkzZKF/iB1B+jFg5Kl0yv/MWnGl/pAuh1eevL7/2TD00b1l/9lz3MyUNBaEw
toJZb1L9QfCY6Jqc+zo8b7fVXMLaW17NOvjbDuW9J6r6QY67WKDM9XHhcwETdmHd7xJd8JQqJRgT
mglKHUZkybzjQzewELSu6BV9cDVvR3wMB6aE83GOj+tYVS3bN9tyCX4plysOklq17IiXNiIEoGkB
Z7Gh5GJuClBGv0MQzuJKq7+ZssJPWDbH/YV/DKum03U64Rmmra32fMM9yW/dQzBeJnMbgwF1fzrP
4tVx3r3ueZlXdOhVHwtR7Os+6spcpGAXKADWWhIOaZAN8BvVxtdICjS8YmyHFhthaU3MOQoXU8bP
XZqBAWc0Sj1HcOsl+lITsVoOkQVy9wzKYVZw4DNEGrVxF2NxgDVCFLCh6m0ySAq2RsE8HsTssegK
fD83U60R1w5i+F9DRBmUQRqbrZ7J/Nqj3uZv/kCBWSh5RQxWBHZqJ4Au5W6jy2B+eRPPhvNEgxeP
P82Z41AqsNhnwVZvrP3qBdtud/p5LHY2aKb2O1yT6V99uxvHfLuX29dPK3hZdPlvP236Ahrxl+PG
NLGESu6CroAsNjfXEO7FVwv0GJBQ9VvIdqIVVpQ88rSLC57n29yewHHhkKc2v73pKHObUbXc4TRD
AigL6jvjsN1qJ4TUHAhu9cfr3pOLITqadKs//3VjdMRMXHZJDN/2496s74lX9Woqx+qU2FtVsddf
W8H6+rIDmYgGwkhYVmGKPG691hARhcolTj+Q9/fc6OzURvwdTATtzpQPCWKFc6ND5VotQOg/nX7l
L07ydVbxl5zoWhCuY2YL0Cpcd6iAtrH4r5WwaI6UofyJXEuqCeSyN1B8f8wY3MEaDqhal2WkkgdT
0JKVVrpXOrVcgjj4OLpmU8deDMw3s+3ClRpO5N+OYGKAgBiuEqlge0mfk16RrlUvU0IdX20EXnjl
+88XTTIrKXIEwweiBd1x0ic0tcgDZXSmxkmdA70+QXg0MXSW6v8IBUjfOBvJESnc1XgxHPCFuI1+
i3yJqep+zNtTyKJS3lp44z02Vdqt5MrvIrtKuoGVwlvRtPtRGnmSLk78Xsx09YdXn6geObzU1bN6
p/QzT/S3fvZLUrMyL3BBqWw1hJg5rsXNOvJbSaruOuQhyw5pEIX/jXcaQhJOSctLCCtKPt6Njr6X
Nml0yzICOG3PFQVjc2GBWOKOXvV7igTySnGzjLReGd41mh6vcRId2nryOEQuWxBHvNZYcawLKl5P
fcRyy9/FLaWYvYyPI6uCAUg875wr4xM5gGtVuda9jaiYWvPQ0kaXGH/aRSgKLvPR0gQCnLHAVhw/
0R7nnxcc32EkHIWzSErcZww9/TdVFB6RUu1bdTDoc7YO7XDhZR6dLi7gpZE5x8ZePjJ2OMXrytq3
dqX2dHSkkEWoZWs9KRfIjWaIjD8K8cGJcmsEJEKXJFrTI6o1t55I8ZQxeWw3RgqGC4T6h/ED80xl
3MZO/gnux5lQktenDoXsTeekjC1hMjNfBSNSTLPHnJ2E1NpJpGRwPihcT9Sx9poXgUbCP58jMoQ5
N9i3jE8hZ7PUGgKck32s6WTc99d4yX07YjqGlnAD8eAgF2WGqVxtlN29ts+F6aRlzY8cjzMXFz8k
cXbIPb0nvirOgEbNFNFcs6CLPjOBVbs2/N/nYAVcLeUcqliXp8IZcubaXDvEi9JwYVy0K8jwH/Op
Aqp+CBOB9R9zdRQ349e8Lx9ud4frqeoxMNthck7YXNLlGMShKq0VfcCwl5Srjb7uGHsZa3/s9Iw8
Q7msw6jv9g5ZGVZusaUjjY66VumTl/UR0oddqiefLQJWnoynOgucOhax+oRbNPcNKoCdiP53+3jH
cyGeP0O5E2cZ0QlNeF9Kg3Wg8DHtSuOJjEO57hUvYHfI7930PWIpQ5Gv3wrHKShtNFiOuPnOCKqk
g1b7B8Tkxfoim5c9IJEwGvA2dIMCktGD4Qyhtl6Lq4OUkourIQ6OrASr5/TEOu4xNHKYKLxh+Cli
B/e4MTnyXVOCYPGERTr507/16O67RjgS0y24i5Ww5GhwsxYDKYA4v072J6YT8Xv5ZaM05C69mAt2
qAWv8gi9GXmoDNukt99eiuHse/TXF+kctqHDK82qL5hq2ISKiCqJQNvY4zYQr3ILTKY2JKCLqW1v
Nq2DhhMUCIR2tTX51yDEKGNXo2iQZ4X5pS3V/ApZzPbac4IoPw43UNLNd3UkWqP0Yo++K3h76oAa
p94GJSPYdxrENk3R2zNizX3p21FGqtUmn0hrYkk1OuiFRA+eCc9XWP7vMlzHyJdo0e9EfUHFdB60
inVqb5X+pI2uuQL7tHmFDcI4H5Ro1SXwhCj7LyfPvVXnFUbiMMHqbDQBySbxEg9z8LAr6/K6fcjb
h5FG+TCSNv5q80Qn5FTRzCgYHhSenC3HvAEoYlxayQf+p0ksV+wsj5mN8t6skr/4OwFoYSNGaSOY
S3cM7pdLdlal6x/NIQfEBIO03t7/35WAovs5jPkPDtbfwCeuvqWmE6JAjXo0qiVjsekv8LgMmaP+
tYVs+zebPLrbCPbdYFItNdt8rbLqVdnWjYuuk8qRVv7gSYq8jECT1X9/0tQhRP1vdxICHekdkfO9
7r8sU+bKgqML8JzGgXNjLpRx4e2VCTUKx5ei0oTd2+28aFq15KFqdvCfNj1tbO/K7G+Bh/65yKqR
C5hk+UdjbjLMrEQ+tRAiztBy9bZNTX17I11W34LTif3aEiL1KK+p5lSwOsFsdiev5/+T6uOkuF6G
xhpvRUpgSvsJ961OpL8sTKYtJFKyh9E/WSUV/4xcrQA0UAnKoD/e+vlxHrxySix0lYIEjW0lzKth
Ju0vVWeCsQkb3DdxIixkRcIoVG800pJ3djcA75x/B7e+BbNY3FIErdUiJO0Ys20ae215e3bq5r7L
FvDsLWy8H1YN4dhpUqyEAPFyphBQQ82amT+FTasZpRUikd8L7MFp6XU5Qh56fI5Rj65z4rrPVKVp
znbExTk+FD9N4GmK6S4tPNiIwhrVVpLG30ZE96tAaemZ0lNImRRj7AFmBrpPRmKWpUU+WRvT11EO
Rg6jbyIoJCse7unG/sz5ym0NsBcqg6G3EI/q+nUdVZjpc5wMhG0KX/jYNQMVPsWRV94z2K63PHZw
h/F5ME9ADq7DEToDyhQG33ynvw9JcgdyyzeQnvWnMYWbJsLMLBkCWZDNCwLdqJ7Q8RsswNFIEae4
cYUTDJ2ub26EV1QM+8jnmMefAb3RAnZz07OZuLuJXjZVs61J66WDY9HdMg6xyCdUNLNiIRLmcArX
kXrZiEmX2ztK2tX4FzLlvh9G/ySLaEdavCoOsElLdWEpcUa4JgEiQnUH6qzI0Gy9I5mxpHNB9HhS
++ruyIlM9Z3oiAbYxek42hVO7Pq6hUydVWAxspwQHcJFbnDWdXE3X+zi3rAfWf2DLeBzCBiooRts
653jiPqCYIO1xgI9H5p+0Kcif/qTHUvGryydDmpdmEB01IvdgL7ZPvOt+0oMzSIZRNeeGt5Tsi+9
ZwNnq+2zym+NmvaFRGkNb+J3YOI2cNnWyHdFEE54ygZebCbZ26VahASV+042VLICbJ4bZ3ukSbg9
QH8D23CUqD7qkG4G+0FEngqPpxSkGxIaoah22pnEgXcel3lRS4iv/jEb7tcyE7RB5LBJcyX7tgI9
++qtphNDZt6QpIt+7fwJSLSQVcvSw5qm4HBwM6VLTr24WZpC5zEFCuxlgE2cI4AZtaYnSKerlf6R
jT8ep+3X2pA9p32I5+oykho6pfNzTZNkERICtkQcMbix0lQ26WgQ08wyjbvWw+BCJWtauEVSS9lB
dfHjjI26ij567MELHaKzdD3oSM8sdrehX3OcJkOQeloX+Osxh6m6bujDoDdgcGmE5IBtrrCdJOG+
Bubh02vOdCug8UnHT9fZjnRTemoVZq0b35uAtqguJ7ObAUgGvW6t/RKp5iZvLRy0Qe57+g6pMBRo
QpCsi35SMP/afrLtfTIob5mKEn+0FB+WB6nRqDmDGgvnNPF2i8Ee8BMLaV8uuogS2JZc5BZ9jxXF
jxJZnn4R5RCnHSPcOMJcZvcj/dNveCLNUpCoIYRJV7PkdymVFFYb8oMVUXTiDEWoh3a8Z58Wqb0K
DHVcqJ0+FsQG2aYBSEwEH/RXIXucS8kl1zfS8zTCxg96R/wfEJvPlS0InpSAFj7+cwvPcQYCKJ36
CwZfxCWpzxQqrO9VY1mdqc7ujlnd6LLgrf+tZvzRVKyeg0mFAu/yoz7LFhAzZZoEKEh9YsJK5UJ/
sJOamkVrXvwGCX+nr2ulSLGWXvsVXACOS2+NX0n/cRQLirNBCxHElbKql6GBEPuJqgatSO7LcU8P
9yHW/E89cRRMqByAXoo1x4flQWV+WYkDDYxZJk2AvN2nB8nZQhJlkLx989+YB0t1uO61rPVt94N6
onV7/YdsXgE7JSOlLalLvl9pQq+iVAgChckjPd2RbbxoGtgs38UsBSUv1MOB6n1+Tlfsd9ymWcWx
qmA7PgoTjearISPW8MSvbIbeD+34LvfcMVVH8Yj5U4sSohGILUPd3MFzjweHGJoUR+hZ+Fdg/9AJ
3Bx+29LWoMhsWu0Yc3OQ5N5m8CIMSTfmFxwCv5ChIyf3A/h+SXh5sWNgbP4uRR0hndrZsgZyt0QC
s/LSK0dliKiSKngSLjktjIDhH2NMMF3OqM2FubqJ6dARU7OOVtg85H2VBMvJGcMABEATipqEFNs/
Q3qtIuwLgygVXgbK3bUxokqpPOInrKdElFBFr3vFAYbG/qN5oZHxKj8bC5cYcIl/CiYCX0OkMjRa
RbNjKnwm9HqN3/GHC4ETowya4foaTpBVfEGGcYCxoCRlzMhDgvVZv6sr4mccxvUhCcMSa5ruLXfn
nvp0XSmx65WeAvgCUho5qa5YC6RdyV2nRf7Eyx0Ug7ItC7pYlKXbJY2ssbp+x1BJuU49TuhoBkOj
/L0PCiJdUnwWmWXiz3OWuNypTG2ZBf3x4avQ119E20OkDEptmxT/MqQNk0lV1OXma8KSrPleRSzu
fsDZ6RLku8ATyjJ57HkSy2Grv6yfk1NLoQ7UbQWuQfYuKKWrmpETVYN0edufzQ+P4omP9HAFMBHA
fhJSP/Uu5efR1RBWWC4RFY20ko/cUN63f4V5ekj5cJH290vk796Wh9+X4Qdw1pFiuiP0O7gv4Zjh
e862CEzt/3FIRdgSolcYMlBGDysZDDcRAAzGAMTyJBUWQddUjD/FlHFjU2olMZxOeFxmaHNpWibI
qsdS8LgNBQdOZFABANpTizsrLlnyOx6JfkrmVkNGz13HPmwZYUETc/ANJyv96h7XAVadvvu9MVJS
IdXmY6rna3CXNKiJiSrbjiz59TvJxXhqIskG589jyi84AU6Hj5Gi+ptz+XwGwyyhsSaD/mtt031T
DYpDPNpVI1/5gpXFfDHMgvA1VWuqzlTi7hPJnLwQROjzfdBrzneUcvIM9k77ipfkRmw52jBDEGWX
PpBEYyoYK/gFs9OCLW3lHo/Ya41ivY+w9bBYlO8u+RJ0MRVTX3TXIOvHMRsSF82RsMHm6lHY3UlI
TmEb1zvO5McN+MligivJBJ8hLpvOmD+rU6nSU3zKg6llvcLXgEnLmbQIbTj9DR08r1l0ljnTPsFV
b6V27qKq1yBqqG6rQ+fQm2MHjg4rTiMPGT00K3iD/+Fi/M01GOAa7qIbChjGwCDfUN2NEQI/KIoZ
kDOdSJrdyBmIVsTaG3wwZ12qB1oMgIVwk1JkkOGQDQLmizT1g0Axsn4Mh8EMRGV2cBgVkSb8SYI2
WoTJdmvQzUMtQOw1tL63McJnr/t54paxtp1Y54f8CzQCvwpV+eP/gmpm7p9/uZKQtG94Cwvuest2
DEG9EtvVZty9qF6FqLFL70FB2WzknlMJa7hrJ92aRwRtlP+bqjxrkhX4E7A4KODCHFWl1lgT08Zx
r2PeL4JkIuB9BKeJaBhI4nDHaaZCZKL2m/lj6noA4SSbzT3XN92czfY8LQmb2tl82SlmcHkOEkkw
A0ZCHYeLETsgr/UgyR4fvvbXN7LFnl2KE+J/1TnrUhHumqJVRpMC1opmHWBraxum7IVf/CrELGc9
KzZcFnf4tOKMfbT9vQ4VLYafGrEUlIRAb0TlrnxVAnmEpRpkfsyooT9oKDY+zbtRczFHtHkrPgLA
Bg1Qlyi3SOSK4UNuKgFao4a9nBIuBwp9Yae0Hv4g3Q2SK0q2Z17EW9rs+sZDCK67oYhQIYNXq/li
ek/qFQC07mljSlRKY35g4/IY1hSFJb5f3KVMFAaZ4g4qbqGLPyj14YYA6WtI3kpON8jaU4HRZvMz
JB+VuYPZdiBTexWDsXHo3jUrYXc/ntypN+CmtyCDR1yAbz6lqmO9jw/CzUZ0cA/Fhu8ApoqywAg5
IVxyduJE7zn41z6wjUwCF5Gjv9WgdiQF6Z73CsHMwje3B/eBJS4TFXQsPpDdRtXJHw7RIwpXMNv6
JYKjVsH47nJPZyDZ5edlQsmLy1Dy/YjpR4sFZ20TQchOYPdFotbpgfNgZ2z1R+k0rXMSgXubo1Ty
Kf3QBrmkSkngxrghp3I5moYo6TRYsP85JFO5GNk+dIZf4qq7B9yR7nU4vFjEp6qq7s4Sg+o6gHSI
fBuYkLOlfhB5uRTmrnVAxCZkBILlWl4B/R0+IoyL09mghrMKZBPgLwGtxcDxo2KQg4z1PSB0ox3E
eVmFt9EGwHrZKV3EQCYNMLNgbc4CxQuPsgnSCZlCLPABdLZURuwpU2KNygdn9ojGeM1TCf/X9CVn
gWJg7NNkKWz4c8Ec/X11tZO3f9JMzbfpxV8AOlKGJWXJ3cGbR++HpGkBvId1Gck1W9SEI/qLLje9
dV818cwHCd+9z0Z3ynXXGf7Z+NaVIk8JFOK8sXG1sJRgZkZNYAAWGL6uHntqYu6KaX+gEffXSPHh
tlug0LDQtcYm1R0SCXtxnqDHDUtS1qQEvtpSL5w9hrc2UElf73Y7TWoqgNnHE2dgVYtLuFfEh5ZD
7oguutRrVnIR8b4xzYsaoPVzBeLQ13gdxq4g+MTjF1s4K+X+NCNiLPBucCDnAkbgZR6Ruim8UXji
wg71AS6wPBtZSa8yN4yBXgMJzeZ/43Zjk8/NIlUYbOBZCeZUml8+AD2DQV8zsZu9N/XGOlFdg4Ay
ndA8k0Naznu1cCOIHlG31dmaLfd69FiFhAijVPjhRIahuB92FT3SO0/n0UkoqRXHVaQRyTk/yQbi
VA+ANp+VxKmSFlKxXYxUaLF/ewfX6hMtByPi8ge01D9RmttTAaMrFIRqzNZWoO9TgfEhUI/XrCPm
RCKsyIONzeAmqQYT4qAHbF3Mz/of555bhab0tbD1EFI9RqWX+vxeIBtIOnFdTruzGv8whMzYHQv5
J5QqqFa7IFfsFouKTvMQpSfchoRlCdWP/dm6+i+2c44pIoS+fEx3XNp3H+lccY776Zbt7+G/oiK8
p9LA04zUvTRKenafczt8PUnOfd7KZtbygEMxrOrvEubIXWXTW62L0jpOFfcw75bCvdQlNOOGHhuX
xxLj+GywupYbeye/ED5tW37Qhy5Cqn1f2ODObc9UQJ7fhCKGvZN8f3Ng2gDj7m+q543k/NYD7zfV
6goLvNwttjS1Ijju8lFsBQgbeWx7VrpVEfWf9LhNLQyuBEYYqyAhIYNf9gLNEttepQ5nfV4iKnm+
XC8ttBm258yk4aXKmNLFVbfTCHnYFjGXjtDWEURbPvZAnO6L4Xm7dX19REUaob+8GtTU56gUEMpV
OtpVZjkZf6EgMt8ZglP/JnrHQ861mayclzfRnzdJTEio4D2DiR93hzmHe5iQryIBYAveJHMtcfUn
LVdOe+Xs+uUKqJf9zq4VIbVssGCHLJcSGHVI8sye2bViHlWOb56I3JGX7e5bN2tAL80EUkh3Xmk8
AcGHDqpYh1+2maOhTWenqsUlttT1xXgX+T+HGx3DSYsK3v3TtZEiHif5Xx7KxcI6Sr2qFdPxuzTk
V2sY3T61aeX3xxe7m98bC0A8kSYxbKblnsWRnhco2e5TqHrRcO3W+VPw0EpwYxTwnunfzl5A3T11
WuUjxtEBvXN7tkbJUB9n2KaseJHkVs0+7bTRqO25Cs52YlE3PMSfBuigG9VWiqXDXnCBsNtm0ONR
PGO9FnEoPddi7W4m6K+C915psYVM7VdQmrpQlbo2r0ZeRH0zX2aP7Xv8cEoqozNtzfF3gpCwEj5b
90HPfhOWHT+jRsJRvaVivppJGEN7P3Wor2ihijhXxmjc032qa3nojwJMnKtB2kgDsAw3mH2h7LsN
VAVXA6JLlBa2WxqM8nH4AMGaK5NdnZPpkYfKSqHDnCJBhQz9AGAKsI7ZvdPoXZcB+av1TL5zhM3s
guPamQkPltxZOo0o15iiBKqSeR8C1IV1G0mxAxwiqnu45eUnvukdpmG54kpgsmZkhcne4/He+l3b
mCKwVHhzdupsTL93FX9jXhwvFFRZCwKNgXwQmjNETG1ZwXoDVZQi/IIb4d1b+l2BD4MLa9Turtzq
21VGa6OgDzIl8jEQjiz7vE98s+4+3CcrjBL8Vt40DZby29UF+pcLgXvs5n/QmAsAjywK5ic5xjbr
Ja6FTrujDMMdM77pOsY9EYXl0iJBBH4WjXUDIu9m5BgzFM8JCgP2Wy+xtWi4tnkKI0y3mQjjXO4P
4itvDJ99MmhCkCDWHnq/gAFC3QPNJgJgR2D1ymQ3IvVW4NpNxjQxuPMGP2UIE3CPc+HVqtOXmUWf
6A+xXSwVZ4mtw6Ql/+bYjWCfRfJo4QvDGm0ka77HiSHFYHtmPYTjyvconr4yC4Rad/rkreiyakEB
IxeAYu8GuiR134aufystMconnddea0YhsRgLCjCB2phdrEO6Q4SOKM3ep2eIUTnDtVanvXxbHNFe
LWchUK5IRVODdrzqqSxvtXDFL+31JYTy7lnaMVSDA/ro9vwjYCO8V4ip7LSWkIj5kHtT2u5mp4cB
KMwAyxom5t4/AMJssqMky9IEmEeg+s920Xej99iD32+tN++hQrY9i7CktlFiQNIO3vDEf5vVmATr
YOeXf6ye4Qcqw3Dot2wtr6tjcl2vKMiQvYHlVjxVeJ0Z/iZhqQ2oBdlrgOTMdxlSJdm0pARDQ5sE
w0UT5pm/lUqS12KQC0H77LzWU82aBdV8Eh+O7CBbIUV5wFi68C87X8Ze/GYj3T8T68XCrdQWNs7u
yTQsz1h2yMmfN/UvqrFgbTYdySE1iYdYmrokGRiLBR4s5h7mMgJTGPgtidT3gFEm1QvmSGFEdxNT
zklDX8X4cyEdzsAgQFG1Y1RqgEwEDRDGzjoz792iRpFgx0O5SXOe3+ceNCrcjUhnLu4NY/AJbeJq
jbbyvN1bPfwjx7D5QhX3k0yrQgECOXX/w5TWmHFH+x4wvDh9Xwoo0U+gofoLL/XO201HLcw4El6M
eJWJDpEwVW0ODroJv5qpD9hkvSgY9hWwSbO3nDdlouP2ku/Cu35rCNRH1sBuJ+SzdHbThk64g/Ew
pLdKqwV1gRP89kBw5/m/ZBjjYHM3a6D1q20dIb12LBbTBwrdBtKGs297LXVeQUGLscHcHuRzYcWA
Ey/3CSVAMzgcy5ZygZOxPVVQCyo2G1ape3SjK9Ib5AFxO/HxFBYiFHAgdzO+9z4jd3QgiIpVFmAn
7l6lXE4/WF1FEtq89Jmd619KeSUr2OWW8rtnJzuAAblU1XtQ65hk4QzASk3jHx3Gw81BYvdcgSbJ
Y24LXoona6a+KsY9rJVKYBQqPAUb0SE7oEoXRAmB+Iqt/0ET3IfvxEAv5n5Q6dgo13kX8gpcXSPd
845VMPdTyVMsMBpQjZ8bWjqMoL2vlFv2t6FFPIxAzEtuPrUY09nve0KEV7R1Stc4+OkQoap5q9NO
C50GeeSWa763xA6ZuTWIo6x+ILgxiUe2Ln+utSO4nNb18ogjUccVGaloMOOGuztQGDPkDvpW6CjU
HXMSlLJmjva8V66n/QjEuFY3PBQIKndFeXKCHD2GM5y4Nuq89VqjTYIOJ5+kA+8AP+SkEPM2CIhB
HeTMKD9t65dt+N1LIQUjDFZi6N/175aqnfAjpK7Qos/9PbbgqBBfZafN3qaQ/K/xbG4DlpSpAdfM
JbU/B+C+aYO1QpZ9j0R8yU6XLOgjOBYKQvRoB7oQufLQcng9PbLO9zWPZv+MvOPfDzrZdwCF51Nf
7KRzN8NmRCs3tQqnnBzz1WbtWTL5zvpaj6WV1hwbrDSshkk1cZr5Lj4G+tkTaNMeIZ2S/nPAgrRU
J0Ymcy3jRcmOiY6Q5escJOUwEMmJdQZ8N6dKNtuJtAmq4PdJOjW+YLrudMg3llG+3DzIePkp+zcn
XnM+If0i/y61Ixrb74yD7cN8HQsMiCCHN/Il9OVEejyWyl5RaJTg1YZZKxq9I4YLm73sV81rxtRS
2D+hLcW0N1wmWqAtJHFl5Ldrgck5sMMSVDeig057TYXWtLnn+bo8/jMdud83njkmTWZvPPt4VUtC
cjf+uPMg1aYpHE4b5w2GzrI+aOZ9Q1eOYUq8sOK7FQdzMw5V6YQrK0Pv9hGVfSQAjY8AP9kGnvz9
XK/McFIO7QeMik0XXaxz9d2fhQPNLUKUqI/616koORPCH2BLmuOvCRMI0eSgjOzOchM7QPmKd06l
aP38vi+6AIas22MxkJgQJRhYF3tW/89LzZROvsNLDMWXnXw/h3tQvMM/+SH+MP29I9TseAnYgRbU
DqVC1JpJsB5SDW0IIh44zAu+aK9bwXL1Rex44oPKuj59SVsf6wwF62BZ37n88XHktgx6q6Ki+VrB
Ss+W1Spn0NbwwVjyK+6+LA6hXS/AbfWKdf6E6rsAEGiVmBZCznJQDH/HN/DAoyHetncuaCmOEZ9C
Qym1FNGIpkCCgmmtP/6X0gPczzRqJH+8woMHMUXcGGmyZmG5fjXTQx1/SEtD8cjiGT/g8cSxvgcn
DmXA3MsUhMIqLOWWpFofTeYLQnqtMv8UcO0OteUWkZREtBMrH5fQrOTZYvAdpn5pIdoEEzzVTN5i
MK8ltvT51DHjDV3lm9Qk6mCr5ksADVP3NEyZL8yKKvCE7Sf64CImKgA4AARwByPjB7C6uizKnWEP
f37sHXR+QYYs8Qpwm8mB/Jb+isr2wYBhVBxTMc3kOmk19W9EV+kNRM5ZQjKd2ILObr3aH3rqVj+l
HqkTf9I7mk5uxK/Ld/NChb92mP7wcyLqE9ER6Ev9oF2UYsHOoPvv2O4cDJd56YEPmBKSCaj4QaOj
23zfU5d+czOrSWrBOO9zHJOpkcyLkV36vnWT7RzaVgFjf16Qr85TmyUryqbsfYItSGSaE5vZSfX7
VGVu3//4Z4e4m0mKsOoa4s0bgHMjb9bdd6FCrs/DNSS3UU3fqWKW62mNdnNCO3kWW1r8uHqDaf6n
427WY/eZvbQpJGzZmvbruvnHGj0HHH090niD0d0GQkW3zRiOZcByB7x/I4EEPxMhoqLpDAxxid61
RH/bIBC7kGhRA2OXq1gexhhf6F/uXvP/+PuWE3DQl9AYJ1Jysno1W/hB14kLDZ2gYFJa3KgEfa1Y
OJE2l4CXpHcCMtxt0VvDY17AAOyUC0dO8L8V5NamoYGSV+CWKMedHcpEJpyUDpWswO2vqWz9lusB
KJUleLe1C6Ub34H78aN4BnUeKafyMUNtK/BGc8D5AVgmS/fRG1v9CTf0YRbwvmd/igaUCYZf5Ruq
F/Pp6UUt/TxWlZXoIJh31NQ5DsuUhO+SakKh32dvJCGDQbAaKyvjI2iODJHVOk4bBD77cvxjyFRN
m7urGUbX64w8aYxbFk+ZC/7sTp3rgURapas4b4eZAro2fwfVNBa7l31WXlWnH06xzv21I/Pztycw
IBlqUO6NIFhc2rzbujDM1/BxowdX8Etoi6+3GLV7xKWxuUJa20KpbuqzXST92B24Q1H8lzdK8Co/
8s56xYK0+jTSkTQDVCxiqyla6p4vrt5tfefnMPAS9SUfyuhgzUBPwE7ULCNsLBene14CWCD6UnKF
9AbMYPECp81/iLfMpaOiakIeVAsOnD6Wh+dOHo+5neuaJdBJkpuxzwY/i+MYTpT0CPOlS88UxbUq
FWk4tXfAJyuISREcl+7iAPPJNzITP36wVipvC6jWlGZAU9qNXeVCkRk8DVTfROPRswDhqGqQj7th
+DvaGIKASefQ9j5d69rjGUQXZviJ1JngP8BZe7jqJuhhc4LHEcAnCWsPlZPrstsY5KV9cNG13K0T
5inO5NqUk5ja1GUYpk0qKchAArcqyrhD+4b8CNShTsomOuLHzCWSSBxYm9B1F0ud7qFOFKpGNLBL
ljwFOiakLbkFGtkEj+KPdx5QtgZPUduyeUISSsNlPJh/Gl7aJ5UuVY9UBO/YFShAZlsEl2HxWpv9
vC7uTQ/OSeAgJWpcku7WVqf4Irn5oH8tNNTRMAtAc8/iG2EyOmQ1gAlM6/8SbB7yd6IdyJR6KkTN
k86guPaaS88/UCCGqyDvp++PHaxwTfzJMldb3h0w8IFWnIHLa+GqYjpbnJ11/8HtUsA174b3YK9I
FvP+AfURWrwFTR7g4g3inSkC3getG8zFy+lR5hNteu7wlAvUAsW2JKbUCfMkYZgjqY4rEZLHeytu
RwJd914I4WwAnoo9ZVz8LxfXcsWagdCR2YIzYwyjSEJ2AmYzTek9wXnJ3fmX28uIw4IpTKC/iKta
uWIHl3P/2THe1YpMfYHCgLW3ufUF9pp0YBFmg/JQu4t4cJNC88fKgIgbvhlVe7g/xuSZ+IGOK6h2
VfT0z35a/Gmlkx9yEXwS786u//K3W168/YarK2/NPE4mfD4pGhtHYW3chg2vTHaw1d38WJuJbFHY
OJfAdgQ3HEPCjoOOXz5tJp5nSAQbuI1C6wxn3dyuD4UO9y0wpucA66XFzKPm9QDvy6Pb5agpZ61m
Pjn5enNX2Bqr9wqJvOQNkxKIxE1XaY//CGcyGQck8q7UZDoURbUwj068Zs9ULqoOPjnRBF9ubDIq
Em21FuPAAETJ9flweukzqXRrqQ2fKW5FZvi3VPQZSKEdzYhXF1EDXPXmtjuBdIcHaax1L50XYK1+
k3UgpxEbbNMEn6Edl6Y8IS1cfKo5zZ6mZazVJcvxAGcNJ0Qv6rbSbZjyz0DHHTZ7T/lFRDdLx3wv
OFge3IsBNDnWgACk1Q+2PZ7EoXRANNH+72Dm3v66wNk+jJ5RuqNKE4BhWp+9VFEMhoGpuSjlV5dI
c+OI4gEwFQWLS0yysQQrbss7vpMgH8NrpPMuVaWWNlOw5XFDtG7jkzrN+OYQtDUYBiBNj4Hb4vVT
zk40M70SUZjxj9pHAUJ6cnIRZngGCoJ65ku7U0OGdh6iXn40aU2v7hwcdO3YxmjPYTR3wUQ/4QV1
jHjKfo42AdOvV8RZKCdLJJu/lZw/sPQGxFQoNmG56cTXYqK8yXhao99ztk0Gc7Vp9BHQCJzh/uTX
krAcQ3Uc6QZvVmxTtzhOjPJ0HcGQ9m1Ba+N0yI5PMS0dnR5ZIU8dlditFD6/XajdYShVx3EN/wcJ
SAymiPGN9Mdwghd0cozumxm9Z+UAxpULo6oONMtEah8EsZyRsOWT79nez/0a4o5FVbBSU4i7YOD2
s/4ns1iuiLFHWmcWb+Qqpp3UgwgLrmA6XLPr8ZxFikC4Smb6uePV6skHOTnM86+gflx6QJw8j0fD
hAfPcgwYkl7rVGinsEwNwqXNAKnoIsllkmXI9eb+gssx5AIdKYxvUJVwR0N87jB/llPjGN1YeOSc
6jvuXu4kjwqwJ2lEzjcWET5UhkMX0w7Hzn5eFanQexuXnuz8T9T7s2xKGA4QqZpvcG3xX3cGUWT9
4XGVGvW4VKd8OteAorZfo5I+v/WUuIKG6NOTxmFbw0kGEaVU1BAe/O74jD8GFq8CZwNPqwmW9PBP
eIgVgiSB/YF2NjJgWmaO7WfXKlj5xjnmf7vK8t4HuAy8f6REBZrpRI+v3RGnte7e8ZLx4Y1L1ADp
TYJ0xz+uwPlYuuQRiqKcdNIzLSpR0rN7RixZOoFSu4bwULHu36yPV9surEo9b9jcLojfw6XekO63
DPoTHzkpU4l6TiQBLPPL4NJIpa1aNk9VtUVRKlu8ytmYDCF02GVF+qq3ErIpMPt8+4Q1nEplrz7U
qFJFaEJ32jtYY1lr407U+4Om/YEbj4NWxnYjSdirDOdG0kkvunPbPgpYCseOzPzqnMXJjN7g5ENY
rxymOL3u9KwBrqzZApXv1tjPXubr7x1dL2B506WO13ePgtiBOsvqxL4LHTnqaZuILZapA4l7UBDu
pGAnFLpkKHnseiB+VgAc9tL//+5j8R8OJcgjSDRZ9Qhip3uXXHX2wPGv0MK/pB88vWb3ptYOSqGR
fcrSMnk5AfiufC+vXmawXOE3VbLztiDkvQpHVsuogwixfxqCoYtFbPJp2UUmvcWNAu2JJ7T6B6oa
YujN+XTRm769g8PnV/Jhm9Ve9B5ZZ+kGenBJMl+0OtKg6Nh5f2f3+5xyhkWdgphivnnHpGUnu+dI
+194OCBvrbDPj71yJhLFM8IdMmoVHoXEoREGp10wFycnzON8C4CozBOv2N7k1rMfHea0KOF/eKBc
H4YVZS9MmoRjTL+vlpJLpKYa1WvcL6lQwWaY90SxbVHV73VvTwsY2P6Q6yvLIUcFjwMvyoKFuXy7
3HpcFV9iNQeaPwJ7K2rAlB9jeQHsOzOown3DvgdsP9BFAHNqT9sep5iJgz8aOkAnnzKl0B1AdMFN
BBhJvH9KzmCe0c5lNzg24o5PLBdFPu05Qp8kVejnMHNtXBY+0t1d9mrppU2oEk4QrltG/TieqXAg
7Uu7cFyLI/h4ZKtrKF3N+GXWPE2EW/t/WPbfnRepCxJvaGdg6UG6nGIYO+gTb/wH6kWFTSp87IUa
18wYMeXErjt/yO41TgxXkB1JOkFzki5Y0ETn0ZzeVmYgp5YYO2dCLi4MYc3A9XWqYlQrBbOfGGQH
AGWh2iPfC2l3SJBd4GIh4F+7OgbUv297phVjkbKWpLTOmXhrVqcajYRUpPWsUgd0ofYKJkYE9uDp
boutwULMUDVfAHmG+X6gy0VwoGvntknkuyfthLNJy7HnLAhY/FUOV8Dzokh2tlFz9tYkM4tm8M0Z
Zf4OCNAg5COmejmVZ3tMcjrjiqvdvK8Xn6KW+V96N/kLT5fstYbUKzpGojUuAse5fw+n2mQMdjal
EG51kOcwGRW625Rl4FZOru65p7r3nI0FlycUyyN1V4yL86y69d5md0Bcc9UDl3LSKU3/EAfoq/dQ
/PMHtQc1FR/9s+H68yJ5LtoEFn/kCgctutulQtjYdL/KuAPQHv6FR+/uOHJcjlKkbFjPQ/ykO5Eq
3KdfLKWbjB+ym95fOzyrPP6kLjP5egsKF+zW3O9HY0qeIOSbf6frimPx21MBq00YS6VmfG00Z2Z4
BAG7dCgOmTFQV0l8uVA5RPyg0coHrwjlc1yzdivi3R7kJwU/6aiuA4IXi9cTAEHgK3PRQ64cL97g
H2Jfz7T4p4mDYIQGrx0FEPpRTmR89Cfl7toT0lZ9FRSPtGw4zUMAAwUaLkln8QRL0B38keH+n6bk
o8/VfCt0/sQ5TkadvUckgL18mUKSjoNGeqUvOl5TgycFFsjZhAPVsEk2zmBEDEA05cfWHOcv2658
Goc95siP2pdqfxLvY1sgeWjHVxPKPBleSlfvF84eVAnrIXgkPWV8IRRJdNSlPO8W/U4/4Y14lcd2
/bg7MX9egJdImo762UDrn4ZXXstOAeie4JmYlzfsPUZr7jg6XZ/LyNyLtgwQMEDSwTKQ+0Z1laER
N9yfLw/mZ8WRAG4kkLOubmGvyjV6rmWJUkFgkGQIfK4G3JwMeOQXakOKwy+Z88gmJmvXOY3L/TRE
a/euQ6ugBgT564eFdufaOIWjP68QbGvwsQto++pM/80jDqXXqadeafOJVhALraTl7MY/h1ZVRDw/
qT+KTIq9YHdXOzRrkXCyN8SWNwG3KG39wQalDGjeEnOPn0FrMKPXmBWZ3xdqpwEnvFuy26FmqRYY
2yzQNd0ZmQBAzQqivDQgY+29UbRw1w73v4mx5Yva/RXuh5Weq67HkEe+gwspRCCrDg9QQKIgwUhT
/WvbzE4YcmPTr28Tg2kyDCTupjqcCukNyviNdOIxxUF+Shu7JtSy36g6pjiOROGmViSJJafT2mT2
kZhE+AarWLe/Jn9t2Awr/uvJy6++kOZIgepTyHUF6ZmJQvjvCJ0A6XsDnE26W6jc6JOjbUtExmcK
fxjB1W25LjIYPftfl5RO7iMBVL5p6eZOB+GGXafOqkyZ6tJiH0IUPRIu7zWontT85G0xX4AKfK9x
lKkwljuDFigR94FeDUnB9QbhA/t3fNSYAxtgntCJBJ5ivpDa/PJBPp/NchS3mdGS65EWyCbQuexU
4COOWxtnR95tupJIAe6Nfi4HZ+b6+TxO0WpA67lufkjQ+nPhbcDmqBrFW54Xr9Bt/4+onPKOJ/IF
5Q84dTTxiL5SYWh1ZIUCL/otdj47cwWvy1rIcTy6fKMRUktGnOkbjwsqHCVraRv5uoM/2REsCldU
tR4K35oAH4qF5Px+C+prvTkyfy+16kxvBNb+kj9m39cEvFy6s2ydLLQGgMsGSr6oEu8NUYJ9SWwl
n4wENAWTqEiLEFNEJm8i/PBtonOakPeNjIg+3+y72Vm3tFji5g/BmoGyYF9RCuaDUW2FrbMRdgVl
lqr1sTnj6JVL5AxXL6O3z3LbrXsHaqoebBdr3xab162RfqEQ+Y2GSqycMgHj9dU65rqKgZ7m+5oj
6DMgxzwfCU00W1w+3YKGF2Q4QZ8QZB6DTgOBItjIKFH8mymttSWeqH2+mi67cvO3cWYWEs14RIkH
ubTEMSjOSZB9c6swAGfXQWaSIgiPkr8LFMjJvJNESNUwgJ6cETGrFAe9PrIsteRQ8Udoqyz2spqA
yfytsFz/nP9Py8Hmth6g/xMuOHa81KWC+KvCGLCBjw/sKxMUPhg4l6MHPbZzuEUZOqzD2uk2kcvf
3VsKpmQbwWI5766H6a7VCosZyGuolOQIrCx7+9UQXIaYt2FwNJ0Zcmq8KzoqsSwtWTLkOEOtBFav
pgDuNvpcDbkwaQABaV3gqRr0XFqvskM9zO2aZmHMwK52RBfk8SCxhNCHiJni8C5uB9ydXtXo9nmZ
2bBFF+W0poWpE7mjusWV1bXqh0YsApQFaBOHUBvUw9nRZxxombwx6FSASgXt4gDqcSIBqbLQjlrZ
Slgmcje+3YuRQy4hbpIK/L76UWOxH8h7aYBXdEUof9G4tzQ8Xjb1c5/kFbLFYKtl+8q+Ay1lgtnc
I5U5FoZwAx4+iSi2AF9WyeLwzocNL0E3KxF8hdVRVmwGWNxqtn5Jc4Yi1jnftZSgFQas8aqL7JN3
CgcG1ietp8l6vlCxs27SwSG5vu4/srX4dm6iED9jH5PotJfhDzjNunzBOIOMoizNViVQa6m6X8gU
GmDOhAJPocC4AokQ6LLGXmLJLgxeYViaSFGaZNEhXGv+leHE5wNJtllfETHmbh4MCrgEMHNFGEsA
YzrX+2vK06Ffd/+L/JpWkl+GD2fRF+t3iL6OcCHRinbxgCE2JleT3+3d5EHsgPECdmdOjiYF0FqJ
93YgoJq3WfU5sspDY4bAgUBfF4F2Kz/3QIxejdErgBOi/fyZBJp3TcLmj44X56wvk9eVFSLOioT5
0/JgNKiqgFtAs4LkxrZTWvnvl4aQ5vezNN+cAyEU7loRvbi5t1hvOBTVY+JhDeLCXjLWPxLE/524
o2jX9GHc/3jj0ku/6SxtKHfXjnvGJvGS/GDZqAveXtyPjY4K1BM25hU+wLvTppHt5N4uAu5kTmp7
3hKGjTL/7dDb8x0T148k2SbEIpVz8wbL0ASLfeOCvkXXODRDjeCnF5zUMKFbZ7vxJicivbKiLJNi
9HnWiDF2DQgidAsFBzInDiyR1PrGFc92ok78StHYVx7yb3sL6w8TukXzTaQGaF2RJsuj78glH/Q4
M38ub/kBtSNC6H8xX0Bu0Xb8GGkjX1wOVJSaREldVz61p4ZK6Jxnq4kZEKItLNnz2JUNKIabxCmK
0zgPbdhVee8/9jHAyW6C+em/6oKrELTsKZ7S4qPFUcjNOMX74RZFrWleTNPkb/R9mv6q0Pqs/Qz8
tIrLPHus5POF4wzHhXtT39naLhLjKD3l/F7XsalcvugI0fK6y8H6ot9Dc6ZDSrICEBjTN0tUALlI
Hq0yJMVarwN7ZPE8bIy4N9Mup1IWA3eN1sWbcv57zhNhjHfLk30CsESh5abLY3Hx58MAOA0BDyT6
fCYtYgeV0iXveqJmVfaOtiM4U07AYTOSrm1Ad48/ZWNymc8xGEdJk5yw9I3hZLQT9BXeWeII0MKY
vYSz+M7PxU5sjvKNfke3u/GQ6JWcsHVfWNVcKSKhM0H/NAQ8qOxcTLuaZIQT8Ejws+n6MMFoqWuU
Q4jTL9LKNDeK8pWZGSCriF6KjP9elE4P/OsH7w/2PHbBIY1fx1UPMt/kQFOqDe8sixXWMML+3hIw
mEhYEa0RJD0oyzb+vBOX5sp88uXEry0bJIyQBumK+j7sT9tVi5eaUoO54LnGDUHcXyhyOLCtvO60
2I8U2vrED1+9A6HLuSUT120SpJjG3ZnYU3IOA2A6vS3fF6GLYuM3IzFYGumLDxP4fmfXJSkfzGvK
R32LuBmNJ3PCvtQd7GUnYT7QCq2CbijBYSHnQ0GdUpMtS2AxIKSO8Jn/IzIviuLVPOwZ6cPHyXMC
snpImB7sbdN9JkNnas10JM+XtioNXTMh/CNcbqnMHteR+EpLPDL6GtIzZFdGPn/MvwFWX69QP1/r
/Z3TkTMDK6WuSp7FjOBRsNlles7TOLc+vmHci0Tr5gYKeSMDbUWvO0r0+3KZF+PeDAAYJGwU45mI
Nub5Bz4ErDgNACbysUbQV5DW9/iyCCo4iJYh8hP8UKQykxdwxbo/BgnXCiNYfp3FnrBKepH2uw5N
0gORAv9YokvPRjyaoAFI7UBfEBZN+gHEaIO+kLY5/HxT4UIcEBlldN9/JzSqHQmt75hwYoPoC7LW
V8ikTzteDJuEVWB6SB/mScXn6MJm7JXEaCFTp/4/REzmoSnD7OF8KvDi02MCvbEo75zavfbFX9xo
bZImHLNf6aaWzbddXbPDbMN+qOK9IUzZ3sVUc1bRkFe1dtcwDrtxmQvagW3kUwkTMkHWhZiGQt4w
xH5JUrxbtrybsmGb2JMl9pHiOtA5PD8BpjvJcb4Hxh1zw1O+q1OwYU3IyulUDVBjOuOOb9clJitE
OTk+Omq7GwFYlUgqLREh0Rlkyuyg0OzOoew8ZcKVH7tkbNhRhr9Afagd4tstsCr5+frqrw0N0Xfm
JtQC0EGCtURpiwBHDETeS7YMXjMP4m9SOx1Q6JmvjBRri7No6E6f5UavpqJ+EuVEypxxBXfIrUXO
5XJARnBrBeoIfSOA1dW80v4gZexE5c41JlOD+HHXuasFmTJzqJ9xaKUivjT2C7HJBe6wruO9T9/X
JUQDL++ylUFSONehAJ9N3AJUySwG0zHGDpzYKct9e/Fh9lDgud4fXHBbkMuCMFmwnwlpjDFwC4Mu
LxUixMXskQ7ylWa93+P8BkA2u9Pydvi2xDZochCTqjJ1BsGU/BU7AwD19sKlbqENk64p6uM5gYM7
F+VoSZUKLGsccN0xRgp4BAz1NaMImBZUyIxSjC+GZm95Fu5bZjl8DhbcvTpBd2N3XHaYmLhv5Laq
8yrAKe8D1wYIxH+N/MIyWtXnyfCZn0Js1RCZhDh6jvHiqFHQE/PV/6tTQenRpTV1+MzuJ8qaN043
901sOf3IwnEoS+CAAgVgzM+tStqv9ntjNIZZJHKK2KT6JDQpdW17CbFyUCtnJwYDaSthzbwUr7bR
CpSSIz3K0tSxmHbsrfcJydZsm6ZGZFpyV0YpPlWZookGE8GYvUfHG9TO4qdlULVQCKq4kwMVhCfa
XltnOxmvHCBcFBFoSFGvfEe29VoRVMv3mw8fFDQpVjCd8cWKwnWMBKHz/N/PmZllUH58A8jhf7TP
CchFyJku3GGWvvINJ2V09gelAFwI1HvD8/yrT3mBwiKUJL8gJ1C7ZXtMqsyBCjjsbYTXexTsEJMz
8E6GMMjWA3Q4uudzr+l+vd5IadiZh78ov38uH+kEKILsbybm2TowXgd07d/S33R6TAfKYfB2lRMg
jPxmouLeApMARexYx8P/h27itUcX1xWxlg0FodaSq1ZfbvWrMuokWGLApJydbfH8WlORyeYOq+kl
AVKG5+NOEfcqBLDU/pn5+rzUC2AzB9sf+eVpV8q6NsMvjK9dB3Nj4lo/MgEjUROlsD/L/nbYVTzF
TTvLeIP7sprkOGhx/22J/989p+fTYWoTKK0KzojBn+Qp8h+We5nuaLdYvplp4vc9MBeec3hTAkPX
8k31QMSkGhc1fY9iBh/oqLGEyKL00QszijgsNs5241e5RIyjVwbzaaRhbxDTB7oGD79mLmD5cW4n
zUEompn70kTqNDM+rW5y1Baht/b4lFzKoTRflZRDqyHtoyzH3oY3IQ0caZHfoTAtuu92+LIObHs2
PoUzOSo3u359qp1Gf/SstmHL2gkcE0KWx/BVfDqXzFSpgD8iH1Z+XwBd7gCI7bMhFOVKC9s/zydF
/NYPCe9U6w0aNu8Giq5+AMEF+GgRgjHpo2LOCNj07UgS0RvUSNweHvlfE8i7B9ZomTGxYqe0IUIw
itwvZf+ImyVKqWOGlz+Xi9neHlZWOKAMYzwN+k/U7hbYSdDz2+KIue6iyJkqsK9ul0KwH0r6kikK
WFj1uHc4tJmG+JoiQ64P/+IONhSNyaYE5PMlvYSoZktBDobwxvRMeZzxTRsOpXnXh3cwCr5Nv3Pl
ra1Cz7Ob6DqpU40c65SdJ01cxqgKAJAygMPIV16T54KvF6IhpLSUtjf3LPXJSnWCU4KhGhwEefBR
egwiXalix8W2+jsW+x/UwyBHeV8twVka6bRs4xl8k8OMlEgwY8oPr0hO8zJ0WOVnMKe7MWAGTT56
4YIAwpYe/9ZMpX0flRMCdDiCGqAgF+UGF3XXpsdAnWWGDqCp1pb1DnSvYIUnTVxEOTxBZBHgnkeN
0A3dfagfJIoBDBGGnddg4gthw6WWisCgZC0F4Hp4lA5lXTuoZqDHZ8LgoRZSez74FdMTppwODAas
NZMqM9Co7Q4JFOuL0q7nxei52ji6RFtg5ct7wJWb3789DE1FKKhgDpUxB/WMYAZbbyX561BuR2Ye
TmMFqIjP4y8CuzD1F0hV/LAGYI1C288s+LuLnX42XHRGdbAlE1w04QOTPdGrsiUBmxzh9jJgOp/u
l9SLDq2S9ovGMMNEY/IzPlRz5S7r2NZVVG3nOsxCssI5eRAI/rOso0wf4ixUpW0h+0RlpKwzL7Ro
x476HY9cul+thFKt9SlWzPQ8tJoLC5z2aeGRBfoZ81f1fTTEowZnTnVOxYvvTMZsAzb6opcqp9z/
IJKxBp9TrDgvOP37XzZjtGkeCSAPB1Pz30ueIbgC4t+FEvUslzCEVffFnjwxqaggV8ESfjziNGZ1
Ekz2dlWdVSoqnN/deQjF2/NRN0glCtc1aJTgrisrpVv1ONty1hBIXssx2F0QN4QQMrG1FKEg1T1f
klFbqhRNWy2ZygA4hssXZBk4zm1rjIOygs+hpa8WT19i4z+vNBAqqvCc2iRw+z2bVM1+zF+OceTp
9Z7aRYOzp2qI7ydeO6gyVlvjBQhFTvuQsJ8vJDEM09IE0ap3+N8YJgpHaPjzya3UZfesv2p/uhfa
l2ohKAWdEcqDLG8bHlNCCWvqK6oHkNsmxfMLwUFRXQqMJqwkHVszV6hs/2qybOzlVfSm2e6x0zgO
c95ctE+G8FksSr/+IBlt9T/5F7iikESujs2Xi0SAii5WvuGbYKMUorCeRc0EcY4QzqOc/MeQeeva
dW4DvfjU1nUexFbo4DW6q4J+KpMa66jlrqtSvF/bPNtHow7zfnnMaPh7E8Stfg0gRxgBV0JyPc+c
hcu801R4QShMrGUaMEHRwYXKiK1iY8lYsjUPmRf4KB2YAksFLgA8xdhs8xFZ0k6B3ZQepnELO8Bd
FSqhflX5FZXMg9KQ6keBWZBcGzj8ctEWrs7V/YCQ+TqDyzgU1VPrOjM14zf/KSrsLKHrikDP7i/1
HXohGeSZrFjY5S+lkqzwpYzit/Eo7KWeb6qFHC/rpCFKffOzkgoNQ97Gl7B7Dh3mGqgm/k0pi0wO
BA6xZEYRTIBno7UzvrO/PpDX4HoSjbdpVh01Hb84ZhkYyevLT4NzMO+xmpH2ltFG44ue2/pAbGBj
9Pw/PigmcR/NK/+Tu1M2lVOriMrVDa9wLt2LnZKSr5MQtmDtEWKJUHTUtIEadeOEAVdbBWULl9TZ
TFAruzRTI3Ejm2GYiP72o19SJeEIJzYyZBkCiV4W+2k4KzVwr5tBe8RMEok/jx/ZjkXTeWh80ZrF
OLtPMCZAKYb28N2k0JIszKBeGqUhPNEdN9bNga8IOFttyvucQasZ4fXCj/oR96zErY4ryeKVUejS
K7ImSuBs9Gk24Ith67hSP1Zq1JQVXtM4qYAeXk3d6b/uHOKbAhg68LfcnG0tzCI7oEgfO4Npus3R
J0kcul6UYteTEJICLO5nY8itR0T8577HqJFPEOkC6yazDpML8huxSdTGHr56meYhnZ09PANdYB4k
HYl7monyfREdqtPq7/fpTP8dolFqUUfiAreFkguFDOyRd7SW4IbzM5GAt1XADsP8QNSG5xzTVdm0
1AOsTuXbBp3Lbc2murDRVQmBrdgQ5gZ2cblRm1Sj2SGT33Bpov2+iErS7auEdIKUqUJ2FjTO46CO
VoU8m6+6G9OIq5oI3hYk7ovNkZajblOoLL97d7fA5iY4wvhFRouunT0e8XZ9fyhtxU2xN2ahPmWO
cKjpRzqhmiI0YpOCDBossvddzojnFyEXB2+aJGRczvQfFVfjUifs4WLFjwLFfi3O11OGjjMIcGMO
fZU71TogWHOtYNrBDVryrKi/EFITsvaebtaM2gNlElE/nA302xZzgWtE60mq0CWauCu5Wtch9nH9
rCLLI8ZuuO/AuwADhpkxyhDLnXzlxVCHc6/dH6QLPj0alJla+dXG9yA9T8y1KA6Zl98JWIP21P6b
tyduvK6hmQuxDPL6qT/sWWYDXXzhwcHUjlhVIlSGKJuggVlX1SyQrnl105brSkEFWRmBbvdvTvgF
9qNcS8STupTjysUACv2hMAg0tPO/UjJdhscq/dsTcphIpHzzbyAFaQwjo06snU2+iuVZH/9rXAsk
1/lmws9AnLxUuNFBDLsz08rSGDSQL2HOTJfH7wwhiYU7HIUzhWwFTTz6jVbdfMD79AiPFucvbLwq
q0BAnW52i/kDUIQQ5CB4EoU1/Zp2i7mzwmZCHOjeyNkYHj8toEvKa8uoo6OxA68g7JHEO6KlfzkI
hdNBgdhC21k+Vc7P70A86KkR7Er9OVAu9+D+ZmqsGXInIvAJ+zlGt0VnrAD6rFwfsWOC/lUZYbem
WrnCMbHkAZq2m9wKC3B7TVN65xGlhJOblevurXidQvMEqvmUkaryQv7+NC7Pg5wOvFcGi5DXWjdm
KEZ75MBVr9VE51PbsQFKULQtu8nGwo9VW56YpEJhsIbmkXgaHnGMESHkSO543x3HEMBrxCAvgGkd
ENB4TtRWdkcPpIwqksvmjSqDrPhTeF8pTjtHL6hJecpGGeTKDAKSBiikAoA8AS+9q9BNpg5jG5ya
O2LMy31EXYdWFH4zbn+Q91Zzsjaa6+MaZSi3m9gofwWstphAURziOXNGrEtxcTH+WG8w8xnWj9Ev
BB/OGdKlBnVsGKrMsPdUcifQwY1IcHHF01lQezaFVn5sNDRLulYfdi9yWsqtuRme/bbEGtSTDFYV
xQks/m3C6y6C2gtyULg7MFaTpOTV6T5AZRbHHbGO+f0uEeXuhhKDeR291DZE5SQJCn27cW2xf9yO
e6RTyoNb8c1PIItgd0cxqUI4UWCSi1LNwrHHuUR7qRCALLjP4Zsna30JnqK2+rQJ9ju8v1U2KcbB
fVzU5LFiI6wraK8oP6tgM4tPJAHlaqyciVeH71KroiTx/JypqNhEDkHDgTTQIxOTYjQjV5IxYk6B
bhVvn/TXkZ0eDyOM3dl8YZKpkRECzUC6eqOItccg+DFrpa9jwwNYX8CYO+0wNAHRR79G3tqtx6vN
/B6oEvIdyqmK+h2Hd6/lhlrmGQ38kUzp8hb6pGjbOnZ3H67izeSFnkqBWm09D7S/yNP+Ts3HYuST
UJ9OeZeDbbfdngAYCYcVTYWmxzN7OC4DgPOgHStGbt8sUUH3nJj8MBMNqE8S+1NMpR9aCY65L1Hh
9T5mlK1LR0HiR1qC/n64tTStFhL3b5MS+Pl2q9jdNJBxqsIDm8ByjMYPzlD3KMNZq+1ASsGXyLY+
1yJOUtdgJRfttXk8bfK7AyJcFc7P7Fz0i/+gOqfslhxjpHNmaO8jeqmSqXLABTxwxzVHgE1EZgQm
0TAEFyktbrJXHOZlUKwBtgIMNdoGQH8cgN4WPtxXVyAcQImg9aiOsD2wdib20/J4JFq0BXmre87H
jtGX2r4QaLWZ5mjUYdtGfz91eXmhx6xHqIxW8s84D3vlkEXe2AXy9DzicVr6MQw41ufPU0L9IdLE
CkTldhc5ZHN4zO3Mu65XekNP5PDvE+SKaUKVtVX9CALPZkImfRSjgaDdhKtCbxgeRrZBopieA/8J
MxAT3+gvBKQ9IoS8JAuyGHUS39yve8mc9LI68ksxe0KNy6BBAcQM3z9wMcdrLoAeFn70yXy/DePH
ySTrxmr2kDfOZQWaMifH2zmOrqJdl26pYc66NUj98PLoZbGL+mmvLf04xVK3ThQWBt/5VDl3pNkH
RyxcVLLH8lHCDp/UXFf7ZqUtWOJRPEPsaX8IO7x9OYsfMHQWY/JFP+CrKAcsqdriQO6xHJ8SBKUo
OBGFbdK1PNjBC+oUzh/UXt81b8VhKOHvNag1WnNYxw+QW8maeRAGOcljcwYV0uKbHXT3/m5ThTnO
+GaIcN2cg4GNMp7/HUGQxS3qhY9XP1aJeuhu0xswnEciOx02ACibW+DarGJmCMtKVVssNRCLfqoc
qmuRbT3bJIZvN7gHA2L/V5fGSi7x8QXsJvkd/Yz16QY+Ly9UCzRFVyU65s+PRgvOKozSwZIePCqM
MQ3I8209hwsr00PO28EPamoicoiF86WVllEv1h37iUFsjDBSJ1u47nKa7T+xz25bg5Q9yRG8g9ya
mgp5IrjmumFBtPqQCREeAWLWW6e0z0zxSA8q9E3nokTdUolreoX1gHJrBkQ2+u8H4Or78TFmwJiL
oe1fPErNTFAYdbTze4Z9ax4lF+9kHgwHfZyWCzONVWr/q5df2Wv0rYqTXgkEK1SW1vVhiQnECxj8
vLly4a7Av8xLp/ToVqkkqGyz4JmoHG9UaJhfLTskkTu0yWNXnwQDqZng/wRCt5jqWdyVIuttNDaa
/2PS8SRvY2Bko+cXZaGI9vHzBjzPBlOAJit8CtNUBTZeIUw29P5rvv0MopSkXQj/8bGN8rHpo9Gv
6FO0WprVu3W0FEVjEMTzQNQD3+frwGDEe+CsIFHHfDE/sKa+cCzKbn+VGvDtb8TE2eHlNOunYcnq
eaYV9pOFiRoN369DOvWqF2oJs9cgrTutZIt1KW9mVjgLng91dkqFMqJeHhbkYkx7eS58KguuoO7N
V3W7kkyaUkmqcbKcT5XNYfgu4ojZteWfiz82vjv1uUCMJyxuwzYFiqvNXSvWM5c3fJrn3TsudBJR
J2jx805rLyT7KkhirviHoaqXtxIzmQju4f9kZDaHetUFZAW//kfBLea5syTvhFcB9S62+83Q/8oo
edSU1mWOyhWtEQ1GBr2+ccewB37DoaFWONfSeiT1jBkdyeG8M9tFxiqgz12DGiK1fO/xQ5ZC/gwP
X2Zr0dGU1i5Dj999kJQYKReePxZxv8jKM4OGvX9V5ZXyU9sepNs4UOgT1N33iJm9NBRpRxEBooi1
9iuTGx7VmYwstQkLK0cQlQA4Y/NmwVD4Gidb+dUnCZ4VoK1PxocHvM9RZDjJl/sNyjIuy3afGqP+
LEos/raIHfvXq4DEe4f5AQYbkLJsPE1y2zIrSqLGsBrT9SXcsdyBNa9z2JPgpSARrk9W6fo5BQPr
/I/BGvoQKI1Nbocm2uoEzPTqlu68MSkqExLv75VUMRwX0MsuFbXKTtHb9gtFWsYYXycJAw9cZ2hh
x936V5l5VGDsDEKsvOsoKYyTo1wWp65XPNwb/xycmkvXpiOrAgWcWijvZ3CYs026/iKd6qhxDK8o
9JFvqRWRfYoANZjM/pYvXWl3yPfNA0XUiHD8pxsCuKfxxazILP/1iIgZPaWWNvYT9aQBQVUKWcHj
8qSVx6x6vg6xJMrUEZixFZgsTyNmF6+IxrsNycatO1y4cQ0ycsVMHMRLQx7pUVL0o7iASK4ypKJP
TK7IYIBvPTctHZg/lFMF502BdcF2OTqmCDU1nb1GHEfm409sQCdGCXuSyBbVOsCtyn8b1Obh5idK
jfDGet7uZsdC10wapOUJDQ1D8891cBSBNXTOf4ck5smIRwoUVdnghrI2FDZqXW/XiVrMi3Nlr9HU
w18K/jyt6Ho8cGe0fqOXpXt7E1TlzsBCATH6l8siIBIu0AboinO7Ubc8EOUff2Al8EU+vDJeIiHL
gl4JLc4mOgfwvFHBkT8SNsuHGd+qH6REsq+UaNWeGW4t7X2wwM9Al+ac1PHnD3Xndwzi5eo3iOb7
cZmdB7t2QGv1HZenlLCitgTc1KfxW0wEmbjk4ZXxcYK5PKN3/QGmWm2RC5bjzrdtTMHb6m29kkgR
gSR6wlmBxclHDNAj3Qng30uOPybpEvg6/zMncSMJC1zA+rCbmkz+U+4C9BysAaF6Bkni/xAxpG21
/AhE9i++SMnlexaXkEy9trI7bUGl9zw28FGzbifDX09bOfITgXRnb5YxW5nCP0KL75cjr0U2jRjE
BkpTESz9mnkWG4NyIhT324jPSCt97oyyCIU5w9WGclMA9QhOkWxJDMRSTuFkVIRGu2cp9JrS2UwZ
mvpoh4FlDh0k4AteUhx8wl3YK+QWYUaPrDPSH1UGhkUQyTsVxzlroJJw1+EzeHXdCvlKmysU2Fbj
m19g95LS+iD2YdXoVRps3X40vhS+h2aGlIX14Ur7bG7gTQScRKQI8xGyHfDs82x2HG33ssYc+dMq
bfN0glH/lmcmq4/qUS1T87ndr/y1twDvYDbYbzFv1/TkOUciOA9Xchl/9AJV1/TmTuttq1nwIEhu
pdt3flMyTbLqENfhRpu6PSOW1ExubyTT1Ina1K1X6M/9HY/SQE1xpHrc8/0HDIGymszRsTwB0w0V
VRE5GXdjtx7us1eqbkuaqyaC8ybb3ENg8i3/Lhmo6zUE/Y1YW90QzkMU/LoI9BhCVypmyzDzT/cM
A9A4+2JPRpSGcNb457owMcbrunJk+Dx9XE4gDtG/ygo/TazI73T4RSQy6TdIEprRoeNJpLJluCsF
TBBLMjs1Xs59MndsG4xrpjyGC/pyTbwwHSvsd824MykqQtScvA7MFdXY6JZ7NN6eMUFUHUcW4XfU
9v050SALgDxmiuCWSj3IcVqKnKBWIqDbOKyQQXkvb0aqSRuIeTXXMP+1NcNzzxUbCUShHu5qFoxz
5fIT+TNnb7AyygV9gjj9ZAGjtFKC1SrOAzy1YkNmYh3NlXkIp978wNfIXt4kPgYdBgFT0pYKT0Nv
MMG6ZdhfK+q5887IwbCV77uxvoHEPiAAx/R0qg2g3AwpS5ssIhMnZz4sJLUw629/0wr37/nZpsJa
pppNvV6BHNgilkbMniZli3z7dmbwZ/MAXUfqS84YWz/XZMbOltAMKo/ZBHrtSSZl3KK2LAATo/Gu
YfkjSY3l5IvPUvcxwEaUEhR5Du8YQuwgJDpX9KP38eU7w9JXHMC9xgBG7dtpFh9k/DVUW23Nzpym
oyFWm1PAyW4xgCrkLBBXEed3nkjWm8ZvUZu3BTpzlKh9yuioalcuwD4/hEaFArQYe7qgj1eXvyV1
kizoG8HwnRe5uTfdI2wpYg6MofuJlUatSjmZuMR6plyf1vDFKzqFOqbR6COLEcA2JTovZ4sHFP3d
iZBaECQ5pl3SnlhOqvwLjuEFf+Yw10VNdCHlgXCpdQX+TUfuR4vlZOZk1+BMF5UGaGFwZyRuHLGd
DzPuJN6DtWuuO8Lf2FJDUhZD37aJ1mATzDRxSCzOAWZJHC+4qCvuHHOiY6CKQmfW4ARYmo2i+YJw
55KPeibp/tvnK7AR8g2KMMtnttvapKfbk8L8sjlZouV/gZkHq/rkPIUQhajnUtd32EHMlgEptFcN
c/5RZ4UH71kUYM9Apkh4QhVytr9EYDg86+GIOumFC+wKQ2xfAOqJtSRQzPwe5FaU8+5jTeH+Xwv/
Cgfm4ukQDIb/B/dFWYMwGxqHlv3AwBRtnBnqmeGbE4eemYRdF/TRPOw/jSgSDTXn+6o3TvmaayL1
Jzid8nFDhNVPBiUQz2CQThYwPAukdv+vzbSbZJbcsdEYTtmqvycmGAf/xjYgmxvaa5DUc7eYxKvk
TWrMJfXrCJWrxywgL1mRoFDmD/vOX1lowo10S5bvJR+QQEWt748T/QnU5SnFPcG+d74cEapWwlFb
buDkLoW3ebY6+xLKzCIPVyRUxUL9X1+iXnqRIQX6bbB7SDGdwfFBlGAXiYlVzJLIIwPlRy/0Jlqk
J23FTicmXWHIZske5mBx6p7R+v3v/rl8lvTpKYzjkM1bnoBzmAypH13QlVF+5XSw/YXga78cCRqH
TVUAFEaCef5aDhBvbZPjDcU7bNDKy/Pr504PE6k0FWVMUOQv+9AaxruJgIQF45TQWfsyKnNltIOU
C+nFODqaPpyJftTMcPyYMAr8ok1SUtxP1CHXk+RjBoji5etAJE2LCzKVhPDJQWk2V5OMjzi7YGqQ
k8IMrf7J0L+Askb1FcZAfgBWCAfJkXnok9JEaOU4HCQn1z3eZAqSN4mOx/6ZiaoAbiP6W6Zy2e8c
8cK7zzQU0hMR9bJfjWnC0l67IhdtWASRr8L2JVgUrUO40yP3sHAPN0w4wrQPUJj8yZn+VHwdghnR
FjBRIjC/coM9gTqjnn8k4rQsERZtbo8+DLU5iy4qj/wqyiDY51TWUwdebiorLpkAoct6btNaCXtw
mHvwv99emm3puPF7UtZKP+TmvirXZYvPQ3lBRkgVdztvTbAEH2VGY9PIm/ytnrjoE1Vk6BOomPnT
ugnMb3dr2RQSI6KR/MgLKaUme5zNugERdjO//d1/VJiM0y8t1RQeT3Du3ir6QGE95rSKreWLuJkg
vRSwFzh09RqPjYbKEKmmrPt6FZemKNYkC5qJWLl3I7tuYN4LuP3SHEzY4VN94EAVF57PNes41YPu
Rj0G18QLf797uNmqgtRCIMmNJrQi46ccsq/3M7XEwP/4QHRdkGH2950l6KaLn2l1Td42TZiQ9l0i
WEFgPr6pO280baL5NrWbPtw2xt2ddoWEu6wHm4osj70K8ETK8v1psVvjCoBWGXklQ5ZpFruY6kDc
bVSScefvEc7fbXri+O5IqJY5JSHx3z+MTn81f6PvImRM8Dc1CVhuIo7UtpHDD7hthVEFGX7V2JDi
FVoYbEprO15+UxR3SYTEEVaCgLG0Nd5pV9JyO50a2KSYQ/9ncu5Iq9WFc/4iMhvt+rSB1s0OAkJk
J0LpEWIm6J/JAxb/abN2WNSCXfHS6Uzjsui3HeiiEioCxjHEMfzBCA1LXz7EBmlnvi7oo68642yE
K6Go2mxKH7qwlxVyCAxPz4sGYhhesgCJ5f2fiSuDnIwKUYGxJJmMN9z+XadBrRJLlkCXdjRjIebf
EQKFE7Ee59beA8488QHiGGpIj+ImX5fexqZfHeukbOeERIUe6NEn/JtE/4RUTiLVbcU+t09vIDB7
fOtGLZ1ieDXcyMR+Hz2twm/4sTawDh05dIGKNMwHJdIU/nyVuAfLtCMO/YW2n+RDYEinmmXXD1C8
EuUwMLGP4rBROBkGP6ATZLsI3JFXLzS1KGKWU5sROfe+o4PLnTnkmMOtUnNaUIp/ozHWl86yFsYW
ZVIVUsZT5H7WAm5WkReQze+VHiiol/5ZlvoUAzPLlzt0XCDX/4SWr9DNSO2ko3oWfPPcV36k1SOy
G6xOLlMm4djJe+LVOnMoB9snj1eFgZ0pnVDF7ZEA6gH0uft3GmL1JJdKn7dca4r739c1Xi2DNct7
TyWu8Kozh1F+/54SkEoApFidS/LHzW2X+t/XJC1Kx+7czpSsceXDUcTHSfpkiF8eGSoPag1b5hS8
hMDH40EFNvcpA0dydwQ7vb4M6w8a7GfnXKJT+fMeqobIr3VadU1quf70mhgP2C7jNVfyzvmom4Pw
ZiyPL/VVSBgNe0LLBPCUrR3t8WW2ZzhXAPO9HE/gF7h5K5EjgpJeRduA1zUqOuwZzllKSV0eXWDV
ox0J4q/OyAixuAvVSCb7tNmJLhzPxsNzt7bWHUIdlvsk/7ef2ahycOw2ibIdKDAeTmoP7UhYQKd5
pRWBd3/F87GQAxbKXQQ6oanmBwWCWKNxT9z8OYw4uaxqUVkuVgqfMS+t6fqYagEpGa79FKepCoBV
ZWa9N6JPS4I6p1cI44itFEG/Rfsle2iX6i1LihC3JW0dRQSv6umIA7nX+Ltr536WzRFWzbQGVsLg
TFgjVz8528C5t1l/MwxlhJFUvdQyxDX5bfYTUYOAgYAA2obO7g7finIU6b/vlyQy1PQPvkkUMQxf
de49w2+2tDfI0mipN45c+mXgcjwRxnT5zLuL+FmA4rA8tjEDHpAv7ijcQzJ2AAGxLEMiRkNytwle
NLZUhi8xtra3WQcPdBXP1Rbdpy/ig2UzCREqOSMNAg7PIFwZlt9tB3gjyokeiphO0S3eGGFAY0Ey
H+SWxhPhAGdvKFEK12F4pMitBBaHWpFCfqNCJWm5rvR2Y7zFjjp8HPprJ4Av1CdPcvABjqUOdfFq
A0YFc5xZmdLUroKOrYhyg6bbWTtSXeax6ZZxEhTCvaPMm8bJy0LWo2GA3ln9VpZ/tKmjUqM6qAVs
Odd/g8n069IR1Vlsd+O5HSushRxiS/iw42zIL0d6/pXnz4OD0KOW9joyDaLAGHP+WMO/a2Dx1Uzy
K9Cec/twJMWbaO8EmO2T0sDtnrTQRxB/o0/lESxA5WjDKcGNVPP2iSlOeHRLxB9Lx/p/GoVmCq4o
BiTvR3omDy/77tGYx1DlaCJqYtoxB7AvhyHdnZWdXd7zrfen+KwQuFoYuANT6z8Q3kKShb3Xfd7N
xb7bJ0Oxmo/VFws9y2kSZIZEsApbqEsX/r+Ywuj9HnoBhicogXP1yi/mF8QNJ9hUtVPxfX0YHrfz
3Avz+phX8HDklu7IGW25VNB3GnVtoXfbqQK96fuSI3c+/r/6PJUQ5nQ1yuLZt9kYGg+ZO+qnTWJy
ndp5bpvK87Xn2/d+UGnB7t2JiYL39kYT8Ks6ctk2skbFu5YObQjuMH5ZKMAChS/PP0IhBRI/3bS1
OEX04oOkBO0iYl2E/LTpfhuT/ka6qI6soRfF/zpeszIeBpYzoD0VXuYL88Ldt97Vl5XbQmQwsHAQ
ddab3sIe2z6nzryty7KKqA0DEWOgYqDuVsFz394jhVqelIO3FVzibTkvKJeo9M+eSkQAR2SSbO+x
Uww8hSPu1joZBxsITQ/KAmXkqw9AHEJL5vhVRlD5zLz2f9RyBnGxvypH2fn88K7rmzRCF5qTIb5m
DunGAw+IMlBYCyAbIB3hjd3AcIP+R6lQX6mXShN3/3IknO7/Vtp0a0VQ04Y7HbytRGMpgo1YWV5H
pn3HAFTpGdfm2hxXFZ+WhTuO9CxbB6i1qC9LTHMBPtbnRFlZQ/pFN+ZSXomPi0p8laFKgtX009kV
fi9sQMDRS+qpxE+JMDphxR07WYftAfqezX1c3ActTzPIQsOhcQhO1EQwMV8EMlkfMoWlSeMXiP5I
sDxNJ3ek5cV5dbShhPp4oiSUf0MAN3HT48E8QLFc5yC5JlkqVsVGngOroo1Uebjw1qR70puDO+Lx
T725BsSirYbDVos9KQtF69oEI7eIQkamCaZ3wFq6xGT3WvAfm7tqr4QPeiYCcaLbsWlYx8oll8mc
sPHKs0ByKINC3R66J/ji3RQXFaqb9dSW3MBZSdd5pp7f2daQnzGoQGS1Abuz+08M478KBgMJtzvF
qF+qnwApsvpK4RiB0xSJwFtbqCM2e1L1Yc2oXk1RkYTv5fiNm+RmU6HEXvrtoFz7hUZtBBKgZDtZ
QC0vKS06hxRgV27a/6NSpHEtwp2xwwF5aWI5Oi/Z28odBM/wqJVOo2qS0B2Plv8NuSJKPkgBM674
LQ9UaW5K7LFN6t1gXhClhqMpjtzlZbmKaYLDjZTFlo1Pjr0yp2/PipnhqoThhUHY0rJcePCV2sGy
4JXUp+YVLq4mu68nQd3QfkS0UZy/eS4kmyb96bRplGmLwpguHKGRoH1Kjx0Y/KFEdD8hZA9XSp8r
bQVfI2Vg/8kH0c73fQK2tZkLOePWwwt81D3krzJrxyx/YACbsRvIT+bU0C67ARyd78B2AWN6TArz
wt6hlEqKWZ+iIOX2Mc8N/iblWLNbgjkSNw+Xxtv0Wq/sGkwNEgMke7je73csuZgS+m1X9fq1e5uB
JUOeayqqHUio7dnUUfA9ZYIDSHzaZWOFh5ECm2XSXBiYihnkl9cnBtxq04Az61eUrNVSsMuLWCJT
Fk5CacI+TU2nbsnYBtus+FwlTN2jT9nR3PeahjpK3dq2r+7S8jTEBIQ/XBCxu/zGlY4ksu/hwKfA
Y9vsmmdPVL22IbotrgkwRwN2bd6QkhdiB1hcsyWLCNUFGsUsfbTxMdgCVEPCLJCmw2/mjqNHL3ww
zVkELJC2AgOjyrVz6HeN8NWCHs335xSLbouMu/sZS1j6Ug3pFtfLbmo9djwO184++9FGrdeUEiCV
vGj10qFsP/V1uExPllz9ACZDFNpgO7s//xwfIj251l3p6GyFuRB3dzhTTKu73dugz/P474GKJ1LR
WXP82MZNVUn9wN3/sdBpI9KNi3KcKTADdMWJOwSX33x/I+Muw9EBj/4Nfi20yqV26S91MfliTnKq
Axlhm9TEeyPUQSwR+yykZZIbybUZjwBwUP1dEtFFUBIzEH8C6H2yJnUv3P5gGL//w3flfovHFNRO
a6wC2rasIwiMzLhfkClvo/htAAzH0xk9aV7sa5pLJ2wYbL809hk094jNCSfqnA5hm2TfkDRkV9Eo
qdrf/K5QxlFCKSs+N5ymXIjGghCuyUdTeomE1tec/0gFfcYXMnlT21BnQ2qH/A3GZAnTv6Od4+oo
eBb8BQdeQ8F63KbTnGwKqBSxfiYAb21CRzyCBrZE4Dedhl4763DCHLE7bXOSDfgwn4TM3Dyq5T6M
keKHltwA6QktCrP0g9TVD5YUD4ZGU1MBn7ntVBgCnhB6cmJv41Vni5mw+bqm98qLAkDR8x2kL7du
epVdcQ+tmIF7sNv8zEU/nwPCDhaLv2XEDB16B0nSG0PhunJx16aeZLdq0s1VCeQ6CGrbwVA8EZVM
xEevVBneiBUhSZBmaraDSVactFvzLSzek7Osx1H5WFVq3oq2HLJ7S1buWC5YiW2dqrII6Tjfzqmh
rEtYmD5UWrjYJYriLGcP+4TBQ9qNGFeeG6FtOE1koRWFQ5PgGBRatbXfz4bFkp6O4Ohi2SZYoHOe
+sjTbxd1alH+uJxiqVrAt8G137QH7FflsKsqtYkKtoQTcG68n/hkBlr+fMeRikF0S4W5L6Dg8GZn
o5gPZjRSaYrlKC4YCCbt94sF8i0i6pD9EzitOzs+xZuxW+Ru8ZoeXWTrRq32NtsiN9gOLyf5Boti
jlHR4XiUp1F71yln7ZUvP9FZS+AkocTXe9OHtlFn1BAU9ea9/V5CVx87b0bP+am5FY+rDiggLL08
+38ZHNFUIKQqJqH9cYoeYLrdOV28AVYLQeB74LBS7TjjWrlRSZYZeK2Q7uwtUE5CDG92GEAKy8Q3
Q2g2WWlNZ6vXcssa22Ob67F+vR0DYiCNvRw8QtZFyx5f+eF7MdQ6NNJrX5/SkdvqtgkTntofxvEJ
493pRDZTK0HMlUpkjMiX0pZRl7Yka/ajIpKs9YzzEZcK8QZ6w3b5t48DmdrwHPkFVM9HjLsjuJnx
zRCxUfGLIZHZD7HNzXpqzx3ibomf3kM+B8/1dsGPBrOT8PwvJP1Rl6LjaeYhhpDLZWrJttQAQelP
D9NlhxAUkyrZ8oJHx6rQfOI4LDkhaOF1YbYZV3MJs69ekYcyHYdnKE+K7tPzK1YrTMnOLaQhjOZR
cnvaornGXVG3h012TDWOsku5vRxUjF5v50c6sLl6XK6OHnvVsw6l3XetoVTvdI/2Ok1IKyvMgva3
WeeaHg84GT+BoOnca47eYYKiCOix/edt08Z2Amc8wxVcbIbXmES0VGIotxTieMVo4DD3sCKtnKgL
Vu32m+ikOEh4Y6AG10fyOWLe7JqMMRMQKfm1NS5zeYGkplHFHRrJ0rd2beJn5CCHVkIKUth7NNGo
uwHOLh1t1Yz1ulBnLkh/9kxgwHn3jZ4kiuJVGzHMp8onbBkQqtxIf6houU6m15jOsTslMOdGn2Vd
Rps2uskYkL9OJsfK+gZGr260o81469nzWYLWhTb8Sai2zbuQkovi+zW+CJkXVuxeFLahuV+IPe7r
N2mY+WZ5EbdQqL1ul7MNIWKEaXSChbhznVewZAIDnmoXH5o6nI34otpP8g26AklqKZxnjm5fqgEn
LiDLRzbEpjtc/1z829s5sLENRZhoyVRgOnhcpqvmwKkGFg1n3AR6GJcbiiy2d6u6xLgxVyHJtHsl
iMrzeuumWiSNPdEtaCeq64HSycf448Ou2UTXqzAQyvSc6RDqbhz0RqVn7rqgJxAzpSbJyg/caPJt
XI8Bv08ul6TPtst0bNSVF81JgG2MnxURhGX2t7vfSxeGlqJ8HYdwdOdoD/3y5igR+jVacRLJaEUA
1pH1LFSDXfZ4THhonTk3R5DtD/IJ8uesYoWXeICfjTJURqvR5n1lb+R9PzI2ixQwphIChhBQJJNF
CD0O3W2kA0rG/GC5/U9dI8prS5M7hHJC3FknztscPJCOZzTGJW+D1PQxoOn6Qwo51pvwukyqZid4
pa1y9BWd9Dg2hjJ+6XaV6sNsH9ItBmaIiy9nIGz8jITfarzDSeYeSROsC1injWad7WHf2f7Q2Dew
8N0GyYumF+xxHeM4t2G6iTre/RPIRkR74h9COdW6igQ1GdJQGq5OXJyEjxGOX9qsasDLxwDucmy4
MtVPnKyzmqDRR3xQ8Qesu2oqiEi1x6Fc11r1W5qfjdPczaArcQejhsLYyhtudhX0OH0E3siL80m2
22bC87hxenOpqlLJQZo28X5ab1cYBC19uyS4RSwx2nBAdplCJDDr31YEi1Bv33/wgygo3wdXZP2T
OlllEJPkHInvdiFsrE0UmGSCVEjRyiM3BCul/XMdDFIQeLWGCG369rbMwDMuI1QTAG0sIUm6XeP/
PM9qsxlnO5/+l7RiSXvC1VWnx85lQQTnb/TbNb8Fl7pc1amv43PrSIbGy1vTlaFKYo2tK6inebSE
QjyJdFA+MCfttaF5dv+g8MCEkUbu4arCcPNcORP4DoPi8QInvMPC6mzA7Nm6WIb0YmxZKdRbMJZ4
Z3QkgDRnf6atZOB6CnRAeVdaSdpXxnonIKzG0wsavg144rEGuLWMEmatXPp4VBbGRLsq+ERV3xLj
HZRjAwuDjB5FLXeUI+1Wq1z+i/oovJZPatzJopgxzE28q+DWrLnRczwrc+Yool6sYQXAsiEBzHZa
kJ3/5ReKU0aIIgFdhTGlpgkxIvWjHrKXQskKx+Tt4Qut5wnD3M7LBrjvc3NtfwzNBmYRZJsI/puz
jZRvlXHVkT38CzwosJpQxev0U/fB6hdAGXXHWqLSHOuWrN18VoESoXJipHmLhe/GuhZINgrpRKPx
G5ryRU62c65t/qSfyOmpTKWcYd79HaqCn0tu9FKYBqPCc/rWtL8aRqe/Guu4Pkg9B+3y8Vg/jgGT
kqB8gJNYdbzJCWjGu6vym38tjpiiJrwLg2unqiYMuKQm5BxTNaJJBW3dQqxqWi4Oo7O1GOLqUDLI
qUV01VTIt3edrMSmCpmzlG3i9beRTUOdxCXRHBmcHAiANP0mNfXKElCNu92/CZnAWguyqEeuUNGr
sKhImReYB4htxTlOkb/KJeIuKkKzRJuOyjn9MFn9ojRuxyrWQKFLzF6E/bc4lpxdR7tPsYupGSXC
kpA+JuRaSoykYLoCvty+na+1WCDJFH1x00hbuDcqhfnL6LJ7M2yLDfYy5NyXh5V30bNbJCvIBanf
9ukmZwPWzsV1ULO8ZrbNN2YkkiVN+FysmeQVQdaFzJSylY3gKGp9CReyLGOFYn2YSbFtcaHVpKyU
lIAUI+bppvzOtOWX9kKSwksmBNgeO1xBp1JTzpn0Ktc5DRbN/OhAEwlX3rLWZf1l4XLnSq2pBs4U
dmba+wrXGuOoNjbg/Euu/5f0Ey0cKfLzbR+J+KM+n8zCKGTC35RK3SGjdhjAFFw81BBrJ/mBBT0n
J+7jvGjjVBY3CPqHt1xShn4dcVQitNXgI4w7z0JMWNI2lztnF7WjD3DqBGfmLDfrPK+8HZEiplQq
iQaJqtxPZBEGfgqB7i3sOc0Ure4barZOdsmysnqmLuSYyy0Mw7yohc0y4MKMUjaq1wDqIKAx6v31
S3otLdnvOhF9GpK6+0GAQBlVeQnowBvM1OdaFQLAA6JrWsIPqtZGC+y6XYsLVsqKsE7liv5Z7OT/
DAJnoZbCas7yFKN41qRC2wNlLSmzwhukl43p8xuh/hTypLMBdpMrc3FfpTbGp7dya+o0aw62ROlD
sjZBMYC1VScnRX05jRmAo4N4Z8e9N6ZM6+SzXmV3B1tkO1WH89bVPuKWSRT7/nPvz3MLDihm1BR/
EX0Q65ZD9/vGW5LOD1lJPt/QiQHidjEJtDQl11Ovpn7YdIFH7cVfbpF9PBWxgq7n9YO94JWNa+MU
j0ayZltUF6uavzwMotQZagSNoVa3aZ2GkqQBsakk/cNUFen4PRObYudrIKOrfZzZNpL5SOOzm0nG
+PR+rIP49Li8k7rsggSE8NWxAuV1Hv6aieR0k4VhKEmEP0+doH9nem1WgYXz0r2Yq5QP+tLzp2UN
F8JndiJyCBkbMycpmwQa/PkcVMfXOk7NAE4aGhOYFCBH5rSCovZDQ4QQNzWfngqLRtq5DHXDMIyj
7R7N+oKAYlEuEsCs+UoQVRs3WGirWs3EjH4FQMvNVwTZ/OENcfbQeGDk4YW1F7bNsmcGbNa1BZ+c
2Qapm5vaA0jCSqL0IlRBj0Saqd96koMVBtcCY65SgqlPCEo4ZUXxhylPTtwb5Xn8AiguRqYf8BON
t+4dHyq17vGtZv64HegWLPlHtF9HLNILrvXakubDfiIOFHXnevzjHFuER9pCNpW7LdSuxaF0jJC8
Oz7gDTsPNH+AOjCW4cAUZ/D4L6tQOO6/RchSObTDtoo4c9JDwcVck1zQTMsNuWKX0rg/nBCPUycA
ApRK9isnM3GNx7JSqe9qESeUln99JvxmLsW29up5JLcFtBoRPSswahDvCo9x9z51PLHx2XkSsBoq
3TwuHXJPgeY2knnRA3CB0Z7xEBpyBevkUja+6Glkkxt60KZYd5thBfNLmfRrvXFIrYnoTH3W1dzy
aXcdwMeQm+ShtY7n3yJaRRIVELZj/QYjRswi6Rlsvzq+NwfUJFumFd6y3T5W4PUPjBwJHxspqxtu
cR6ogYq/vOa3OUvDQ1a3UALrDtpRfj8Otq8qCKg9j56vpDaE24iFkoLOf9cOqyTEn4G1Y2JAyri+
DWLlyJ1mpd6S4QbgnWC2krrzK0L5IdAEFOvihPImw3qGNW7wknm6OkPEmUiWx89FFWWocdZqV/tH
LKNlR8H/L80JT7vUxUFC+/xBwfPt6Nw0eoGhP2J5OojikNtwfk5JdNWSHRe9mcIx7dl8VKcIpr8Z
16dHdq6jXhTKUHdYgI8h/6mXaJCBrSJDaF18Dj3eMqIJ/vBNsDTd/X2wioTWDSykC72t8RvVN/xe
wjDBdZ88lCsljOpj8X13RkHELzGYfRdFpAJfac35/XrwX8gAOOrAlupt28adyjH2UWjdbrdOpqWM
0Ke1X1rRT7ycOfgDy1f55WdO3pGW04YGXPcjk1WYQWKfE3tq6YeCr2bkFy0evMfIocTN14vLfgOX
I2fH+rD/udcSybZA+Q3sVBLw/904vuR879/lW/l369rp3ds6Gw7KVZVpxWoRpXZpAsX89RYfLtWg
vHGEB13pt3/95EJZl6vm1h7r0UhvTR5gWzAmDlOUha8YuOQVuYnuGq/DBZ9aCsXET3sPKoBE7LAb
mkN4Z6gIG51jXgHb1JKjaD1FJDUzbns8aYDJtUSL7jrknyYqlJlS2z4phiEeOFktjCyRyfddR9sX
MGjuJnbF1Sd5Ky3Xhz6dwUWJvqLs3CJS9NRMY+ws3tZaLYz/89iJ/rAxw/zAdd6ibcHMhB2EeE0P
ugMCouP5R/IwJNB54rydE6EiONUZCmTSx6zcjV8YdpkrhW58bX/Wd19o254/RXDk54JW9/4rJqa3
2UOmHAHn4/UhCVD6/FTer04X/d7N6+EHkCKcUHYdKM8OUNGGmTHhBPMBRzsIUpQ+88KLt54ksOjy
BGWO7btDPZjBrEXaXxqA4CsiuzlGEIz9T5PSskUry6eeIOvvc/QYlRD4rKrnR25tTvTL3odg3XR2
iUIg/MXRctRrUUCTz4lqGH86lDtDq0xbcuON7FKRRVf8IeUPFcxK6msf3TLFKa2jjDt8+rrkbYNI
Fgye59EWVZIT6Rgd+Zo/HX9L1elQmgrSS5yDw/ORdXPlk8zIlxmRvT9/Fvf7H0fP4bYhM67L9KYw
Mik19NPblPFepOCek1YcNMP34w8EM+MNaSrfSdit8jmv3TcUtZ8R8VI6CI3eOvZvb8lDMmWG/YZQ
0ekTV66QjOlmNnL6sDXm8isLYGrOM/f4Aqes+LXJC7OxNm5mIYc9aS2xFnS3DlnFD3vWU0Ed+Prv
ZIu1PfqOBSGY7WLkEgrhNX+8OFyoZJC+l+etVLR0FMci7sHNT1yLdbT9gJBhrT7O+BKlfyB7L47w
1f/WKjU8w6WTKSh2XbMCwkLSRGF9vakYFsEAwgZmj//W6JAIzECHqDyWUr6mXRXzXncfC7efobsB
ifBn38b/mey9HwYOuwJ7GerzSNXlrBa41SKO3idncg92tMOvlu964uf8u83AMsnXaz7ohVV1S4fb
uAbMEgrKqj4JJ4Nt4yjhOakjTj/33C4gUf+/h76Zrz0ooKaxGr3gj1zBUqhNY55qAFEUOyi2WclN
9bvSKXEGLGIUBBAufWJmr8Wane5mSkgLqU8SwononYIIAqoyfnasu/kOlWIf/Vze7Mxt7buoB1CX
MakAkp1zyiJjHKYEYPF3+UsZbLV7A4igUU15xURSVHWmObr4nNGGyloCok7MDn24UYBVhy17jJlf
vTf/O1VS3FERnK7HPfK/wr4HMmpzPc0i/uD9oqWvm/UcZ1b8JbM+13GV6yqlhOF8Tnno4FKalBF9
U0wMPRX3VyCusrosK0jn5bIJhFQuMNjPzuQblPM4pMeHilDDWHXDYdRhzfrAKkQemJkxslw3/3kn
3ipp80vDzhQHMw55GJZKOyLWNbOSmJImtkciSWFJdPJ2KOhgQk7A8bt6+GT5FlGOkzxcYAXqS6fU
7TkwYFa3ZAwbMK1R6AC672Rk+HVr5sm+ftT5uzfLBjfwG7atS42TIRPgD5XR1UgkQR6eNkiutKL9
pBFgmPVGnRgmGmoyWgCALXMoGyeTGg7szOEvsAFEvKG+gHycmpQAHakxlxzjIfFL+X4FWryp+h1/
jR9aEflMrQDl3CrF5P3RbLOXpXVAWF+XJ47R9haamyFHquqNW3Wysdcj8cwfNyatDcfkZDjZrcJ7
bq0nC8TPwJv5K877uoy3L0AFj7qZj0G+qdqAoMi6HR75zoWyXSFhmXMkkpVfH4vQDL3EVw9lJq+l
hal68t02TFVAbA5uH3Wf4e45kTQq8YQC26SxTkibcoXdU88GJYiHHOjmX9gRvBN4GDS507dPt/EA
JaovGeyfv0VLSGTTSxP5PYvH8ak9uyNqctI/a0UEpzxQ+xn3ldlO0HNLIu3eMvqwbuaA9glYZyil
QOiAc9udF6bt1iCOyGvwZgyfDwKSjK7HLysQWvwIyJ06Ay11MPKzLOCRnThToBGIQEA3tQUcKti4
+TpP3mYu72R5uJeePTrUafEo1XUXuSbeTkiiCoZeuR39htzc2yVh54dKvTkXtCh+KUXVDF9wfzSc
94ZF+21nO6ekcIvAqQp+GaxcNPFkNMJz4MPRNSxGnarb7ulWClsyOoRQgZdzlxyzFfaCZXNIHgPQ
57dPTPpZXCshRj69TyOkLOzT92Auwp7VKoywkkBmgtqRmQlvnjvNY8lIfyhDo4lIof2sPzWTlbFF
wd0Ro+zQKStdy6CfyuQ686R0W7t2Sd3so7nazrMD7TU6/seliCHVI73tptjmrEhUJ2XtYpTGkh1A
F0I+uF13u4BfMRtYlxM4E3Ow1eQpP+xm1fho+BZr33gWsm1ttAZH9hG/9xCGbQDI03O4DPXHdK3B
e/PAUnwor67FRLkMt5esA8dWQ4xOJOeArQQ7hH1vfQpqjM3YaMjxE5KbeYAixT3Sqy7gQQkHx1sL
6EoR0vAHBculx1VdlMRkH20xT8VkIVUk7NEpyahk69V9+O/aY9B/seJK8hVnB484vMqB4ac2ho4H
1pqwlnPfEDIyxiqh8c7kjwwIcg0QrlcmpLn4lmxQSmIH5eJWwlrBzPAS4/+J4jOvCOd0k9k+GQGq
oIhUULIZEYuTjNYrTgBcR1bkb/aXRuX9J0rc7LgpZBZLNvW0+VKXbO5QRutQAWmR7ORq2LpBf1n+
x7nB5hlxp6KXjMsh7+6dzWUtW1jQityNWsuNBkj8JLzC4SF0K60KZX+H8am+0l7dMaYx3jXzyylq
pnIVwvPB5PYrzJ4GPLvxqCQIuwEuq8n0iKbudGg2+z3fxsaj1CqvIocRPrJw0zz4WJcLx8IPx43U
a0kgUjG35Q1e5azlIyxJxdqBjvSup4kjJ1dIAZuhAPB+MrHGjnQvcz285FU5SSskfUfUsUK+h72V
zVM0b1x4LS6AyOQ4eT7bo2KUOdgd6oZUMtCJmU/Z7h/d3itVLD3r1hHtqATZvkHIcTVtr33fGpaw
U58S9qy/7MLTpaTf4udA7hdsYojdcddz0qGSHH7b3FcuRGB83Ku0rMO2+XoxO86cTxhTrDtVNwx1
ddlmakmXJbUYon/jJNq4+6oi2m56T/8CL7QksDoTSKvsgHP+o2si8U8dXvLFwep6vNLXpxN5InIX
wmUkRYABrpaIb3k86s+kVKyoA32/6fzIqrIwPuk70OdJ3dx6INbOCQJ+Vz2DliXQHKqD7D8hNx91
1aLnK2gps2YSdPtJRpp1/ofnSfGYcTg4tJyu2w+bv54Dl1R2XxKBvQ2anpqVPG+zJQpcGKwBSyx8
nExiN56w2gT3NnsQl6roKXe0epsKCZ9l4BfEfea+FZu+inG/5/gSApSV6i74CZ1W8KMaOIlqhocx
8O0SVaeAYGHvWN9D0ecOT8KYE4VvNxDIcGP20jahI5IOemshypzH7IiMqJFqIjhhXfDrPnJFSYlw
ixwEDuhZS35RqYkj/Epmz2K829POvTRWBSyvhkOWFoq6SewOn5o00NKLmMA6qV84Phu1CPhCf8PB
2sWgnm90UaeVhi7t8Mvp8Be/MdJeL0lIF0SfH6/wRJG7SCkozzLYIEe/8URjPR9YSxgv0XuMh8Ne
4F4z+ORfww1+a+iS+0GzmyAdQAcoKNuuvCZ1s6ptGt6kGR81/NbgUk5raDCyE3UpjgbbnU+MUkbM
9wQ+ituhG51VfRUp0OY1ecANYPS4cXnF71Nw8p9gThjL+YkFHCyt/3Drwm1PQT+VMXLjj6g9j22c
vgv7m33Vg6DBm2VkNjc9P+U+ProbmfMcMfWTfjHGuuB005+D4Rptjx8W+Vf/pAMVjqyNIBoKnjB9
HO9EkUoOUEqm3e9KYhxuF6OK2AUTzbTWVNnUTJw03hxWEAATgnptgw7/hGYK4TYC9gb4xSNdp7FM
ndT3oEUyai+zRaLUDWWabH3cihTVzQ56Txpp647F5wPlHPnm0BRLL/SlO7PydSkg0l6SISvntSHD
q/rJOycZRBSZRpSn8yYIkRP+Dt2t94FfhFZm9f8l1A6uKVNHnvFhXakANspN98ZmPg6ZhjlEryHR
dPUixHSTyu2DjGL/vTkOB3I34iR9H3uYADAA6kTN00TST39WOAyFnuazQ9hHyef5gXrJnxgFY0fU
83+S97E3WryEWWN8l6HmkD/KMsv/xz+S3KpRR7fVF6YrY9suJ2Y0r5vGeyY5YYq1DOil9U3tx6Rv
+CxiDAslneOwvKpUC9B7mDo1VGkPh9gWzNHx8TCIbPBm1ZKX+5ceXUGsXwIPyB2TljMzlw4PYppn
qRvbpV06DICQVjcaPPTznU8nBWZST7qqNPZQo/Xonr9oC+/UrpcMbitJV7wYEiNdnWi/HtUEIxWy
pvdfGig7pTLt6wkDcWcUjM4vAGG/QhgksZxieSK9zS8ID7PLI6wviRopT9pGDMbj8mthSXUbGiFo
SRQJm+bqnVcuhGqYzJdKfOULD3Zwjl7Utsz1rLgEXN4IMJ9qua7uowENU3NhLob6isK2dgmD3Vev
KHlHk7YtASEyctQuQZTPKzg/KSIBPNRIlfU9n4PdFsa2XjAtk3+RdfJOCbU92ly1jHIfMMD+MeE9
64qoaH4IGN2BojvG5A67QjUmVH7AclRznE2uR1+cvFlPP80dsiimLrJ/uSIFEBFQ3D/2g7MWg6TQ
X1vHTQQaQJjuF2pwQHOYgUCWbzB0veeND4kMydSYv/BB349SEVxDgzCtjCs2vImRoeAznZWb52GZ
n+3z4h6TBG6HQMFeNUfHC0/B93+Y4F8bBMlMlIIfj2y9CB+5fD4oW6sl+wZD5oNb4Gr95Vj7a7X9
4C/WusA9MM+tg7SmJX6jCecw0F+A07WLfYkZ9U/PKmsUb4gWImnk6bYUZDeJkjWNOljgKZjQfDrG
e+VnxeEgLo6dniq8vN8nApp3C4NCg3A1HWEnay8wBjcvAnSHLEcRgFKiggwz2GuzDtlu6ZTVlK8w
L3KI+QX1pTHGS/pRvx6memM3DBuVVTLs5o3ZJ50rbEyd98GQeq/EWhFQ9FMNpkr3QJibT4V5dA1E
vF1X278CIsLaeatna66r3FLNZ/94eY/b9kzjKPn0MknHkirQUQORBTtfP9dGp+v4ci6ezQECAzGJ
IAxiAbEVUTdYTv4RTf55O4V/NV8PPkX7rBPpoFpnClYwwtLrmaqWSYKYBuyFfmXuq4jvFhH5sPLj
5x13QlkD5MRLgLR0JIST7V2c1YqnchmuloKT2PFQPVj/ykKK67PIyNFB8NTefZMnqUKUXTrR9g69
0Bm/2G5DjtD+oJNu2EeW9doDpwRBZ/iIkPJU01h6+AB2knoIyCNwOIRXL/HGLbw5gyr+yGg0fp2+
HKL2sBypUfDnmvlcrz+k3vxaGAM+r8NEXOcSx4I3Cw/dJuH3yjHzcVzKG+IeIIhQjl4Txm0kUJ6d
XTysaxSDyLqLOsdqGJVc+23YieeASOu8p3XgiTu0mqyHXOB7VTkYiKBjelrKKrjCIxwT3qN4CsQz
H6+rDauBoRBduDXZQRoAFYzy5DaXRx/ifzcZkJ29LMHG8gOUbwmg49HaqEqI6E4VtyyT50VqvsQ4
CdOKg106hPGiOwtn029Wan0Mak50hBnYNeTidD9uAJkq6zLHQ+rQyIpToCUsDmbVAMOAnLvPcRDN
4b29o+n/G8atWvmaediQzS3sXLeg4hIbWo+yQe/ciyDVx5R3bGXxw+fs2Ulf6iV/GT8g94IlLHzD
cZLsNgwBHKer2wUz1m4BOFiv2OOZUY3mfGO8RIqCr3s38S/3LzkNPD8wKof8NvosPNi4X5S78REz
99jlSU5ZVXwt0NoxDHbSEMoROIHsp8YIfsSP60Qq2D5FPZ6D/3SAR5BbWfdbTmAqa59fpOe20CRO
MajpYlpTCDXuHcOeRCg1gfrIuUhBXq5kxYhPzwMMx/j2n6rFoJhIUWZv7wy5b1OOvZQf7VtPu3hI
3E6hSt2jLpOLVtbejJr+7Ts0zmkZ0oQc/wtaytRz0d+cL2fH+Wx+JTB5aKYTMwfx6HNlq35hvdA3
0ir+nR1gaSnJPisYVo6kkDS0YIXIMFwe814olkjeVzBGgDLFlrrg+cXKvl9cR54vp/1T3SBYRqll
x6XmVerPxH1lrM8+F1TI/V3wW54wzoKCuc2V09lGXXnzFKEBsDk/BCt6yPvob+4ur5xf2idGBRe3
lWFaJEU26VsBRaN7M39KV+AQAae1tW6g/CNhlBHYnZOGKIKfw0r64Ze7kZm6plZcfcXp10YewhIs
bzt6Ebz904U6nNxGQN7vRtFPo0TeEYy5wobn4Do69HmUTCdF8QQLrcUbXMOyT1fPtPhBiArBU0ZG
FEV0dDbswIHxXhmbVFIJKX22lwkoRsZygBwY9G/Gj/or71KCGTYDHbLDpj9Sh3sChvzSLe2PS+2t
Yl/XVkujBB97kWct2mtP4nXoV9d9cdt1Lv7JauxdoKzq0Tr9TNKuD7k6bd6T/pCo7cW7GIqQXG+3
wtKwnF/u5kiQlLyaccivIjW7VkYjX54NvOttkcvw/GYFXRsbI8i+fdo55PtRFIB6pA/xrmCu9XRY
yJMghq8FYy+NK7BKP8PGaHX2c9rEM5XmbGaMZ+1rZXzuOiG/l8XSkbw5sF61OA4AmQcUpblSsyVM
5xjNd9wiIPxHI3AyGTiYwC2gnLdnNLlzL51NCIgNocuyMstx+Y3iZhxNPHYkHTRnN98HthWEYbaA
drIBqG+EEDCfohrUCDZCv7ptNFlL1Eya7ACqRwZ0iMTNLHqd7HqgnWLA+HI1/UwgGT/fyyznT0gk
YhsGpdS5zLOssO5pEHeYHRXHeAN+LDJTUQ21Z+QUt/9SdfLUsthHEFFdXT81kWX0SnHCA2ooRmPQ
NK1A3pO1/4gymGROwt5Bv8EUTiWre1D6Wp7/8U4FeDU8ALfcizzgVXnUkX4I1ACbR/vckJ//ewTY
hKwudmg54LqMP0MHdGdJEAhOoliMeuhnr0nFenmhBG7zkWJAHjbxgcjdgwBpqyrCcw3uWm6j/Ghp
JQGZkEmYWCWjcxmTjnDuX/fVA6eUMqTtB0MLO5ESIbiE8p+6TwKWULMp+Zvsj1ztVKgBNJqTNtD5
o4Tja96fEkicpn2h1CvVp/yPUz/kLpegaT0gPt71Ef4QSICjjMesOCYFtRCKg0JBPS/zXxXuEAHP
sQSji4CFPgxT9iTN8bCM2I2NT1Sgtg/Fn5B7knt0zy0R9tn+c4J8cB+8A7sUuzyUGeAQRd1tMx8o
MVw27QLCTLxLt8X23drY6kdEDwKXdz0TcR0MdNfEX/ecjevPRuvBns9alhBDVxidjz3EFv6BRqiW
MKoCcB8Pr7Yn+dNxah9qUQ9C9Wl1iSv83FCb0fc0A4yEvTOVpfT6Ih4m3BtoHN9jfqf9UAlwyUZL
FBK87VGmS+zlcyiHIZ+16u+CVb4YpEzPUrRPCARS8BOplhtevJ2kU00VvIEkjO92r/14sgRiv3DN
oEOqnddCcGlnklZWzhT40AwnuIOcukfMASAdYmlDqPcUD1qqBxhaluluwLQAkF0Zg6TIQSFHeSb5
Hwcl76YRsNklfPa3kWPnKOm0x0ZqF2c2INO7f6/agyrWIWA16vBrZ7HCE0SozTc+KBcUIK3otuHP
TebiNXLjbGiHZ/1wkorfuaQbwD7yK5W+D80gsNCBm/qysuqGKXwxi8C1/OVZzrn4VHfscg/DjFW8
ODOdACCnIu7Rvuu4P7tSOTjGanGDwiCMkZhuisX0+uzXguusnUEemzW0Ofcj3vsWt6ATHu8snWOA
uAfGMXPpRdeOmbdhZneHnp+UIeP9Wo2tg8VnHRG5CCxA7G16wdw0oYwhUQQjXLg8fo02fWKtUEt2
nR+1gFTgT2SnP+nTk/FzEaG4CvCYpr9M788cvrMhcTBfPpCcq+CSF2SMXuqwFVFg4yx1XMefuA6Q
WO3wvRKDjdLvRjFzia/RJxOxm5hY7aNLgwi4x2BBUAX8ajFESQtH28rP8feQO/4w3XnbbW0ZRNxo
LKpxj+ZwZ1ANs96zBkI1NQ1nef2gNLaBEBCIoYgK3sgAjJtDlxsutCvsuVPxOFvTr6x6Eb6h0Ewr
HtMsKzpordXH/RFatwwx24g/3tnOJsQBGqUTbxVBumticieF9MpBYz3+shpCvESW5SWkkFLWta30
o13uh3h0pqKz+9Z2JF4/Vw5i734YBWcoKO1dMoj/cNzaHyjSxEaYuLsE4bg85TO3D3SQiXCJmgGP
1WMXYOGbz9ExN4rJsoTUZn+Edhlba8VgpfM5HQeha/v+0ptMll9gm53pvKTWnHRMSTGs6xJfitkd
td3+pKgmaII81g7qVzrAQpAjRC3VgGNSJgKREkiKP2u6kAAqoOs7DfqX5XFDZ3E0T0mFslqeBZ0E
bMYrWdGn4+wsB20vqy/2VR2rvoGmliKZY4SXbR9UQn4KDWqvr/7Z0egNUWlEVPfIqXj8uU/28NQV
wbFUyQ7N6yptsg7ofSH6pK1rKzFiqfuJyRt/gsOvsOHkaUf0OPQ/djzIT06vEUfn9jcLeQKQS++3
BRkqFWqaszFn2U5KCrf7IZQFO2AUA4Sqyo2VVE3AS4+xwU4Q/wQTNGiPGvZ1VyGSpF1FpAEwQQ0r
+If8VQRGdBFOvlXG6tvovkj8MNsPzfnIfBy+HOmfuZpo27LJ5Pqo051ahOByAwwLJ1K9ussi8QAM
NhKmQ7mJB9Wjw57ls9neQsqEYd0QYhMh6oINMKyzS/rV0f30XpxhEhQCr3UqhVWwnIqQ17dEDa/E
hn2NN/H+zEh1mMNb6zwwf0A340fq6vrE7uWs04UBx5Quz02m17lBGoTPtCwc7jXRSoPMRrNByOto
BeLkpgLW6dtQfGPNdTo/jrUP9qPNpJf0t0VPndcOg9GH/sSJBj8LVz2dElBnvukyysuDYzEjcYbX
6j0Ae9DYmlmBCdA2fWqZo0RzwRJ0ko0iCcPDaLNFx56n34hzaaDbBmKcPt/gD6bQ8sgKSibtvFVF
dzNUDg+zm5khjV37ACvJAw0j9+31LpVTUL9M9TTqUMF406Vhknf7uK7oyqD+S6Gg6THCBmzrGhKr
d4nE91JJ3NBhyNirmPWVeMktIx+6PzikoIRo6zsgrY/tn175gCb1Bgl+sdQslQBlIBjg+TpTbmrx
aNMDMqKAOfZKRuVODxLpL5SIli4a1wffbKEqs+TdBswF12Thj3+1D6b1Z4+IYJtPEaKXaL3Ib4gF
P9Chycg0srAFRLuzUrt8MU2DtBEF9Q9UUmOm8KhD9FoiQZTIvQckWp2rz6k7ceey1BoUKb1zBk0t
HKXR0CQq0os9yq5ZQvoTQVK3B41wMtZwQphX48SF9ymFKZgd+l93NudX0jHt6SIx3a8vOSQzqop1
LAHq4wtwtSMomg3UFOhMu3r+rzdwBo3+dCWta0EgjuD31AE/M1sT2YNmtwVztv2FV7S8HSTYjgHt
PTJHL5S/R7/Ns358s10m2xXLs8SZCGeTNl+qHLonLEGCfI7X19Zyk8u+hAWViMFrz0X5885NOMgS
gHvqYdlAuX8C5sHGQKOwYC+Be2V+PhTxDrsfY2bBAgtNm2ctbjf/sjqFbUxFhowOeTYBEzdFYrWU
iD+2jbsSaJUhlO3jI9SptFH/hnzhYL8ljIy4SOHkpWtUeYAakNQtz4FbWz/aXd9A89kBW0ErtCl3
LzlmLi/TuohRumKLDcl6taRX815yO+jqtKpR2ZMCEJoBNjbiZoCalLu50XrRUcnlXnuGEe5J1Y0a
cpjNHTUvCBuu5wKIGk9SxzF5M/zf4xzZm+4fkKNzIItkcy2v/5HJrF+p7nqQlM5E4xhfh9j7Owjd
arMAxRahVc/bgaE8UQ0aGtdfarPfrRtwwTXo6TUAyKKFs2IiQ+9cFfV/KQUdVWzIXCideOXth/hB
k5D7ttoDdxR3/7NDtMiT+jBELOH+YBjKOqi67evGoXMgOFUvVDwhAzW2EC1fWRII1JjON5bVE4Ao
cdnyvONKCxPA0urBT8Qy8ZCBZ19jSUY5aU5Rz8ZLYNPM8hepCOK3FLWtvTLjicJYLg4d7aQkEAGl
cQqrXaleZdJDMZPR6THYTtUB4IGFOeTZ3odnCe+kzYISCbNAaMgGvbPgyv/7RJWoUIuPV5eausue
FeqVB8eFvZOxTmlzttTKawqY7tJNQRenUlbxYZBtuzsljYU8cS9W25nF93/T3AQ7ZgbFMV146RjO
+yZGGpPT6GxnovgYvVHw2XD5StTfxLBT1rgFtNRjoOPuXlHBz95+iN7CbgQmPnQRB+Xg2fUKrtRm
KmRl0dtXK6MQiogeblFCNm4Vf6oUoriW4RMoRTHdH5EQOAd6tv79n9tuCVFl3Oh4/mqmi1onTJwt
XrMsGQQ9J7H7w2eBeATTXWTzeyzOT7XLInvWUm8YDbWt2sDSiJx0r0B7jcFg2NUEguwHgyJP7cfl
L6ZaHX0dUiBdvg4MQc+eBM/X0w0v9CAN5n7yPTktc7VM6WCFh/mQeUvKYijBJGl73+Q/tA5Xms1N
gIycbbX6rFXjKkKdFghNTBm4HMcSovTB1fIOmikbYb791iMbsShB8FxLLeKxW+NFSHNqeH3QnJVe
VM8mxlW/oMCYwJjBl5cUT0DvV+2pYpTErOa++vHZyrtqkKkK42nF8KB2+gKypW5yVI1ZfMiOs20c
HKylE95DOdN+0OGYZm4ox5mF2MoIgAh5zfya7aqiNt0iPCFHokmR5OsftgCmV4Ii8YjLNhxTNWfV
/KzLZmkJeg1deKpzzgMZfRlc+N4pOyF+VTrCNZRzHrna21/pwBSOJl7Q253CzwtZJ+DTjqfHa17b
KtMz4rvwyJgNOXl1m/GDOZUTmZmzKa+fjJqpW6i+CnQ9nuz9GrEmVYxN9MkXh+eacHAByz+8p0za
thLVRA9lr+r2qVByKExP0pM1yOA1zffknR0HrKCcS/bKTUW3WqThzE69MI6/X1YfNRJHyZnIXWAu
E5kMar3gPYrGGoMCE/6KmmZSqHEXBT6I7f7S0ItgnuSxdl3tX+2XmSV74O10tamtsWJoZGwsiTLS
pHVMl9Fre/h57DidP4hitrIQCxOJP4Tm0H4r/WOrIOHM5I2huWYq4hlTqXv7G9JyVevmbY4Kte//
wYE1HwO0Go9+471Pap/e8x7auLwaxOhgLsutXQ4bVZFCzleVWxUM+3m5+rXpAP0QMrQWMuweKHA7
xQPj8jefAwc2+dI10+9iNjdGefUUhAXsmY/1wAa3shVx60Dg9Wrlg7Jhqh5hcWk3NMfSlwU5QeG2
jKVOtDmETAZ3XGqnNHfLNYanGcisloYRANDZicKckZd6CbzFaFUBMatNYQxo7G1dEGtHkbcfUAzv
7pG6gyaEZtPTz7u6yvceITlD7OxB8/slzD8szb2v1YU7z4j5rXeeGuT7kSAK1U/yzMx4WNE4Hv/G
qb0HdaJC6Mqz8iEEhs9Wl9n1WMHBhFkxYkiNf1jc8qusyEuOHlBoT1ROcX8IpQk1jzmTvqu6/IEF
O/6XZstVH4iitRQVkeSvY3Rywf1HfSBDRUDsn5omLBhgukJ2oPD/zuHE/iOPhE4lPK/908x7wmlh
VQyrkD9pEEcSk5c3fVFQUlygvcgkkFrNH6MJkaVdkDdPc9Qo1Fn8U4TD6jHg27m6+75aK6cOnLfE
SIQzJ9ti2P1hDp5bKum5QFdArny+z1LkVGYYxZJRwzu1kL4Ko9y/xLrBemBoKM56peOm+jCWC2/P
UE/AGtN921aM3G8sxEcIhMGFXxReXv3Ic55mzzAwbahupIHKLJd45uocGz+YvT+Vxikfs2O/D6Qs
mdthjbAtaucRxuBSQuQ3V8aN3NyyyCgJs49dA5FvZnhloCzUE0FSEDAp9sBYJ/Zniefm6V5SWfO1
NPBpY5y4xBLqh56t9bb6RiFhx4FkGqaidASSaRyov9pr8s5X7TbcOu9vacNuVrhkonYoJyxp3l9+
qCCEqyGYRxTDOZNJ3LGlTnpBuvk16IPCfTX+r1L5abu4nqq7K+ArsamAnxXTfh6HdJejd0tztk8q
0oMvgt1T1A0M6elp2pZ2U39SZFFOnlV2EaIMyecXw+4tT/c+FzW823+9Ue3BnKcJu/nfHI5nLdjd
0JRWKJtT15XtwpXD9IuZ7k8VQT3MdyBlWk2Xayfubpy9/G1sgB9ekLiDSwcSWk/uDvCqvDBP9PzR
y66JzRltBPVqFopEzh/x0bcAvuHGXMyxr+LjsJYokXrCQS4vRXRsqwEctcs4mfOZW0HRDiPStXbt
AdK5F9UN4pQqBm+4TrUS21VQ+j/gXXfZFRo8Nf398dKs226IMbs/OiLhoCVcE3RPQQ4wzRoumCEm
bfzWzb3w+lhK5LNLPgvrP3/SWPAE30xcRS1K0jjsVDCbgr/SgOdIT/xnS3WTlHYfjmd6HbwHWp28
zCUq5z47adikst/Col2sx8IyS3Hv3TXiDCqkddxqdOzUCJ7ghyH8mKKWcAM1St2XeZgy3NC+3cs5
e7f1BfWSuDSgNMoI/3+VBwBaIARYUVT8UxG5nB/9OFhzZwYCWQ6uKvDFI0VFCAcNCdhcl6MRXwvN
xUNuyQLDa5YC59iODdCLXcE2ddeKhD0PCiTRKtHX6JzC3wdoXQgCZ4pHhVO6srwJTU5WETiWwz3x
BtdfQyvvgatJ9VOsqkkIe/sMHMM0rbkJpmVv6HHfufFiIjuLt8tkPIl+xndrfx/k/14obKDWco1u
ieELzmt6tsXQXF0eQlUeokA69ESaymxNpJLdULi+QztxTuuVGcK3QwSeYRb1r9ndVAjtQGyc83QZ
nEt+5c3sDTa6VEeYAUpxk7LkkNzT+WmRLEgyvQWcCwI860+BpHCJ97AEkw1XV4twQvSgrxybW2zV
2Lv0Apjl825/uJVk+eJguf/RPfw7cQK4UlLDLTE4aOY/vAgq+4TwSw9DfPwwTvUEWa8VC3TtAvD+
0Kc0K3iwYZ9dsFcQ0ty7LUHBR9lWsW22wKu8wcUaBaEi7TmP3a49F0KfXQlrslyqW2mk2isBMe84
96avUrQ7wZF+VpLm9yNb6q63VrOw5ikIVcmuWsimqVnQxA5D7fOfdLseW+0BZXH7r43aS0WlP8SM
xYa+RF4CzLTKEFLPLpFuGvQZlknLwsefXkN7iVnoOUy7fFryfi7m/DEjMGoL5Z3EOvxgPCYEHtQQ
g2WmJmG7quwzRpkLAvZZ1kZDkmAf+BnPyH7v64XtC+vuAghxBctstDHm72zMeGidZxgsDH82AqTz
2i8HSZX3sM17KQbfc2BUnTh7yQuiFCZyf5nixX5gso1mxDj4e/acOgl/DWGxKABbGW+sYTBsNwcL
/evg5jQl+Bqafjop6w8gcElGS/MimuOj9Mk6d6MKOKY6jZvH0OttC7tQOvYJO0iMvKTcU6LASzwq
DC76J+sbyRxotkaKyrNRZlkgoFAg8b9OLfGHrkzZkCMHgisUdAEd3QuPBBQk/a5vf6AfaQd4rsLd
i/dLWlCqjMUkBN1uuyY6h3GTk5n+1Kcdy81dZUSYyZiZ5eLGWEfq1lKRmK9U7w3NUlcpKcmbzzag
egwfH3F6MTGbF+Y2K16Q+KYCPZmubmCHcRxIbfUeCqQkvFCCGSmHZpoR+9QhyfUKmyGTN7ORluK7
jPRL01YlUi3RX4prqyG7z193FB7XnldBI6tiJf8EtHqSChKx5bbYjrcHhSbIKZPpOkU8fJLFPOg4
NlUeqLnM+DRt4s7M9hSa+2QnlmsEqO444h1QXk8bjX6XXJS8rgF9uFMXZ5I3M2OCvFFIvY30D9GB
wHRfe6MwK+WcmNIbOn5l9csuXaMILeOBfb6pcelGIVMz0dKIgzhCyXBCHDZkSTHfLv9rQr1t6uvJ
n65SO7qh9nArUfRuxAucQdlewp7M98ujmza+aLv/pMYF7ut2KbLqK501T40RmPR/Ybr9JipxI91Q
LqxFBa8GaL38JnCyjCWBY3T8Yhgz/TGMjs2vEca57Ciznd4OfeE0y8ZrnjGtuRD2aic2TrkiaoJv
wICHjpl6X+1ibTkuyue8ia8K8re1sgYE0giKBKeHUrdlIYvdSnKs2ZEGdb63ivYzqMVb0/xBwWoa
VD4lUjH1SzDGaCTuGFnV3453z4j0VXiVBLu1m9QqcvaxMF6xXIlwUpvfadpBTWTKt9nbWyDrxb+I
O0IvKdIIuhRS8F+TjKA1KFYqwU0i+01ACykankTyk5jIcyLHzo1q7vH9SizzHR7lSZMM93MOUO4Y
+o/D/n0T4v9+7Ults4j4/LkbanMC+TnW8KH5PiOmYpZhYZX0ZijG8ig95N8k+6JfIIQfqQzwBX32
i61IA1yz+B93jSwQX6iewU32MER/bZKQ8Tswuuu1b87u4srnmObzQgccZEKbTXwDe48+B9yCXK6N
MI0M5C06T+wLs1zn6TmWN2NFsbur7aO6Swrj4tNijUo684LDqBuO8HAZcrX8BknyMmqcsqruK7+a
OJfSkLZjRe9cgaCcFhda/nh7+B67l+oW4ri+0yl3oRkZpi2fE/2/1nS2D6mxSB1emF5puvsZhCfW
9yJW/5Q5X47zY/2sq7oc1d+ukflkOgznQCwkIZBlVNn0Nj2hUbrzqc4Qss48KK2DIf6znqg00Cuc
ns/Px8aVCxqtvX8hlEKAw6T0wkTehwfdMfUpGljpAqWNJIZqdQnrjy2BQ7CMH0vaqFBdinkfpA0n
fICSh/BDNHt4PfPYzs6vD60Wf4IPJ6n0szyyIrSj7Yq1WJdU9mK0Gy0dn3rThQPcSGiMH6u8ENcP
7w8iV1mO6Gz2g6yAFY8N3eLlCEJm/mgBuZOoYskIncWF1VZewoW2/8b/MzDdPNj5Bx4sRe+US/y0
vxTc2OMYYnB3PR/sBAy1ZJd4OoRC4iXZGIpP+4mQhEtLyiSkALyRWBu45clhV63KjA2mxL1ID59q
63MDWTFMurLQ8IJFad1OjPmFZ/ih0Pnd454C2s/FafVzpWDeaHfKit8Pgls6BZO5UScEBYca27AM
J0OAAgs6QV2aWeUFc6A0t8UJmM2rf8wGgb4FE6AOwAxvUlr+gi1gLEuNEOvdoJvu8qOw16fsswH+
hVbtYXHMP/hxGWqk3ahN15mdApcYkudp4HgRqA7YW3jzl6nBLfDhH5hjsNcFpxerjGc3H7MSv24r
lLddCdOMTOdx0+f4tG8tTR197ajZPdBVviKfllzM2QVOloUCF0/c1n5BcVUduVH/qp4SiVib4rCR
I01IoExLHODn4nh1hVbG2fqLmC8ffwbSpp1VrqKNwN67DwEt9eBbRq0TiYHs2aY4QjBkZ8qrJmUV
0Uw5ge3pgpDtuVhuyn57URXXWrgHo2vCdP1JrLDyQLF7yhbCwpSt4cycv0rFTjJTm1yskyxnjip6
En1Vb7vJNY7MvZShw0A140/CsKs1XZ1My0TSuWAO72hF+6PEVbzcqrWKJu8h4f4dZdA/RVf2ExA0
Qy/BJH/KfFvvdbn6S/Wvw1qnYYfDouT7nxhB2dPqPab+/HwrU0Mt0JMbJ688VWkzJkQl88frvb/s
cOd7EDuErevLMZ9p+zllMMemmzZNz/lM6ObAUlWy5xxQ2/C7+KLSNbWoYnaYQqa5CTzDWmZPoFpd
GyvTzBIHN9kkoYOWLmQHnerTbI7d0ZselxqkkPAH42LDxiMDuYPpDGY8syXIkm7+riFwnDc8iw2x
Ga7dY07Ca4x9OINTefOY96lQtJzMcTJT7YCj2KVDntFlbfJyEILj9943awhGruv/qKBarUlK0wAL
KLntD9/NWRFreZbXftzdlX4eK/brNbZxw6ywtaIRlR4WNJ9Su8ZmC3om/0KDwAVEV+2onXVk6aLY
etiN2c5KCoW7+oZhh9VbODwbvNfKbj3BWM3sSoAy/WfR3vX+8exN0LHAlhOfGa4Uq3aPM//p+Rq4
pZ9IFIvgaf9TzYoNYRANdQKuBcT62nFz4hw3z+JV+uWNLZZaVsjntI+cW1oC0ihyrH5IZS1p0NFV
orfLLkaKOGYzVZWdhkyy8HfDnhYL/V5Zj+cqOUJq9d8m8wmpgcGT8ERWgvs1WsZyImso3U1KtHc4
RDoCy0haKrFx6NU094ZWCv3VTI3dS+K+nYXfgSfpUoG/y4O5rftUSP+cLijUtxVBxz8S+wAdZkNT
6CutoyUrpCWRHM0pGbTh2vhL4taqXr4l6SvHcqRrSVIbMHItVpK0Dc0OvT7B7npX/YPd8azyoTXQ
GIp4sqEcFkqY8FZxEwGXJYaS8Mo1N4vR9pKP71jinDDc20HuxWiprANZMZHXk5zIW0wud7ozBJbR
Rgx9i9lRmRBygzkqUHs8KNXwf0QViu1fYQJxMAj10lcpkAWPyNOSkwBNhN7xYJ9KvzTw7nFwCua7
KWMvKaw6JhsvGAekg9de1aYn8D4o9jNFNt1xYam3hMMRpAJd3SIOxZPkkZsyCfwYEwkmrAKFF3sq
CjwAMlL2PXO5vBT2XlCH60bHnY8QY3/vSuOHZlBgvoP+xjKqcHUIOvdfunvPmU+ON+GVzt5dqamP
LJVhyiuGTvezq6DHMYnjqHlqoQpStMFeEwzz+ezoQX7F+y18+JGlxR79XAgRQJOIAQpb8O3H5hyM
bgmsMsrAyBl0jfJgujEN5hpkywSAXCnu42Od3mOJJ7Yar8JC6mkrIJwrAcTDjwWK10G/yDCTHhZ4
Uc3rFVXJURpVctgG3arbp5tMxoALJFUAO1xKGfFCNBbPzKcJRApM2Ow1kLbKNXZTSmZhH4HoRA5I
n6yh/jrUfFMtMbYshf9CJm5bmsETBM1iUfMs2nGq/17yd4QXjRePdKRHGLTIScgqvRgw7d9gavh4
HSZrBGiw5yyN7k6lAyijuQyTQoAhTKeL809pniWLYfYODTeqM4gzJbvNhdiXpHLKpSdHyh3NetXD
a7QLzsTWAJ2zYMYjkyb6DT4KBOsEVVtzRFzIXUIJeHevu1q2peaaVjq4cHIxRLp4un27VI+LHogn
ng8o3G99Eoueda6XENuALaFYFFZ84BD/H+Et41OaVaZPIDNZMvllWHDJhrNX4Pj+U8qqlizi8mRY
5Pi9q5jxhBPX3JnLMSwco0ijK8/HgtkNl0ksN10loTXYY7y/L0irTpWL4Mj3QV+D19+0HrQnruYB
TRLj6MHUfRJS4VoukH66ykYTTM3gUFr8ODwzE3HsSrUkKc66nG57CM7pXNV2XwjoL2VlBzIVAppj
pj87R/hRhS1KuMp6J97TQFqCbKSTQPYy4+69/vtZ5/y2fsDR7ubREeBVLPl/x0Q+XY3BZWJt/BEx
MCOByKfmbN+n4P2hZhv+wuGCx8X0Q0D6ljaS0fZ5tnuVILgBOCbMwPUzX1q6MMZr8zOFwUqZItuX
rzwc0rF3WgqmfwG8Jv+UKN2ega+qHqgvYjPaS1qJjNpQNFREVDgHy9T4WXX/GjFVMA6mRqSrH52Y
Fv+OwyAp67MM1BMEJbdLZtWRWqkar+TXJ0eigtMSy68Cnq103it9JHxkkOQXI4VdZ1j3cKE7DiDl
TlpzCvGrivxIQhQ5o+vFeUGcDsYqqdwdCtK4aStdct8fuk/NGcid8uMzcMPatMs7uHjpxjWdvTRA
Y24WSXh35Dw9XDmehT4YO88P9M/cyfORlzHiXM7UUNrTskag6NQ4kwsqJaVjVCfDdwPo3TNfIote
M7vge1yFeJAdnki2IUfXMBRcwVPeDhKmFfCZac+QKeFzTwQp5C5Drj0AlYJ4ntRrB0aLwC/QY1Qq
rrgE7zrMVZzlEGS9pRBXazS6bVbiVkHIQiTw3W9jS8LWUJLkIhdZd3tXPGsIY7y1eqMLlc4LRUU3
EEcnGgMrFrjjcB1FStighQQrTyTaVV7qwcWVKQwiibiENAUDRIWr0HYuNhilaVK9OMoQKa5nogxY
4O0sQN73jSuEUJ0l6Jh3zBtRI/UbZt2gud4PRe5UIyia1q92LAEik0gJjpc3hrEcVSqaBrBu8LYm
t0PJos37XRE1DoM44CPszXLtrdeN0lJq1THB1zD2z/MLf5RJCZGeaqH2Y7PboxDALSRFck8Kv8Yy
19fjTkQ7o5ryHewSBd5dkZbx8GglvzC26SRxqKXU10dLBuoV05+JAwfYa63mdT4E8NnRGWqnb2ir
MKudbKDcGXriJMgZoHyKUZiPMHHRw4eAcT8hXpVFoD40/UmyQTcXJ8e44GMY0LzH1P3xLlB20ToZ
eX2BVuPsKceMaRqJXkfTYWxw+EeveUFZSMpmJpoiSF13+1rDVzBeLByo2CCHDp5eFbo9jr0QtnQ6
ssBVXp8j89EdgM0/RIwSWJXf7Enn2JOag5YpZzKFlCdLNnTqFxaXO7RHDqGX8bgI16r+5ANHGLZC
GX78Rqpi1Kxe+IgGIqOodZOe2ucD47AXoKfwkpOov8ovmDknyyW5O40SibmnoA8fmAJ16A74ztzy
w3WyHC0ENKsrr3JFTpSr33fLNBZM0usOWI2MQVal6l5JyH4LnF8tYGMBJFo0RTwEm3nLuuRhOGIZ
q5t+nlw1pMo5vXk5lec1sHyMVLIrRVJyHLP6pdwewgpSpFbkzN93ePlgxGBb2Ci2IRefqD0lNf/4
/0mVDJkZ1bg7Lb4v+T73ltoPc8SKBxTVS+qeM3I0xWLuk12Ss+8nAjE6NQov23YZR0un96NOR4vH
c1WbBHY+eAz0MT1eOfHHCr36S0vwxic//zw4RfJXF4gpW/7NjaEBqW3J1Ei1pTc3BHZvBapuEzXk
UuFGpEGBR4e3343B3+Kun57MT74ISt4dxROsa9UWaO9WPUd60sllIO+y8q3dn6AVV1zuA3mrC/us
NYrB9i4nVrsml200FT4KG3je1WjBJw5oiEJaAvmVIuTLA9WlWkKtdPi+qxUT+riZt7gPv6eKkpIW
MRCuw6yHtw98puSibAxpcwxNB4hX1UekB31STvEddrpSdrB7zvxo7iVKvyIasCJGiEfa8wSRUDLR
LvBdNkWZdlxQ0r/LjJfglG8afNX1ACBa2tRIoqyupdllQDGyo4OZx4ZL5kIJxYpQTzVHvvo0pcBg
LFmdbUZlX6W04ExyrATBFjfQEEKa6iePUXG2yQ11+Rjw3VIHTaClYdc0lK93AXaP3UpjBzMXXaIT
9MuPB1lz+XWYrmB9M7N7DKYwQxcKn2you069d/vq37ZBjljmk7NkPPx6SZ6zJ4RZT75oTFZLqpv+
+5uHrdlclCBiKIZrsP8ADVVq4GajzYxSM8MXmoY+viK+XvF2oI/i31ZMb3HHk/UVKBdYprgowdvJ
sAMCpKEG5JLhWN2v09R8Lu/756J9ccHMZ5sPlh1RKTUbdFAT5rQ5WjAUJ/tA/k2/DM8LQh6QAkIG
UAJuU6X+aq2kqCD0XkJLs/FO4+BvqB7zOMPiOn8cfTEWmnGHnZvDrL118eVPoy7ws6ciBMtr5yzW
gXnI7TqVyiTRbM4B1TsIlkaxsxWA3Xb8VbxnfMDWHAsQPoSuGaxyAc0JMitAO5ax/kcXwMeiEqqt
+isoLnxwe+f9AHIdGC1xamQWvBkDemIrgMl45f6YpGgT4Eb2jIlVxlUAf9mP5i+VODKeRpgWrZ5K
m/IUEUyE9k4CEsvLmYaaV69XYnqTmdLyVuy4uMq6TJGSZGJvST1IARLo3j/bIONUCO4Nfdb5hmgg
0+mEhk144uWjRWgdj2Gq3NobjpI+0THBkbZb7neFWKPzSY0ux9KxKbRYdERCKkMHC+fkVo1SGfkP
/fq5+C9BMXyHDefpUBl6+bxYGoAydQ9JjDAP9x2adMWSYef+cpTTMZaRHCyhL9S11OmW8XoDFYU7
+fh7Z/rw/fKUnZVKVt7C6F3EbHrQI2G6x2Cg+F+6+W0ksTUPkymnlEbE6hw+/tr4QlJPzelAqFiQ
yZq20004UccYYnEneIEe/yJgGDXadT5KbIRkIdI0DNnhmXa7Yf1Mcfdh7OgQib/KYc/2f/WLlJfF
WF4KXWMus4ymLwmMnAorkBYN0/wHcgsF8ZhHCtSYk4MbcDg730mfPBtIq+MhaRoQiAX7yIuLC4Cv
sT6jtoYgelKe+0dyl41vIorpS4gb3vdD6zL8goetkDs2U7KnB/q9VH9dtguCCT1tD1b3vgG0vRHo
mc2YSBsfEF+6wJ69WCjndE7BPVnfM/aH7K/cw5mOyz/WLS/XRgsmgm+du12aN2YFxENVRS6lQtFd
OZAKOAvW1icYHmumVJLSqUeoE3J+NiMRT6H6QCbwKMA9ly1bfODPDNu7BO67No5e3biTSZXprV8J
RxmZ3vhxrn818H/2fx/lgeHudjSovrTgfPwnLdiDE1HExRu+wIhBXZGkFgJSTX9n4KYChO4Tu+w+
8MIIhkabtvtPXh49rCXng/46COz8Vp++U0i6vGyQtGLsTtoZxj4ay5+D3gBjzlq6wmb3M+1gpJzc
9eGEyXwvl2uWfrjvAq4gLfeGr1/cvB8HgwMUeVtSXVVLmBxk1Sn/JR/SmLizhw7hKuxHGfY+KDls
6JWmpIxVVg4C+L14209Xf4hJ6Pjp8DLMxdyW96XxAxkHdqWzTNRTxf4+zOINJ6IZBYEgXWqHI5fe
5fYJSQx6zGdCF6b5eeJ1sQS6InW/0hO8Mkf7SEE/MzSZslJsNl9amfWrAgUHNo8/8FFIBlWuGVfU
naVaOmPjdRaL9ehKZQM0fhHerY/MI8VoMscyj8Bb9Ob2HPyzbMRDcLmTbsOkahcCHAAma9ofDdeo
Nc/FzCtQZBmVD9CYgcmQ/1ijZC7mDNAlyqAkJnvT0Gy+H5lq3zCF4V7wqwx+AgpQUnqnyrU+He7s
kghEef5SonUKc/E3i7/P+ezeEafU0vN9LsBnxEN3KJsZjGiUY9u8rXIM3WVH/ulNuf7LWVXe3gnm
IAucezSelUquodzZPBJF2ABC62nDq3JDQJLiMoejoq2q+kHeYYclQ7LN0FFot/FVeHwNw81M0Rop
+QeB8BpmxBpwcO1funnbIV+HteWChvRBvcz5EIqy3vz7+esT+WABY4UK6/BypFWrf2jnxEz40ylf
l4l0RaEC4gwHXzTmehX8JGHge0tvY7BDTp8P1SR7W1ENfG7ayqs0jZkSDPvV+BQNp256QUxODI1z
0AZ9iwJXzJEW0pEGNgGatbuy0++ph6iXIjaQwQ/hszuuyiJIowFbyvQaYMyjuJEHDExmgbX0GjsY
S67q4vIFzO1I8xShINYvLQxwAz75RxbXj3O3IYnzVm3Pq8QJDsBOdyj4u246ylcB0S7gZU9hS4bO
lZHM9DW3FaLCrg2wE1jV24h/vHz6NMHgSESqxbK51/orgKmRCe7THfsKUC3Lc75/oG2jrDg0bnPI
43//7g8hoP03fhn5cx3SFnJLLsxvW5RbDhd/w2WEGgCvoKfMq0LJeDs2XU+/mVQ+iWyPXQFrI7Vo
wTPfbREHbApHCSc1CUlqp2byIedeVuwgWHKY49kVShVpAFg3KZmm1QHBvm7nD71sprNDLV6Ca9ch
qgRYng1bS4nMyWQY03O/+e63Q6MnO7MtyjOEnizPMcSRKR6BZPdJTvt9yktlcx37fBIA6lxD/EiD
BbmUpUzlYcF/7jKUtIdUeAlUQAS5dX8mmVpEVz5ITEg6PledXi705mKmUrwczGdbXxwOYQvHAFzQ
t7qwFQY/7cr7zYrPWao0MAa8J1umG+6XUsYpQgh3/1Ug6hqnkKVPjl2/Rz9kIuaFXTmjob+uGSCv
jeng2qxh5SB+rndzGxP3FbIpn1pB8m5qM3WXky1mSeITipmsM9mHq2MwAdRxX+yHB7poFRNQ10xf
0YtknxKeAwsNU/DMRRDj8Pol/VQbFqCQZp/AF064CJpzb9fopJutZWBdI+xQIWiUUevM1S+zYNTe
2mu7C24dGv3sf34oke5cTDiFTrrLimG2fNUroAixmsrcGjNc9ZsvshueXLIjuDlVEbd6V3Zus9/U
24r3iei4Imfr+u8uzTibjt5J3F0+os50vrdYljBPs216A561MB6ZQ/nLMoqirIqcB1+k6MlhMU4N
h1SMU5vpryxbpb8vvK9PHdIBZPcEr9d6PZZQHdbWtmAenlWYHerrEzzVeLcrXUas/VngvRCVWs1Y
yrZ4QMKIXai07IjinSmDwwo8MllRxIUdnU6X65xcRVnVC/rrzgB7UJb3q8liR0xPpCnyrVQY7gQN
VaM6t7kmenI2lp1SUWmjQMds2mjqUg8O/dKfwAO3K9zH0ojoqf308T3WsRX+Lz0wIPX0xeWoPg0P
8WhB6xa+wKSssSooQXhH9+AqoOUVzRX+bYkblWJhUiyfppo5gj+8W2GDVaJtN2PRqbZa4R71ymrP
hqlzRsu9F330USKS5lZ7JphmaxOwJUp9O7sNa4ib24jDbujvdcbTmgdm1L9cAHVUcUL+kokfcH4y
+xNVWJj3Q8tVlyC0WpoZdsJmM4s9W0mDmY303BPYXw6j2ilEeoRJ6DMl2JmjezkZxl/Ih5Mw4lVq
h6xCltOfLtW+mN6ZPwKxgmk6vchkfz+jJo8kxh+pwMs6o9KXhTp4lBMUcDF2Q/GcaWo0bCicRXgH
x3GRADvGoicDBTy40ejVepssny/KYCy+zkqQtXf9rRXp1EagZyD/p+8dt0RQu6tajUEZUc/1Cos9
Mmb0On4DW7pm97brEw4rJH4cQksnMsmXVKR0o9JU3fXCOiEf9c3btg2G02CZ2Y9m7AqBi/uoLcq+
eWpi4pZFnhdDZs+tEnvXHQ0gDUVrDsaiItoAHOtVmyutcx9prtSMhn03Dt/mMNe51tQGeMOcT8p3
jFbhv2EVjbRlzUx+UY14Y4IVndOYTShO8leyugVmyU3UJAwNaDmHM745iwIMMrwOkwj8zhK60cBK
5NOSy1MvkEVr3lXK7FyTIvf0bR4oOnt/kA/SnRpxs2o57jJE/C5Ue3Dj89/70nc4UWX5KIrzVUPp
BJTesje9x0gdr0z0/XcSnTVUis+K12gvUVQlggfsl81xdbv/jWw2wr95ZDGmw6s7aqDjWXHJQTGR
3il9cSMFB9OZOOIuaLlU0EoIfyJ3LG/JhklBv322G9IYpzrWyz3mX/xKzw/ZLCj339WkwiGSvSOW
Wk2lKrjZCzlYaOC97g1NZWWzmXzBRCq+jjpTtrrSez1c90VwaRe3HDTq56o4SKeuJmUxlZpTyzpq
G55HusfCqKjLrpxH4PRZ56mY3rEFxwpSSuxcq5tCFJ+dQglF8ZY9D5QPa9rizl3mu7Ixb/jFyF96
q7oTFwrYpyJ6V9mSOmdGg9fsm+MzsCKLPrsEovbIUcdZcIQ3XG0vpUqiYVdIfqQ3oqSIloUmngEf
svT20Pgn+0KFl2q+/fh+fMhK1JUT+BVEoL5toxGHjI0E3+xYW9PLOYnO1MNS2K64UGasvAnCFR/1
Lhld8Z3Lp8pDZyGOlWeI+BI1E+f7DQI9YfGELapwZCHmuoQ3nhASahHmeScPpqENYtQ2SNZELwmY
y+ApSEkKsNW3EG0lz5VxWfeRUj8zBil2ZN8fpCODRVW8NJW/w5ErtnosiXiJ44UiUT3JwXfuoSYd
SuqTHGGPDRqArHE9FqZa31xiD8NUw0NguDVeej7RrDVfvG4sLJ+yQQoCIhmR3A5oMdVGDVHwAH0/
vewmhOHIhhtJMmr1q792xE6si2bkZ5C23LjTt20+UkhETnRW4f6v2PRq/oE8EjXGUImL0kN3HBIc
+/LvLK51WBt0yCHJAkpjUrYFBP48hdYeHL2v62FMlT1BPgGh1w2V575zhRYgmB/HFqIsBsrOiUJs
CTjvpNVgeGsW9Ro9Y97/bV2PzPL2IVhdqdzEQqXcqeqmfca+vIdCuHNufHEx3pXJtDdBhpWTcm9J
Ur4n0zM7jwe+nbbCLA00w38bWb16n4u7AoORjieStKItHOOG5iz7ZiBR4HSXJiL/SpJQykna75Ty
6Chq2PlqCzcwH3splQ00NLfd728sWcGv/BGnge2ixMxL186AruSSPI9sb/e3ErqGXn9Pc5uvevx1
1LRsaRQNgR9avKFb0V7mhN8o65jHkEt+koDn9FgEW/omj8mX2H/BtX/DCBDgu25swap1TtLpGFPP
X2qAe0Xo1fABIbOCP3MqIerVneJZnz9X8oIKrgZ+7TXJ4srEdeSniu8MAdCb8TidodqWKQ2Dps0V
TfUSf/3JNu6MHDc1nU9Exs9ZSyDpSnHzlDhj6SL3j2bRhTz01gq1jGVLBfAo0qO49vCUXg/u7/2o
T99cBwPrk6ioLBiw8RdhsFsL8BMtrydZJiGm0loxJhv8QqwhcYHGc7l2XOFPlRc0JyEywa1P9wDo
8z5RVDVXcjZyJ8R5khWtjPxCyP1a2iCJ2hpNEsQOqPR+sgo6ZVwEqIZwq/C0BbWdB+ATFBoOYHqH
GaV47JpMBmeLMG+akNEx/4/LRy97tZ+5AQw0Dtjf0yaf85bJq23aXDUZDv1YtgOEA7S6nRStgBTh
ZaC3sntvOxNJ2XwtWVC/3AyDNGNWkMVTXD84XBwEk7CSZwEWMQc1lwn8FWEbt54W5nrwrNtIl0rN
Tihn+OkJan3leYobqv8sryKlYHkq0rM4GVOReHkF6Xmaezm06UGYXKQ6Etg22DnazUfzluA2YFzd
r/9dgWcus/s2OrWSMXw/lw6nKC8yLSZnmqQUV9RDKq4UKKNE+TNW17NXwM1+DjVWgqE4mvhOhlwV
REiIHQbm6cmLrd8xxiLkHz9MIj9sVDbkL7zgUqHeZTiIcBJ6kVHi93ml2kdwvcmomXjk4n36eXey
H19k10f18RwXsPywwaXU3b4PxRhHv0n5pqH8Gg7Q8N7VqjRmzX88PiFpd8T0drHciC60jLrKhkUL
ujxcXsTAUKgBzkZ+cNgqOxnwV1ebQQJbpHIWktdd4+HNO/X/jJgK6D2NDuUdQ8VIIBQsGxYuqBF3
IoE+97PGwSwSseh7ju2V49rtyRPt7sd/xASHlnUKfuvN233S/UfupqO+mgIOzGqPua7l9St1fipO
RNN4ou3ClTnqK+KotwL3YS2CxCO0lQnfA4MIu97ZzdLRi1hMpm9DaCsQzMXWlqfNmRdptlJ81pDK
MG+kA81baL2Nix/8xdQaarJ1VrgJ4y4czwcrVpXWCWbdV6b/+06x6aLJqA3TZv7qVl+HSUnYnCZi
xnC3vYgLlP1ogKuOPV4Qu7R/Xocu+UXmz2TtaIbsOgi+eLCvmobpUB0ABp5GEaGT50hVb4KYi+LL
MpZk24YQDffnNJV1XYR2VmpKo54epiz+NbyOE+nM8NJob3qx2ShoNu2ETiKK34MHJ9slbah28jHy
lhr6Z5v6xxOuiNL9qkAYEC5rEgdVmhtC5HluzlBgsigwB1ZBYUPreets9OSlODbuauFeDUlonhG/
Jzax3XQNlRS3FnPSHfIOR6c3KSrFdUc7I4BA6RCj+xuOo1Y1DinblQPUY2dmAUxHcVCcn9g9uLd7
kCR2qVJ0DU2xtJPSd5R4ACXcAnnsyKKvKQwHNiJw239uP3WRJ/z46UHpPQFBZI9mixDMznb5BlZa
dp5o35LBpm/zOMNFkxhtQioRQ51B8rPHAByR80lUGlYESCOsF64w1Yh6UEZMDhmWXcTx42eRx17O
fNoYm7YvTPr03LAJUcHnWlNDywJ6v+1pIiMMuUNn3o9lpekXmRGkxUV2KPk8CizUbDzunDEH3Rln
rTBdQGvENUjGrQuLpreQJBM4dmbaKzmGeedoAaiUCQt5p33uAMzzYd4QEnxLwP48ryjKP+GrYEfL
nInBLReNaNgC0smgn7Bz9/XtkbUAEQSggOeAOOmGp8ui0oN+UhBrLaYeHd9tOFEnsy6/X2cFPkvR
VmFvF7i5knsTv4RzcJ+HMH2Fex4wWD+onR4HID982/2U7EFpwI80RgARvyqnvXJFFsiPwPBko/Jj
4GDrCnnIo7GZBoSPP77bScSHREK4HUAlbYkSB2TkPrp6VXKeqEpipolc2iF3D5pivfgf7wS9X1ZN
R/ZHVsnR8oYNZdAkAfeJd3MCNE/sn0+o6nX243Dep1LhitxgT7KTPwcCpl+6gyGRINV93pHP7BPw
lfJ9QUh9Z5yJ02t29Kv+5Lh5+WC1ecsNyf5myOpNiQzGbmcGU1FGxbqb/mfDQlpOnsQQxbeZjonK
083qX/vf+i5PLOE+AQnzRNHF/P9L3uxfqleVCGlIQCeLB59ryKgou7HF6AdHVAb6PB3IC/uRIvu/
R59cKyVuED4AlJ/UKkfAK3fOuCE22GyW/nOJdvoUrFfIKSNeinbUnkQONR1JX+Kb0hyY57jmVFuU
uir6jLHQoxKQaXm/uAC/NsgG+/fIfOVXdYK25FwK2uuE1OgXmGN5ZKLSaTPzDuPu4MCr++wLK254
N3q3etVIgpYdw6v85u47kY1E/+jxsii47Nz15wrFkzwW4BZbrJ+rwbfdiW1gNIc4rhT5YL1gVlHg
AU8RQ1FjcZDO9EW7ZsA02DgOU2aBUtKWnrNUMKmhX2lBEnzF/ntJ4IBqmZywS2ZYXvHiqpfyKHpu
tP/trYHbXu7I5A78eWdgjfjZSaUTFQUCtqCyqJQF1Lo/32l0JiQAoLsxiDAYkk5tBmQWagZUAPL0
XtQZfF8gx8Nk0o+zmAZFiSzlHTawT4+LY5Eys6nHknk5v//Wy/dvYQfJzG3xv5PZfk+FMj3fAtZj
YWNDv+LO6xKjooWMYFbxEtH3t+XhIuWXoLILPu5hkw5iUBobbxmnqoQxJ/G2joFjR3aABw+Z1Dww
P8MOddUP8zUxaJHGomkeWc3x4nlNcsdIX3114y5ehxHq3itO6JYv/FRQZqGAUysFtzaQqdWI71PR
f7/iWv0oCdSwqhkFPkPgUZanFpM5XNP8tu5EC5Zka1jnJ6rB6tTZNdoSsIEOjp3LcFxmrguacQGy
e7jjWz1rFkOUDrNEoFxnH52CpXTqLrF48PuloFhhSNzSWcGAZEofODC6sOil0k0dc7pM1nONsPB1
vNf3iwhCtJlzf4EKtuiZyGPi3Kv8nNIQXN7hoWJukQ62aVO6ZpSM7scrv6X9FCZ+wJRPinMYp9Gc
ABFPSPQ6NfRC5KzU5zcnI2EV08IpTAXa0u1Pv46Axha0AXt17d4r0844a9sbi8Lo8e6wIInNpqwb
TCQWXJ0axgBceTFv+8Xpyz7NuiklVzLoklbEy3Ef/p9Nd4Tn0JbrPuW4FURVHggHxX4aw6ltfjoi
yZhwvhdxNWiRMFRTm/99D0AJyCEawWigopr9dRCAz2i2za1edTz8xKKorIbj1H42A8Mzn4qrf0ls
NVJowBOcM/kdAMrt5LNzAyJPMK0v6Y9Vel8zd0+UON4YzKYoT50mkuu9Rlq5j3ikYORDZsP6abYL
zlIR5bq+/dzDqlCJDDwwJMNgaw6ScQOWJrhTpDhYa1QoLvROivytVH4A/GAPqC/qe1T30hzsOppT
OVuRUGNEt4ScNgWKk0/BBe/OSV0WMnG5XRI5GewmGDDC70RldBnX0X56taabMVBxa1fMT8HuiRKq
hQH0Jjsw2OoBXmbS66QO4XPwjL78DtXgVZNbxNoXEs2tovsu6bpjstzwkVrIT2gWduKy7JkaP8sI
Au5SRY2HT6ASF/AhEEiJdPeQ+IG8N19KwFmVWHPbYdrqSv5WfcurnEQ8JDHEtEUFSVP45QfPeOF9
RW5j4gt+SEnhbroa11RCCl/zmWaGrMGmY2gLMxLMvy7OXYmdgFKQOQx7+YPEOOejn4pLxOHnDzdU
J0QE6iuRyvrZPiwgfFS4HJzZyhpPd1Oxpsu7Euq/PcJ5pAz58fjkA+z1CT+Vhwu/5RwFMEEQ+zF/
+XPfoPZYFGpiSHBKvZlhrB2zbnOrvWd88glxDdkeSUbO41rCRI7np/yyMBzVg5nKKOQrmtu92TLh
q94swlOf68DJxddnqRRjj32G49OOCTyy3Kssf5Au4e/iwZPVPl5z9tubb1sm1UarBNYz4kQ4gBYE
9bwXhGKNbPXRApJPNl9XBaUpDb+Yv+f8//wW0eVuZN7jDaX+3ooFsbpLxVQ3SNHCyDjl6Kkj6v3F
cjJgAbJcDeRDjrKQ36aiWal2os4F1cmfzyJIB748+ZMW7MbbPb9jNGr9l1ss3YIZGuDxh4SZ2TKL
/W4opo+BD9Yk2aeSh7CqAxqSAbW7C4449fcGj06crtxRKzMGwCzASL44iQwMrZIrUkNsNeFN5RYS
yNGjedSf8FiJHmw1LUmNXdI04r4U2ub4nV1h4007qveJi+JEvEQqMA9HVT2lkuzfsyWR/x9vJoC/
rBvSAkbuLvk0RIhBA9VZUYoR6Up6K6+HKg2ASx0cLH9GQifD+uUW41kvDAaUVb+Ydvd3FDI7CGnP
fYGXcf4GFbF/aioaZd6ZknTIpNMN8+3SPUMzkYnDrrjS9myxGOapa7ygMGCtLGBed1RR0wVgs2Ix
iX++5JzN1OhQDyjuV7ymZSWAJbDp9RfpU8W3fBqXgw+rTLpTdOLRvdeMl2v0+tiUuOU8KhFdgXif
uKKZpfX8lv8pr9Sukj6PoOatB5cnKwKwAIlqFzU3ClIWR6doXQXCX3DsoFuV+nqcQQ9ljfwUNECp
tuI+b8aAs8GBlA+cyQgyxIJpH9/GrtsrYpGH0NXn6WZ0OY4vOZyXP/EVHFN53h5M66EIhiZk2Vs1
SSA6PuZa/QtK4LaLMxymHh6ejyu+enj764e5ziNkCJn4VSSzrjznDtdveFX/8oBH9l0MbF7ebZTF
4Uo9HW03fxXCvgI+ILydMaV3LEa/lfc8MNvvDLlQ2BkqNCwTWn170YxEvhx4FMmAB3gkCV91Ea4N
S6Z99yDFVT+LrUhLehV+e5Ga7pbDW1M/nd0MPx41HsP/+KsD69cAHBns6rZOTNzjkNvOz5QIgyrm
BpyrTgfHAktLP2TeYEVWinBoF1Fs+91NZAUwooHdUNpZthRSgimOcO6jGdWENGY6Q0uYoiFv98qi
hKU+Egz+u3c0ifW3A2yDaelHuVuvzNuEcxePdQibdVKB5PrJ+8bCNwzHOI7Q29GfjRiYobg5PWRP
lARBQSaRqLDMYy3mwuygpIz343uVqhFim2m5XvKH3AV9jBsPWbCMGMKBBvZIlAMkHO6S0qr5jd7g
UWgbfqsz2FppAf/Rz25Zk/hPmpQTzXr/CWBP7GjjBMSwMr5UACSYNUpQUNU+JmAFpIymtKwf7v6E
zsXn5UivVcoj9usd+2zSJlcHMHDBFRMI6txCnqmqFaN3m2cotgTkvBE5n1ZNws48hpIbGgAbLbwD
yYlWQUsagn39J4wPPiKycuy6VRTujq9ncIipkxNRKlnO6f9Mtj3po/fpiNeqym49Fc0VLM1mCRA8
nCPq3XNRW4gpNgqKBIdTi7LBUdtsM5PfYeqrSPnNNtsXOMRfp8Od2IvrQseOvhg1kCWHZyb4jFfg
/tdlVhSWPIA0z8d2yEFCD6rPJH+BEqHivCLKUnT757+KY2IUARg5s0DhpQ3Kt/5d1vzlkcMf1VGJ
5SF6uttojXkBi/dYs97qxFTCLqeqUE+ITKfgmcGiDLpHLHtKqzIZmPPy6Av/SxNvnmQh1PTSm0es
0rr5Utmd0S3oJVU2XdwJipyoo4S33ND9xC4i5MUxCbFt3DN4QZ66fDuC4zbYUkcApdHc3phmfEGq
NnAjEhfxvK/OudBioS5EoMQXu+3nPRQakzmwT+Z4S2uBuoQCgBL/rHi0RURXoKFc7e3/UTVoV8Ze
+QOmTyKjaKfLMjB6EjCm242TvoYb07FYjfbebRCh+0tpJ/HXXITcrc1shuRIbXTwpWEREpdR3i3N
DEK/kYuojcNYyoP17qOun20CBERBbb/6uGVC624C3lzcLtz8/T7gdytmLx4I6F+s/LL/YIlwTfnd
naXCwJz3xgxgt/4Jw9z6O1cWDIRgKOBjrQdZt/a57iBBge1w1P97s/Tp3mY0CclRlKAOovLTGNJr
zwSPDd+SFsEJhy8ComnT58QzCMqqfYdk7orCuUM8S/s4FZM7WRPrh5BerPVgqEwRs5r0h3xTE8kO
yc29K+2eWluL1F6lAGN3PYPwEb49LvQHpzDVfnMJoGMKznxdTyk7h92Ks7OyXJIqt3QHwxzKymVe
d9fcRVar6uWyV8ZK3GNNbhV0Xb8AHJI6EA4etuqwbxDmccvYzx4ZsMifPEOEr2IDb1v/bx+FvNzW
Rm4KuvKIb/FjLbFjCbeADYVGXYw3NBQuup6OngNF3Z5gRgsFRAWdaWVGD3+gbY6CoyMkcDkLPhrK
WSSc210AQuooFRMi4YqTetl3umF4rFZpRz8EEZgkql6IL1yKmxKghv/bLXcpLJDIcTT+/v2Sjmx3
wdTJt5zDuhholw2ip8OypgUdH3yWKY4mDwlNgk5wNUW7Sq+QFsS7y7O8QRcpEy/SmvCsa3P30ual
IFrL00qtx1xwLxRcqyUZ5h8iYiSD8kQjlDUCHYiu7ziJlc3ajbnhwvvRubDQ+xSJbslMst9xX0Vd
EUZQLPJyfI3c3rgCbG1/3t1wgYX0Q+sdjFyTHYkU+7LTuqrsAXfiub4TmSUcLdMfJ9CTnP55mTp6
k96kT0ouRJe7IZMyIoNtI4LKpzjmHCkDVDc2oQdUdq4HNJedP8pIBDb9MwmNveTBxl5b3bcAvNQK
NjXIaksuwyawDiU5x7y/bPnN2/HG7Jg8bwlr/4uMhk/pOVCSOFMBM5k+OPHz6wq72qY28HTL5xNl
8gA1u/gbX1TNoBYHI9YCvidlMzG+kKU9XBCD6RDQ8OSPCGUsC7zIhwUz3Cy/BielGIxit73b+/KQ
QTisBifAUFXJ0ijDw79jwPjdV4vI1ufaD6SokBKgtRMmQNvf2L+hogQ0SLJaqAeDC2Bg5/NSkSMU
l8O5Xb6EgGm+iotavN8G2W1r+enXGMQCnnryhKCKK6ioHkMHuEe1b3wgFu9VxBywFWD1FB6CrJtx
g0sV7VcnsYgBS0fKEmXaKFj2lpxazYW+vjfTT+rAndvDboDYY3s66qzO8ON/5ms5nmgm9b0GKH7W
Y+Gmr7769PX6qgoAYAFBAeqHyTl5ARI5HZ+s2XlLh9sz6rCVprE4k/cef5z8BHqCnJUGHsCbkWWR
FQYw0XNh52OQlVrP7CFucfaQ9Kw4ctsNKzoWkMCLom8iqedEyuFqvLpFZ69zKAeqhLmJnKcB/Tz5
iz1A84d+ntaCWww1Q8/F2CTrk/caOXdH4Mvr6ofXw8DuwmRiAZhcbGFzPpRzrQmWPcOT0OmkRi5Y
KnJX92GcIgEfeMwlUBlkDhnqQnQc/3qcHe87n5v6JsQlCqtPw1USFcV5JTUC1dk5Gvy/3Us7xVrt
/XWdCDALpuxccYIC01NbOvO3CUWYV1CZVvnJu2F3xM083UHYtCB3pDXa8F8EEkn5dfWaAQPvIcL7
JOCX3lAPeUCL8XclUD8P14TG7A52MKual67zH1mrIg8s/nYezDDUjfH6s8/cNnF5lDsXYwvEOBah
JqLBttKm84Dxp5akkzXvccepKtWp7phjRfBsnS1AEaxhJC4SutBsLHBSXpuwxiC7ZsPCd/1t8+9P
QLPHp7y8p4UAtUJIuPGXwCWcUyAkcjyPMp8C57Z4hehwIEsjNXLK36ygAGPOo4rfMEVQmp4QvtBm
BAsILNLD37hcoIV1tyxI9OJDDr4cH+0wvcVYRhmYlv1DTuaEFOdCO/l+FyfbC872V7Py1gnuxsD2
7CzCEXyAzovH15hmVlj+3ncBtzvpQkHbZi+hlqUOImtPKfnCqRxgxB9tIczl0PPy/3yG+z3Heovt
6G5H+PJYKb5f8exkQe8QHmFq3uoBVrxYeBHA3vg98ZjKNgpAD5tGZavv/e55oiT/JHVXzeqg3q1D
3QH8e5WVZgwB4nGVHmuvLz5JvtUzjOVgtNYWnoZKZogyhbStoF1arMRB4E1KiWP2BSZOquS1wWz4
GX4T7kiZFdIev3XCN1HIJfoXJ0i4yvqY5ojmxl0Cl7nBrvJD7g1zjG7fGt653OYUOAmO1iwk3ljp
dUJ8MTG0LBFM0eLeASGdtsRCZu2trThzCxjwbbSX5u5mS4TbfUA1Tku7gWZADD4rXDJZch4JyFYs
Kd8IGsBp6TmUKCWAFANEK52NhzL8sh4htPlJVDdX7Bpz+HLxLYM5aYFhe4ly2y514HZ1Tg0AsEPQ
sG/BVcFUTR1Nm5Qj7bj+Keja7ILiGq3cvDpRzPk0YiEcpL7Bh5HtimsYhHszuw4h4pnx0x4hubaa
Ih7IBdHkXhZkmmDjJCm9SsqcAJyIhukzne+nIvgbWvIswNHEOMDxNPKZp+X0Ju3oDpBY9KtE0hVu
FyXF12yt2x7rsajUalWVinAbBrq9+7Atdv87ExcSMiI3v8iBFzVRQ6/IsjF9dQpD3AJyyVvIop6a
bKjo3P9jwG3fKr8KJEq/U5Tb5BDT/ef6lg3So9EoC64gSYv/NR6vMviSiSVEF9Vr2MA/D6u1oMNe
op43SWukMyk2xomM7TzL987tNZrRLvbFoOuox4RfZBnZZqCQxDYba/zGFEO1MYrxy5HIEQPazer1
nwlUOUVbtFbs1qHlayajN+Q9Hv0jml+LKLcqMnUmZoQVpjz5J/NmIu6rVF/PBAIU1kiSpZEMyOQK
ud8kxBXNmdtpKkDPTBOG8tKmedN5siNsOI7tnIJdb0KKtSeyK+YwYMmmra1dyw5dWnd4lXQnn+I5
d12E8bIZ0VGwlUM35OrwsxIhe9ZwOtVj2Snxp0qrMdSAaApYZtuRA6rIlAXqNfP1aWqm3DEiqzAd
/FaZMHAdFHFdYlM92fgQDz3J92kmQE+V/4odQsxisUfem+7SwGk2TRNcVRao6oCV4+aJZVoincx5
xH4t3IWcCjzRKE10BVn7y+gM8rK0S5i70+zHEavHTi5Eefw7pkvsISKbfRht1L5ek6wdpXsy55kB
esMe2l8wM/fyuTPe9aEVIp6/leMfMgnG0RoVwMUgT48Xv0IA/NRk5lZPlt5KN6jssoY9AvB+1bnO
xfrUAHDv0ZPrOw6jHnLWQ/fpxz+rnJOEA+SbsHO7q8Fr0wuOHi49Av5mdjW+b2mtYMKICHPFF4Wi
/NsPGk1BLn1pH1vK4rmw63WXiOdzaSbyij4p3DmuXMAuTY8rwIQAFFH5abpeeTZlcwangiSTqFZf
M2kEcNZodLbTxVLgOkBW10Ej8PCdbWTyonOZEtgafkSxqp6wfC/KQT0reJxDhAFEVdeEV9mdSj2E
cH1oT0OAyFW6lkjxgvXYxoyTUkt1H4y8EFbUD9SplywPdS/ju3uWVRr6Pqh14xNIRBDDLVkdgWAf
RU5GH1CjBFImqdqBbaBSdpvmkJe0rDj8OaJ3tPwp1BLBO/crLF7K5QYIXC7nYh0t4A7jUEncZ5G4
ST1CDUR8tWgtc93eVBKNKkGVb7EA4Dcl+PZOzLVPddPJ2uAMmduBOjpfL3BSEGIo85+AzMtWb9BX
KDVxE2h4ys2I6CfjNEEEv7UmqxMfBVXaljpd5hXYAJuV8GJYSLENDP8zZDWHKitUPYdSROa5PbY+
znPv4qKBGMYh7KOsbvfhhcdry/XAuNUeRZ9lULVqPk8YLZ2zxKyz4xTBN5A82EUxz38DFH1Cpai2
KKg5T+FfH3Hciwl6GmJP2HIMtmfPyq+bFuppFwDQDV+kS62EoBQiUgnrpwVcw6g6ybZswrqW7D5Q
fMBoz5Xre6UE8VagclAgsOlqGY5ToRA7+WRhUoesotO+yZu2pKb7jI8M7mRgejSwphF9Yt1PSSIy
HzJ/nFsxD50IB2Jm0dxQFX6zs+uoZH/xIJd4ybKADKXaC5xDRDJ1zpYn28aAOqVZt5u40SoCt0VR
wrVAw7FF+iBAdSBtb6yozWm+8P/0DRt5dkLoKaUeuiZSk949eh55CdEeuzIDl3JTFTysylJGwRnJ
PjfTsx6GJONWYyJ74fjuaw1O0PoEIbXbZgpSCAmG0DM2Plgg1NnwCCvq0uyEixqJ5SxladYffvtE
Ha5i61IVqgqoG4lCPIEPksRAlM06fjzzbJEtm+O4itX6euAKgTyu+vEl0LXeKMYZDnlY9WIDTVeP
1HoS3B3vlWYbcLxtIkKTFywZoralRgkWW0a6FpOXD7RQPKqJEaUWo2TZFFwgg1t3gPMgsxPZVV+p
KkiSs/dKKYUb7Ue+5pveoqCfnkAHX+X4CDDci0b9oVbs0mZ/JBvw2G768XTOmh4AazbzknqwtgUu
Q/eDw+y9OPQYjDdK9HcefFgeugnZlYrUGyDXd8zY6TWV+GbSHD9ptbe46sZNp3JSMdjMZluGdWWL
w3QlN6ObnbaxaiUTJQPrsA2UZLLatTDl7O7bvJ+LsjDwtYqiJonyI4B7cku47Mj7GUojDHjKByn3
TyFRLiZtAGse3Fmw8aUw5R28+6vMjjvnM2ww7TXrz0cJ06HwMOkd3QLX0cT3Up4AsMueFHTgAlaQ
p95aeAcTykNESUNg9xUlw4md8sTNT1kwkua2S2neExq4BmKrniyayTu58ChQuHMO5rtXdAN/XqMf
F85VJSAz+eT4+fg+YwsV9uCwQBKSLUTIIJ+BpX3+JJ/y4Sbhvrym0kTn9dImGUx08C/epkzEnW0c
F59zXrzFExsorc5l3YdJ4JxxUAGT3AYIADv/qBENJEKmLs6sPO5jiUQzMmbGMxFj/GV8zOBHTe8v
r37G9n9X17t3HSyLtT+B9kRfaxiwv9jE2bW8U4TsSe0Ip9/i9yaivtNbhNw356JgxjMahqV7lIgI
7HRNR1KPOwt6yAV406dhQcFDmRK0THZC86lfC4GBt9HpeZh+nqHLPtfcqx+imvo1av1XHw/233GB
1aTXJfZCbLaIB42vmmnRRPpOmY3mYg3hUr2iZL0XQy84uIcuajz587HD/mOjAV+jyCzTEVxQTkLZ
QgqkKeCy7ehQpYXlxeaK37SV1gPGTRhvhh9liDGI0xXhqn3/y44xKmrH5ehwDrtyj/O18Jdf8Fx8
4DkW0QIlM3lxEMPpuPEnmJ0J/DX4KCuFC+FOKhi1NX/ZCd4fs8ZLqcoWGi09a9bUUNbidOG0XXRJ
rRAUO9x4bdgosz5tzSaOQWxZtkLVurdV9J8L09/6FRJBKjUNDm80gIMIKhs0vgNgfzmQTbeswV6j
vOHF77ZsJ96ccqAGGSzM1+k+4mEz+z7CvESeKdweivLhzmwbzrnK/pOFTlCkPdCN+swjgh/JcaNv
YSUsydEiPcjsw21hdB1Qhmam8zooJKouavC2h8kQAKUdPsD4bt2ilTG+eVghDYblaAI/CGPea2fa
hvhygUfwI94TPyXZUlMJnzscCTF5ai8SXUGf6IuFP0WzvDnIr7OzbEw4wXraJh6+jqk9Zx9+9VHA
BI3cUjJvF3Yjv7A4peR73kVW3yqP/3obKRU79pIdF0SDjo87kczScLC7vsnlKyRL3yCdK6/PEXfF
RJhEahKbvrlYQgR6LQPrXeUFoaA78lGBJ9x/GneCcYPFJxoWGNdwKK4oYH732GIqG1hZKKv8XBKg
7sdCjOU//fg5lLP2YAdzNPi8BIf04zSSwpBFYvLg7cqtshzxSmwkxX5MwZON7pZz8xwcIesBLnQs
QbdbBWz7hy6XdgSeEhgdZD51oTQ8enlx3koALU+kQjx8cZWkIl1ni0Zgiuyd1icdkmf6swrXRRgZ
tWhkN7+L+/jzqRy0V0tF+44gvbp4OIRBWPLh/spPPF+tv8rQveNoin8EPnRXxXLtcxkLCuND8t2M
mOKS3G6gPrPpncEZGhE7Zy0Dd/5gDfpEPbWZKjFE+XI1+vGPsXuk+M4EW8XC3w6aHjP3jJb9s8f/
f6cQix8i57UTVBwJ0xI1KeIREGnUb55gdZjewmR+cot1vnQfKK43bxrSs4oQnqq3W7zisiSzu/ys
6HZbwb48KDF2Zg2LcEbMyLrRzBlv7ZXDrmlIdVNmWtS16flNi0DXwhWsFH5On0qZHZOdkmP32adG
RKecLk5brbbaKDf58dxjvuCbG7NzUrwY/2lwYzagOQHxNR1F67tXlXCACXipdNdMrF570+FYyZ2Y
0oJBE+zFsSd/J+lJlbYRqIgUwCNw6ETqqXq6FLyfZ8RsKY2Q7YLWqragQBZt1Z0twBhr8bcyOQPv
sSM66TeXWikPYg2X9coYW+IdiQV+wmpQPO6cjEUg2bDX7wndWnKY3xwkLq5jULWEh+MGmdMCJciA
GLMwaPDZOGHTKc3e5tBtiLeCNzLj9VlpE9u78jzoKoTJVT/fAuLa2XSDm/cSEc4DFR+ARHqR7IKC
bfXvUK3/MpOK4r1OaUs2SDPuujyt3F60D3k3/kUXTOEy1qbQdQ3VYY6hl4f1TZlsEbGyJjTTekdH
bF1LAmzae2Nr+rUov+2L6T0qd7LQfpA5/TXhX75xABXCBiF9Sx5vVD97eGilsYx3PSyeafYu7Xol
XxLzVAP6xEscDwP3fJkoByrlMja8weNx62odvOs+iaCGwYGpTWTwQlFKN+l6RueoYWMWIMR3OVGB
0tA7d9whymnxxYr/iALvMxQErTZA7vaM5KHjTZpo/pfg5PgYz4yTgTfjXQv4sp05soFXXgHI6fCJ
AGiutu03quIrckCrluXQC9BwYQRTkhMinZz8D7YhOcQSThh2BCqtZJZFDXMbACtLmj+R38PT2IZ1
z+7Lf7S5IPSEdssKzBqhV+UP0tYXBEhq0mdleySZN0urDmmzSo7/RTDpigjxO4IKLh4/xZdE3RtH
eqUgs6tQqJZyUupiIRkQ1WVpoxNyq5TQv8vMZjGyYP50x2mgaSDhJ2RZY9Grgxe1KUz4hgwtlgyL
+hrrtjcVxmzMpAXL5vBSaWtXrF7VfbetpeAgWNFSym2V2Nzg1m75Z0arZ/LoJsEpJsIx4nCuWJCe
d+mdQWWYZnWHdPJVSXeD8hp6YeLNZDE4NxLSo1ZzD2hL6Ovb5iMcDz4cVICEFSo7MCK7XdpzR7eh
dUaI0PXWsvzl5NBGDLY9NgmgZ2DmNBg2jG+P7Vqz8KpMZzcHLgy+6DUKKFVbt5gZEyAwIAMI9kkD
t//Md7sAt2yugL1eA676li1+feD/bxzbJtBcqHSydyRZ4uSZdikQpAg1fyz3s3WnceXjlqlGDwbw
vHjk29A0rdgs43FXXftemBznU4rt2O4TaFLRpn4fbzJGSMyLm2hVI5R+BuDs7PaJ1W7n3Qf5uvca
F41a5T6HCmaqeSfMSwgfLnQagjCD1ZdR6yfu3bXyFwPBE00//ZP85IB/4yxEPJoz6eM3p+K1RJgc
A9q4PJ9Cm5q4kz9/mg4F1cwxM8ROpHBg0XD7r1gO2hDnknUNx6zWR7NHGVtTLXQrRRCC/5t2lYyq
7TNJrvsEWgNvLqz9HcLTE5W3dXUPThvnzBE+DnxN3a7y9bnPpWB3PP+5mn6FUgvjPA4BLDMe7snD
x6gpVe6dZbgQlwc/quKEluFeck8ip6kV7102lGsrG4bht55UUx2uehTmghMWTqL1LoVLUVKcu3HX
7eqUtwKSiY40IYaNM2CWVu4NZJnBiPKery+crJJrjgHnLTfTcsIwm3yfSdg1BnySdLiKFIQ6lKH3
nJShK/Dl+X41L8vrEgF4zJUHGveUksIW5bzDo4Fha4XFceMISL0AyKR2LZMlexrR1637G8vQmoiG
kdVWHYXsH9sxytiR3+8cMZYhIKRMwwIu8IzCOc//Ssu/Qq25niwxVjZxQ5rwDnj6TEA93sm9yBIS
fMoYeY1llXgigC+9bUZVcb+yHjC14rPKuG11NwHJr5iNN5hLOgB093V72VEQbKvWrfIILEpBMJEQ
BJxQfEEukcYPBdXf9snDs1NuKab5L00Q7hTGGVrtmI+T/po48IXQYt2oa3ZakZi2/TsXDbKc9zuC
lXDhKb9OWMAW0HPyTex7bIe1gmzAGtFDmU2s7319AclApn6R0ZNYYn5BZ1yFob9Whk2wib+oRthr
LKkj73gstuKtZNuw3zb7tZENUzKSkIpluixZFU02X0z0zhaP3u+/w9dF2BeLOqo4N2FRPsNEzMjN
zH36doPPL/cGWVVhdDiOuRlv6kcjwauR5Jzskj5UPdoFyz5+klyuw0ak+SWDTOa5fUXtIjX7eXzZ
75UCEJ0YZmOMCWa2s05DCUUh98gAMDmHkXNxPay/8CAQkN97qurU/L3spBnsVzZbMKnTGo9pmEv3
fdy1IIGCqAT/c13wrsKp7MSggcSAluLPUKatKCYQO8z7HlgJKmZ6RBL0lp3preOuK2/lugUnCFVc
yPGmZ+EejYDMxYX2XYlyQkSsvJZ5+yoMemO/pXTPqM28tSij8SqrKIzRdzeIFogPatlIgQ6CLrRs
biigatYfyd13voVxc1ygpG+Lqpv1QsKXu796+/5le1Wb3JSUEDbQftbNpQjsi3+JWCsBG8F1iTPs
csBfmS5d9jE6GOy7ux+fw7bRABcXQfYzH2Y0HMWdKtRF+6ouXxvObbkbW4KaR1+mZdpx55KdWvK9
3658e2yTWbkIDr/eVbmyi6k7sKHGFtCxe1WjqwRMe48DAUFsPD8SZBcyAnHuLQFP2ETGudlAe418
0Y5VgGIML0/CnooIbOHI/jgrLG0Dbqa/WU9RCbFdBQ4UiRYfHG9Op4s4yzRfwC36xI75qgl2ji+n
abV1SLOQvCIKoH2l4MY8KjzGZMiovUJ0h5tlz5Is8LmZuJOxOstHBF6w8uWvxENFjNdEfmRJo0dV
zHqrlND//DyJDoJrLyfia3LYTi+YWC/E/XKQHKHXbOFCleDGw9Egh1c49TYetUX4b9hNatq99t3i
gW7etINrxQmyQZ0MUn33A59Kj18RIM+ygcPjJe02ANLvP9FqhzfSa1vpQzqciyAskPcAVRNZtX8j
BLwI7ybwTGsoPwR1gHm0nRHMb40Q14o8ju//7vNYBBhYNRZO3eWRog9gWvuURNYvrDS0/cz3e4Kw
rE+6VDAswKL8QwUDueT0UbdA7XRhsxRsLHE916fvCVQODBwGOONp7qoVtZGe+gTy/OuipXie5c9z
jk8RLkvkZOHohJhXYNnb6Vj/OqsxWu7P1judYZHboqg9ZPaxnqwUDECKRGsbLWTrIEsJeO/E+ZRe
JsGbmC6Rv37jr348bMHInDSuqg5GWF9BPcoIaNX3ULzEOwncU/UXHarYSN3RR5pFoA/mfBZoLZum
IkSZElEGun3HRCF3WT+zgX0Lu1fu/3d6/8BkTFM8oQ2CSUnXlt8UckNBYK0U6GdKUacotP8B9HnY
ZCF6a02qwxl3srcyVTPvrTyGjqGPaizTge9UYxHLO1BKUsk7YaQCc+TkFe5YJWBANogmdDgJmcX1
mP8Md3/4WJX6VKj1SUYVQaWtFT1WZWY+6yf9MfdpT/lDLZ0r2LIJLcCbeW/0xB/aVMQkx1I9fNBb
Fy7paLCZsEzJk8/RwD3y7bwJ0hJtsLYgWq57ymcA/dRnObLY7JLbPUjLLZIB5L9KsB2GUFAKALKr
yPW5hG30SyFLwuJPIAkAvACuNA6w5yud8hBSkaGfTjOY5ihM2QUxrTIVWYwsKiOlrZ80RghC6FcZ
byyM1zyO3gwiVNYyy2yAn30gVccJ1uWpmnXlqFhXeQudT6wSS2j8KSY331gfOzBlrhTR1u/feZqw
edlRZuo0PBLprXw7CZOM8389Uzcc99yNqV5h0z41jlcvfGKsvMPPeGK4NKj6U6QNzzyOnUt6q0Qt
gAjORaEWJdXWqkHgOzQq7BmVkVnJEKYrBIEA65xHyF1QAbYEO/68CF2LV3xnGxI4FE1lDadVse4E
sFwp57GksfOSyKHb1P7DNhNSnTzaQjZJcy+ExBZJdP+wujaRXsrJd7Dr9v1N9QdXcjEy8AHqY9nc
vuCqrLe4E1Qspe78KgUVSlNid80Xm+d2NN2u8NfzwvZDsIIg6GcWETqeGCsK9gDD+61oM0m0d/P0
zKim1P/iICTFe6umlACE4Cu9FVF2YA/FURMMpWqbCfXlXfEkbxhNRBZ9lX+5U4ebKP6mC6xE2CsI
4VZ1vEIGcj3F9x5f+XotBOeUJ0GChX+MeMLVP3Z4njST+HjGk/9Wzr71+YHjCfia6js+dpAkXCwu
OHvmjkQH+sRkJBjUKFHyzZpRneLEWM0xd6fzzzXy6Ls5gAgsIJvOqvr8bC/HQz3wOpJw4f+aFXH2
Fg2nTM5iWq40zG1b7Vrx49pCPIFP6l95YTaKryxXaTCNHBYsE7HOpwJqRAIKoEdwL381d46hq0XQ
jOluDTacSVikbgbPboimH7iyhCpp4l18edTGi2ssj7Hz19Ba7J8BerRWuce7oCAh8cUISG+JY/h5
aANlGFtvTnyu+6KfpA5AFhWnpJ3upr6pmqaNIuECMZHdv8Xfc14dK3r41xufr4N2IKmObOxamOgq
7hwPvlnRuyme/xmzcxmR6X9sGLpkBsC4Nq0UFqDjSS9vgzlGB1gimtZkN4VQu6BV6z+WcSJ49MQO
U/2mN0h5/JRGowUMUF4p8z/5cvzaAtglMhOXsCmFO5KE0ryWCrarM40XIy6J4qrMfa4rpHW8o9Cb
Ih/IO0ALW/+A7g5XJrgKPEfromf0b7NZ3l6XDoG0OuPpzthsS5keEA/T2oT/9JS9r7pbjM0nLzvh
lG9mjD0/iwwv1w5OhWGJBjkvQJrauUHAGOGTdq+rjdT3iHxMWy6fYoI2DzWatlmep2yDsj5iLjXM
Uxvl6i10GC3zprtjqR7X+E9OiuYnVa/jed1iheK2ikaGyPBE+TfVilnk+XVFAwuDE/M5P84J6+/t
6YibExDMGAxJWTQLPYRLkgdbfsmeP0xKdkgExQMUYZ4TId9rG+6Qr69GqqXmCL65VFEUWA6+evQo
k4yRucFGD3lHZ3/wj4+RvjephyKkS+CBWmzQEHs6EtEFcv3igG3xxB74j/FMYGvoLnihDADtXs4j
FetYa3D6ufh8RnBx5A+78kOSOswRpGNBktAlQWyy2LmAy5F0//tLFnBmuD8e4FBvDInbt7vszDvK
MorLhZB9YodjoqmGNyCm/WtO2xcTu2a4C/9kq+M5RGkOMyg8VXk2if7iaE9BdvuipyLaJ+bHKiBY
o0Qd9HUzRfBJicioNuViGzaPaGKiLNFg2n5XYL36TlA4cHdxpAqr/uLI6CfHytlnpWsEIulQ7C7W
E2fVxkSrysTUobz3bXwdei75ifkK+urXSW1C3FAXq8kQWxM6a2ozVWiiDJrSJnKCSnn3aMb4qv8f
Wdv2kjyPAwqpxLhvC/EGtzf1ClvnXtN+2t6IlWYgbXLXlkfSJiXDEdR9EW0b8er4ZuCHf6v8SRlf
DzAJYx80TaU77mVgPyRd1ml49gp/3lGROe/UY0/it5Sh6jOCK7xpIfvqyM4bzwJkjBqh5T/x/Dkk
DFNakzUmY0zT9/C+MfKOIacU9rFfj67E4pkG3M/LRjPfdl6BKAfeDytMKwt8UblXdV/mHZlR+W3z
7kDLHXxuFVwvi5YpAfaWhgK7d6UlzFrFSy16F1ag2F7QdAdxZCC/HoIj+NkLeeYjLKZT59x9NQVI
kNgtz4yf5cQu4X9Acust8HqjsUyu+WUl+3frtuCiuiI56mFDR/e2FlHH97zDonVZRR57aZGtu4wt
Ct4dPawzKLb7dOinEv4wzhcKd5B8ogkSYcAXjynE9WnEgsBvPxqZ9GCgzNc1/8ZxVihpOPtOxUfQ
AivySrpp7OqPLYG8kiKrFvXfVm598/NgOaf5exMF9/vXz+bOn5MOhtrXkCA1pZFOK2TZcQyDG8Vh
+3FxT31inWljesN2GoW9go+30fqR6eJen6EjbvxvKPPI380+dlxMyR1A9dSi7+b35ULl5AvK+POX
CPzaygf512Yv+aDmXk+qUWxrFM7fGgeN5XuaNGgjSDmaz+Qpbc2xuxuom/Im9/7Sb2BZut5WSobb
/zxbKT4s/ZKd5Ew2GtcQiNcbOIY6/vtznlCRVprFUstf/iRvOLG5UTU/SWxZhtA4Onk14Dv0a7yy
8MMGRIfTOYFcuq1dQOh4jl2fgCUdC8gSAX/Erfy3lZQjEj95LTtIroz0FUMwBuQ2p6mmFvDlvs7D
EHJD/GlR4TDuIKvfSYNJLsCNKd5VU5qyLkI9pdbRwnCDeYhIyKwNjagdxQ6QW3pqX0H+/zjp1lmN
qTcu6esfFQqgFZUBsPPxGFPZjpS1Drgi0jqVT7ZKpAmJ0SZyKv24/StYrrCR8tRPTcR04N5z+1AS
Gj3/WiTwdH3iOs+pW/CyrWJpaqJZwOFUq9AwQBpD8MBMtfT9V1y/sAnE6ZXbx5Yc7jn0glNFnHRz
IfH6yk5FaHX84ZUe4d7X3nHqWSlRj4148XU0nJenUKVVtKeuRAIiH4aDABqysgHYumW4QyOEyNnh
Ud7/CFgxYm5/B7PVW0psTEQqfWF5ZEX4og438U51WamG+Ji3dyJa+hQdZw/t3mcn285OGKb9E4By
xjnKMRz16KZRrW6cJ6Ut17JpitcGGEKdBQMOCufjEZOS/KzgX5Eqe3vNPJ3anrUhZuOwtu+IzgH9
VaKUmqUTCKbuxuS+Prm5JCTkgwYOzg1/rTz9JQUuGFIW2HDiFZpT9xBI1IZOhXdQXKgGQyZInHwl
ppJwdt3bAnAHwC47yM2e7puGLa23nFefMf0oOrz80k5BH4OWRiszS/0PKmxvCCqobzXqMz/dj378
teNxU1DKT3doFIGPJ367MXAfq3TJhfZLrAfZZWwTIcdXcNb7vQXADgaPoNe600Q3yBPkHqhS4D0c
tAPdAjet3ouqZrt5+nFb4S0vDWE25q+ev5YAGbN23YXr6mkpYovvHe5RqkHN4/y6pQSZ8IXHUBpU
wECOmo7Evtaj/Sw5HW88QSTmvohQLM2trOKfSwdgpyjLgGfEwTJhE8+yQShAO2eIejpbmh/H/HQ7
bHH5SatO7nC723PNWB+uSdK91IJ8QWaXbmzaWzPtC+jxwijyaaquQDphOG00ywi9HThd+7CmgPno
UZ1QbjcOQdi2Y8NdgeKcXcPslVZ/zdNkaVn/D4GrSMNXcwGBtRdzuvTRrXR9BVBKvQv2YqZuygpA
MW+mQW2YOOAudDgC9PKeohYL4l9Xhz77oMKwX9B2l/X0bmPbpdwWGkIRAtunfWTsb5W5u+mfDQzh
iDfvr8ZLKVL4NZNAuzmIlzPSqxUJJSpcmU5bD1jDNUn5I7XctL1ioIOokkxv7ewiTLSE11mbNG1W
aJxOCEFXb2WtSQzczXQ8gPcnd8MgJDpK5Zq8+bP2jA/AOLxvL7VjW6FXtSRJtXrVmQydUuVygPJq
Ojd/eD9xf0KtsN0E6Soe2JqxCNOvTL7YVnE2ELqo8x/T/M4trTRkoX78vbq/FxfT+yZgZT1zI0BF
+VHXh+/4MQB12L2unaC1dpZlWSWcjD9GN3OhHc62LBBlyDDV8st16M8UARV3uEOG1xPeQ30aIDtK
dLvXp0/QdHBQUPIbxkji21Ssa5uczsjzH2u2cQovWNyRJymfw8Ix0DZIhItlK19vJb/bTjWNBD3v
46OXQ4pTptKQTD7/DNPkYjLizWl0ZqqA9KpzF4Okb6O739/aM7fixoQQa6HaNch5FcSBjYY8VfUD
eq741W3U+H/viYKvP9raqumkmSCYBGvx1V0VDdAVki6bRS08nsvNztO8/5ynB83n4khQdLEnwRUQ
C6uww1wpfjBy0PZPrivcRVutySLVcRYAeL6oRxSlhodRxVpz3Xt/fH3wZqo9ljPKK5Y6AlscwO9J
MaYcaeJlFNW9vbNlaeysV0y7SXzUSoKvXs2Jwm4FuaJB54NEQrUKWSaUyhIT5vz6cE2WsL5ykSMc
Fvyg8tDhTBQe2u1/TFv2rRtCBO8ZWUDKqXsO+2MyuQ4nMOZtKXOabt3262lkr9ya1dbiO4s7yX1V
Bj6WgDiOmVihkNNmqL7ByB//RX4kkP5HUvF0R19PGzX8JLVmspne8oYSAq0lYxTZfQ4zjmywKsgz
8L1Gq8YVeCpaHiElphPOlrOhdL8217u1k7JCu2O/FtBkjVzo1AUlIgRFouRLonNwSq2UNo2dNvLl
B4RkcJAvZEbsrnLHZQmU6NhU2CnqnIC9aVC7XAMOSCvsQ/FqpG5y3c2MZ6JY+PaDGlc8aFyx/+HD
moG5rA/CGraw14OXjy9zi71yr0V5yp/VPNuFkH6V7y/Qrku8iD7/Mp+nxqcnoyCS1jJVYTlHEbxo
eeRHAmphz5QY5pmEBemNQYMAQdeqwq3DgnXIshX+s59vGhqTX+6yc9QdeOzOyhTkJrqYmqaJ/UBH
WhZCy+CyHv/Q4u5O9CS64We+lZyzjVCgeE8a+FLif408y5TwNn4oLVk5WCGp9wWsA8jE+rXFxxhg
Hd1lw1znzpvagAvyMSaw2Q792I8KWQKl9auVqtee+YXccZhvUiFn9bGORVo6DVi/mzVu0/c+jfmy
IZeyDAsdqDryAfuCqr8RgvAay58e6uUo1lVdRknCCO/br98EZ0+AnGRQGKETfFGuU7hqq2ZFrzwu
58VBit9Fr6mg0vumkkDiEjv+s/sMUBzbTXaoWUvp86MySVCXWu91RLbfyjqOik17f7aFUjSKWQ9n
N5gjul36jg0m+kMnpgy2G0bn18IRCndFzObaH5i1vd3Lh+c2cEnQ6EPc4nW2XnqAWRLqFX0p9Ds/
vlOd5JZ4wxzWLVDdSbCWV2sybqcxrAgS+gZxgLhZUJqKDZmhT6ND4ignqtrsG5h+HOpeugGQaSkg
uMd2d3PbmVuyq+HtyNu1hylhILSFpwVblXrNLy41CfbaNLvMGxcV2DxV74QJb8FzdfXvLVU9nyj+
U5Pbqkjqa9XrQ5KJzTy31kQLWkNb/Kyz/f1gjq1RqtzRM55BeaTjm+xbsYolxO524LY8oaRXSpVE
RPPwP+aQZen3DvDYX4/YnG/oRrBPQDkTWqVVNyU8iC4kN7ZYuZobIePg7S987hlg7fSNJlD5T9oe
2qvdDxFHkubc9JVKVBjGW+uYm0sIL9unnQ8Bwn2+OL0iHgkhlu8HQPEfvQfqAvJ3f/HuvYWrpdE/
+/dUfyB+RusqGbmaHrMchT4h1LUWHITxVd0lJ52A4/wLgSnSOu4GDsztLSDIafB3HUfYxd5cGmQM
fTsSf1+2F+E+kWyAqX/CTJ0IBHPIKBQugA+iNutDku8CTlva26a7+1Xf3PU534NRiUEL5JZiECxt
FMDxVRU/1AK0kVIMXdCZ+sf0mcmiVbftB6FUD1Az2aDhwG2TyBmez13W0+EE1ZxJYp5O07pan/11
0/C/6SQpcxcT1HffaEtnW51xhomTPOnITdq3F1LJAli/+1MwTu04wdE0lMgnGWqcZVhuTCEeLrgN
sGmB3bbmlupHkHCXQ+sIXsgmIRwODTqSmcwn4MPCRxLTdIEMdaBIGbDsfo+hsyHKBI7DEsPJzMUH
wRC11uFYgZ+crqWVNoV9bCAYP5ze8EXv/C5HsIRCgBJWLGW3qed/6Djw11ECjhqKuV7e21z4hbaJ
wJI5R+kbNhiFqP8y90TDElpkW/vF5joytVQchoH+MVX/0nZh46rVBnzHsEj1UyB79Z5rxi2g+1O/
XeQXCy8zLUBM1Wjk48TQwnp898aPdJP7ndsU94Dmg7NQDFuf8ZkOn6Kj8e6yYaEEDk2isiFjLDk6
r6GtYuhULuGx9Xsmsi0JepGc7QCDrj25LrUUKzgmasbD9Y1S26crXPoFK2DCP22HDpY72Q6txiyO
Qf5H3iB1AH8JmQ/uqFcZEvKsY2yNg9xQ9EZnmm6cwFONz0t+wlgG7bwmQNXa6fw7Mbxpa4sa1xte
X0I+b8OrTHyKnPKMUH2wb7JwiKau6kkL8p/LfOR3vaexslX21uUaeyuUp217+m78mzXXyTVCdaJr
KDxP/56+YcOaWQZB6e/p/njlFLLrISyzew9VdtIIVQp02/dQTLZY9Lc2gEdodya7/7s9qfzAV5Y2
xPtHB42S+avLz2Cv8N2BJgQaC3WWJtrkqhPl3C8RVZ+7gjYdSjq6zcRQ+9cHN7kMPzT5ihDQvpet
966HQHm+TtSt9Kd04g3Xa3OK+jLFJ1XcUGZ99qIzPzyV7aGvWjb2EyOZ4RkD+p1U5FJaRZVGbZ+z
iNZNR/rWtEmKee6oEo/ReVKA43lfskwkdypEdp7ONNV7iLJs76qxtomOqi8rnqZq0nlO72QzZvAk
V8exDdrjbPIs2YNWKAr6skPWWmWh0o85SuX1rEJiR/ZxC+babbPybOs6u2Ou9PLTSVgv/AxjYWP3
DilGlm0PEXLkR2G2OAMIYv1/tSPff1sJZIGLA4FmfkHM/87l+k7BCMxMGEoZmmNwRL8xkkWLR95N
4LAbxawZEgOBpoFLlbPSsizQGef3xLfdxprN6eAhwC0ypgl32YQHgxwTGAnlWIBU1m0mm0illjwE
/YgjElBDgQKKxk9UJPrNHPPHi7K/ax5hetipDaJhM5RB96GkoUOMx/sNMIWIqBCJK6QJjNXYY8oH
ih1bx3vd0Pz/vPYQ+luy6dXMoy+GrMFWC4h3HFikz44w09WHB7mzqTRSKxP9Vads/wM/D6w9Xihj
ZhgfU+oEnt6hb267IClMyUdBV0+aL1ltdL5JSTzHx0DntCBRcak+ki1c2cXX2K+HPLCn9tyzNBfm
22k9eukSG5eyKIZI9OtZgQ7CMryaAq6jY2z67mMXKxM2sFNVJis8XHnFLxvuLaTu7k5raDjxUXns
mawpgbMNNOAIUVi9xJ3IHqzbvFVY8iUARP3wgbcH+C+IolsAdO1B1QeFOiJNjc3puEpLeIpUBzkA
Y5pg8yRagx0X9c4Q2PZpx30RbVdImt57ft65bmdsJOkJxM/hg6dwGRsAmgbW01rt5sjpO6C9lWB8
TM0A/3cdRxt7QEQn+K2Ai/isuTOfFpQKFmlJxihZ/mHKnldr3k5stn0Q7CfT3ptSV1Yf1MUyWpFj
kvxnhZckl8/d5jqgCO+i+Xhfchw5HO5fsN+XM447YgP6UEMzFQc3uaJmTSx6ce4Mu2/JLUN8M4MC
fQwqtAd6km8dVeT2JOSabrbaz3eMNwEsLAAaKBk4KH40L9W5SMlUZ9d20SlWni2tzeXk3EKVnji/
bVYpFJqhb6obs9GsIkjkZcHcExXhEk6EYtCWJgy7RtdCiQn/Ha3ArtyQZ5XulmmHU1kMHXySTTp5
uW+CLH0ObUW/coZcJiB0h8cOZCyfoRZ6Azes9+eLZc2uYlyk5H+cw5b/fiRYqqcfAvbJ9pWEZIk9
UQIdr3UQOpQrf9y78ktWRHdqg8ErBu36/X2Ap/2C2xNJGZYOQlX2rI0kfKoPPIXcswQ9prQqxOzc
dXNCwX3Tnc4wf/rQCk16l792Qd44OppsACyEEZImNRsDw1n0+QATYGyG25HLsQHTt0dsnr+BF/+G
GfMFVISLRDtjozRR8zYgZxDHmTRt/6Ng6tkCjvnI9e379/e9+TKfuccigdBHQu576DvDVEfOgDFN
WYT7WOwxP6fImRQnAKZdvtX3+EHf32E+IeWAb1Ghmfz4ScWoaIBe0HGEN/UhfHGoswuiGIi72yg2
uXNg08jOyBwf0dQi+531kwfY+13QTsu8YaMB+Lp6fhKJNPG7wOLsEjNMvIZcr8qAFBBuHl4DX1JP
NgqhNmu92ZV+09lyEZF3hMZAnLaBL3RNXmkqe7kVuu43rBvmHK+rSIg1lDdPeSSjZsqHaP3k1hL1
piEfyCmXQqu6/euZHQDHaXR0GkTiATURj8Kn0hFjnfV3YxbXnkxMJzFAB4cJVASSWZWYmvrw59dv
sl6BL9Lhao8UP0OysZ6HvIsYM/K4Ja0ruzbPMGnMALOlhrR3BqPU8iAWqoPOOVi0xN43NpRG5Tcc
upH9j4MapaSM+NiQdKaQMfvW6VXOo2/j4+uTwmJ39iHplh/RRVSXdlKR+39/Dx99KmwH0Tqm9ckE
iyMPk0PCB+y0Mn8VhHheaMN84HiaB7ayf+ythu1kRVtsVdi/ZCh0bTbUe0wEHi3Vr5uKF27FkvaB
YkDaXGSEfP/jGxnZtJjs19/wAOoiBMAOlDDLEbyPVTbD8YQRaUzEtAOpCy9AQoAZCG6/L9v9TRQ/
7evPzVIwpuNU3R1yAPTCCQQKgCK/8DPIIdLWkkHwCfbZeFeO5yhJbfBFnGLCoPKkWoxQNTVfUIgB
5MpKxW8Sgho1obsuHKPcmDl/qv+E9oXEz5tQH14tqlOpBKhyk8lPkSbfZpUnoSipq8nCLCIw6uWc
AeTpYRrmBIZmYixVO8Q9qeGuDovAlbIXJlRotopQKgOhOBeaoYFiZpzyOK/xIdoka/tFdtTbYDjo
hBlHWNQviwL8LumnIsvERxgZYo85jPxncqKgGUoiI7qlp+lQd2QKgdlZFmGpmrVSzqxsa8uqQ3xZ
18zanmkuWvHwmcZQVfRiIOpOs+FPNbHtEZieSLI/huMuoo6Z4/cSBxmgRQknTwu30cvxu7J/n8uP
7nI9eZPh0asFLQQkrHU/DNMotzVWJvWJ5PxvlyFoWEGR2wnAoO5tccDsedshM0dt7KT680+d/ttS
86b5pjNZYszjqPZ57+xxu+svxdCdHuQ1MRuPl0rhi1j86QHhIWXaSYRSTEXmmkbE302ISroCvTXh
6fiPotClsdTBGXJtUqXVbf6RdDQkbFsAytVnm82sdEUHQnAYXPnNLoK57mSUXiRWuuAZJG5x0t9Q
cndYoWiqlh8I/++SnX9pbXtTx2RWVfRloKUTkXmmMIyF/I5cBl0hr5ZQK+8KkR/Zd7w2Eu/xn5D4
CIHf/+iXg5Wp2Q+HzL4k0WBe7wJh4XcJV9+t7irghEZzcI/7D5hMxqaQQ/ysML3Ax2LbdEMb+q2h
OjW+s4elwKLFgoBrXHukZtbZEov67abphf8iIUL8AeJsyjfIybO5l9yT1ihWtvx8p/ZkeNChL2mk
7r50TzhgnRFrKxrU6UekHiIb/oKo9Js4959M7gfVEpb8tDRYwBtqMOURr1aqDq6q4xOm4ayISnL/
FU2b/Y7n/OHQdYPSm1TRSfpV56w28NtJ/BBZAWN/BSSQzrogDfUXEb3Q619OqFE0VyBt+aDrjIom
F5aMJcArv5vob97DEduJpQYYq78+231ktABsv7k857W1Fxsng7szuVPLyKPsTVyYH7aX4vwU73DE
EBXN5/2hJZAJZAbnG5FBpyDKcamqg4n7UArBSKPpYdSNIG0IBhRffU57eiTchiwaUYSzI1TpFsFj
R74iiNsGZrcRDJfFqrL7UihY/uPrFAys9u3MP6Uoe+UBGo6WTidIxWYjUNrrcsOz9+wfw/NKJpCy
wc8a24JJh2MejwHSQ0Z9s5pVaL3EuWheRxIirby08XUSsHCDXlf/vBmiKdAo/G2TiQRxoISjZNWz
rF0y3ubE0GyseFfv9I8tV0JE1nJOCQHzItkKv3Lz7lfHZ6nAk0NN0MTEy8n0+YY7lo8P9y/dYbzh
eGDpPsg2/I03DJXwuFpUOtk8tJKxkz6NzVR+a7tMNI+dzP8Rh+BcVbb/6fc6rnSAamZWonFS143s
oyhpAVFGm4lbhcreygWVaYr+zlSephfXdsUflKbaFbQvco1K4iLSCj1VDjxT7nySRAzC6eBuVLnE
z34JQBkYC0mDXwAXtgiKavpOHMoOYQQKVr1ymrBlYCQmBnk297guErWXb0qDAtPmRIa5+X1TVWjz
EXK7EfZw/8l0aUVtH5qjte4xnblu3F5Mx2JWn3w4tijuPr/GhLDBTKm+KfLa1wQ/mvwkHjNaGaBa
jftFuLONKpwesFDiR/SMaJq67wnr/XoCZ+Vo2aIKldXo4dS/ppm9tJzrET1UeZEZs0x0mu0GE4UT
l/C72hzJHaG9M8SW1BriLV8cOVGQ/hCiT+ODKFgUueNTEJQeuxxd1938hqHFgpDtfyo3TxAIOsxb
/FeE4sSVgMcYZaoaaXzj+228vo7xi8FSoySEqECvU5E9ksbhfs1bITIJ5J+dSgFHmkbakrDLm67z
yJ6fjTDjPag+u02exg+Rhy2kfbTVNiJv1cB7IdZQxIptLKpATA3rSCI9Au36jCOHnblp2qPw6aIq
MSPEhCRtwy24vGa9DYr3ak13xP57PCywcw7EzaIOgl7kGFsdu0iD3aVfS8vjuwN21w0krodBFhkW
m/eoH6kcrnWIQYKQK/RLGOgDEqR2AeCqR7rUAp+zLVT0UClNawGrKRqxR0b74v8cWH98Z5b32I8g
LUFv9UXiRJNx5+HZrXnH31e2Qf7Fg/JC6EsH/z9OeXTCccpIYtLyyzZFDGOe8D61elwCq7JA75en
scyYDM8dZPjspe8FSvsLZeyXxBBvyKcxReRflSRI8AfiVswCLvuFC2D05ZrAmcwmkOiYJRlHu4fM
vzU9zA1Ag92YcUZvodNfOogjYtMEkn3CW1kBpxtRoYJQ8F+xbcO6LL/tWcGgoQSt7AJBT4k6PcEJ
WHr209gvvV+uS2Mnv8/gVat3v4Ii9hv+62S1eRWPP20lENdPy6iYvC3q3FvaYE73OXCUA6IPBCcR
DIhh0BQcRzI1Hv09GZjtMHNRobtexi1ZcM0FrYy5NLhyRVCxbED7iK07IyJfybyw+mfKxz9lOLz2
tlX3MfJDm4DZBb9LYmtJAi+A64HxkO0Ped6/HQdAIDpyyXfmWhr/LIDruJUbeEfRJvptr+vpL2e4
qOhWhPt/KiLKHRnNozmfSdUJJRtAo1sT3ipzC6qHhK8Ieg1UUOZoe+RMVnQ8Ewy2YasaPf00Mp0K
y5gI9sVnrVrn2Fs4Oi6HgnSmlJmhQeehZ9yciGfBwhDe9jwIYLYZOZrpxI6QJY3lYqIRhvZtROzX
n/v5mWmsbFLF+5Gylj9AcEaKcP+LXjJ7W5hqJu9dsXJIcKbGVm6b8DDt2Bodlt9Sow7+UtfFq0Sh
3+MotUHKdfl8Xf7AxFYaE5EEGcKVpSv8zjgBUuuU3EFWMsj8xN5yM4TDCAq/PBToBcZdXDRwRN+c
T8EP7yTCN+Y+iFsoKFQaPCW09lu91JLVJl4fEsYHprxf3j8PoQxg2QuqkDA0DnxxuYDrfm/HA7QE
ojdNvRMmdqWxYxC7CVigPjJvMFXUZL54JOHSD/eU9GPdDfmReCF5QWwye+pl+yD4T2w+9YW56FTZ
tFyx0NcaBdhCI7R8hy2DbUKCppYbt68lE6b7HegUnx31K6DNb2076ocYp2EC2UYo/gre8BQ7LKRq
zmogGIbxMG2EQnxYFIoSPWxXie8QKou/JyVDYeosFiLA1xXr7zmFpq2MderDTmt//CSVlFjKxHQ2
l7Zi7Saw37hSf7lwAJGmk5j96lIdp61kqiByPZfw4d9p2npnaYqio2rGNxQ0i2VDWQYpqnpY3soT
2zxNkDSpDqsW2PKhbwrfZvRzS7yriMmEf8IwUV36BaFG5Lgo6k8ffb7v50c1J625MAim1+YJ+psZ
DrO5ngz01UPJqCZU5hbhbQxGcUFZu+Va1nPP5q0EvL1J1ept2nb2VRt7PgXumTbwTGpDyN+8kkWG
Gvb4ETPxvQOQ+tqnLbzYJ/JwLLBwujkBInvROaX4nP4Y3nP0QQnMSVUa15/fidUN0sLNFR99yg5r
YNEDiAfNyJWboktl8sgKbRiw/u3csnqZpT+pCr/soZbz8o57nYg9GJ+BPh2qEllpC/pNDwfOkSzj
IfT1Ui7p8g37YJ42hMsX31yGIpoLAB+sPty+VEdFLOssxcsJY/m0FDG37BViUMujXVkpDDwDp5UB
CfrKRv7Fp51uR7QF7jh+eFwavSZbnd0B81Qfk5Aqq+Jd20IC+8Le1XP9pjO0AMpbqfw6HxkbXZ+7
5tuljpCz9pSsP/Av2wVnyCHGNj1alh4GaZYrY1/CZhmxosWEnU4Kdz+kqgIxSpfibzzuRfc5n8Uo
bSlXdGMWX4jhVZeemaz31Wp/IPhnLtz3nrYKk1YgiHFHbykunkPXWTR1EGwK8f4F7dQpwkK011xl
Au0HugeqppOwl3rEVYcDhAUJb8MPGL7wQVker2n4PgcrbQEHJWl2yWTpVTIiDtY7bN3jHVLTRjrt
hIY9aVza6XgYG2ld63c5yetwNXtTXY05XWIfDCEjWStBJHq7TCNtdpH0mkaxMjgit9oq35wY866E
givERGSWoxiKWlCOup9FVkn/CJzZo//sWeeQM8EZfiE9ipUMijXt8QxBC/Q8EVkm9ksF+wv5ltV3
6/o1pzSsHGIVqabH+XnzuDHYmPYVOaSGguY4uwjTvnkETfXrW0b7TVsovU1ziNuJNGeqlwZyPyJC
S5WlO5HtvBVfR73bup+htGyPKAdT7Ywl9kWuUVO8vO59JwMENrQvLyeavwUCNyRP9ObafAImceRS
PLg9ADoqW5CpXjoLOSvLV6/DH3Yg8uQXStuyQx/V3kKwLV6cR0wcESjI8aIMty3+HyoJb7y/9bwb
K7ArwAND1DfBC5yz0SA6uneImVtD8Wf0m1pQYnZRO4J7TiDikVViF6Rkg6A6ixZUQ7X/6g5MRPcO
YTEOEgxdDAKawk+BpjXif2s2jTaxR0zTtraDJJ0wzW/uXaR05yAVVhWnRmZGVPRavD2Avm1KhCAo
xvdY+KcwEsK0bk+yJwFoAqxAJcxqluCPw/Svud6qR96TveKZT59HZkylgj12pc5jPUjXVkd8FhYA
BA3GRVs9n7r/r7W9OM+f49mjCifISgMvvn/UtuRJrBHtNg/S8k2ap7y2HUjfSnXLWUdFmNd+5MKW
nxfCY7c6ylVrt1jPdKz/zRQic5BRZCrHX//0PzHJSo3W7INDDPCTd6IwYbI8KYp/fe4t0ci7s3wb
RhQWoUrBL4gYuvau9FruY1fle4lgurCRdLZpV4RnYpOx7xaCdq6YqPXA2ae0DuJ5zpEjncxDpCha
VLkfGUognMfiPtBYeBFaAH4+bXOjKJGmEszds4O3wCsqACfRN09VuL+RyTNMSuC7glSqX0sefmCl
dijSoIrEZzR2f0JeSfgdkwY3mLTnwaHgOxIuYxo9luxNo9l6LthnpCwz0oE9UCJ2YVRhv/dczwoP
ytSHVifzptoWPM6nA27KrrHKHkFlpgiTc4Tvg88Vg9yZU0jP2MYBsD9GsjZp6MI89QUXXJ/TTsF1
ybFppQVNK6FDQ88PAlppRIKwaee0hoN53OJVE+qJtGvFM5ZU79TNMzUheRDiRtU705/jCSEX4gGe
ohjGK8B8GZ5eqax+JW4SQDNMz3zeVl3Zx+NX5Q6ZPrVU12NW4gwKlWHsH8MGJfprG0pukHJKEmHg
ukZR2f1puTTnLJuAIgGKH/imrinNswwjsWzAEFPeDfIfhIIOAqEZ8OCFAIkAqD02fwMPlaqouFuC
UvT4SWGOrdpqBE0Lrz//N/FcUUOMpVcYp4EK22owmYLAL91KKzikSKlCEL55PYaTcwgty/u6hHC4
fK5i5r+NlORCDMffP9/OYm0+Cz3rYVS3NcnRGSWomZSMVnN0KPDWDNdf/BgLeTchEcPE0x6FFSrB
q00PjQhQMT3XOCs2lKGGjSOmCEz0h68VjuhxdC9Jq4eoEB9YWCASNRt3QEIuPAQTuBGiSIXjh9oB
zmp3JV1tQoQXV5hRcSqUvCHXetdgHMbaR+rVMZTjMOuoOBsoTK0JNLsr3ar19Y27j83ehmbOQEtn
CgLZAFbJZPEPQcytp2jPcDnxgcAztsajfSs2Y0Q4S/JGnY3HNfz3sP7aTBCgv+MY57FrTqAsdZBo
3wQWVYeUoIqaRbGFhYNTgbnYhcaZWaP8pPmTMP44r6PM8DOEpFwcWcIEXAwS8vqn4V6P0bcFEHYC
cxhjkj3y+WzDAvw3iYdlqDMUzE51Xcai2yuAvdtxDtIylF0dA4GqqwQDfGlHdA3S0vX60cwAmmbG
QbcdcVNe0lnBgRgGCdGq3Xy27AoQdF8u4pLem59WFNRGduHPjeK5WsEXe1/r+RS8h21IpD66nwha
ct8PBQgGsZ3M+j7KGnTxYJ/t4zkQ+wwDZthwafN5+yZ3jXh3wS7KLzDsmn7dWvHRD39igsGkGcc+
UrQMZTpRVgF+smDLdele5Yqf/0k9dxM6NrmIKqOyJTSadOnlkGvShuWLkjXe29NEQ39tBaqFHED3
iD6bsnCGpomE46b/zffqUfzcgwuvWkEg/VWXyzLja0uzwrsGLACbmAMQ7P71CPSryaDcDYHzOY1Q
SUrGxFL86MOaf41CVglb3osTpYxMXkkJ9cZxNkrzaRs+/iPrrujigKcr4w+2cw9Ebnl0SIRVv1wq
AHyCS9uJtO9eHXVFCzWDXYTTG9NfvYZre2LrA1jgLsXkBRbJ5zTYpsASf8PKybChIOzYXC9uc8io
+MlmmiSJL2iFpmPgSLm5kh/vrlcF2Szo9p8djXkCP4Zfj1uZv40k9mRNNKWHxvj+Ji7crHnIzIjm
G9bHlALzGTiWgGVksnahqU8ygk6Mzk1akBm2gfCjKMpncUx+QxxglNSuHx5DY4gjflNzmDYmtH+D
668TctJZJvnAihNrXh2WkjQ+DsTE/teg460dciVFplPjF5X4/YadQetGrrcJGYFEZ1OuRLR2Z6jF
H18o212+/QelmZKdYd/dX28OV668flAPZwciMxtosNDVVPvGZPP38aICoLNHRHqlPdZ/EeK49jj6
ni4uLfnvC+vdSUY8jsVEABDRMO7hFScerA3c2KrDviEWzRU/krFDhLlIrXncumodDvXqhzBRt43C
pbcNyj9WfuvX1z6IdE4GeJgA/3PwSA8t6OHowzL3d/9T0UdlY/gjxQeMOyKQH65ftWa5VKNAzLsq
GKo1/0K08wcMWGbgOt7BFisDyQQ3Md5CL0NKQou6XJHSo13oVhveNwBizVvnOY4xpoPvqoIHz2+L
j8IudeJwpvg+J+U0QbKCoico/8bEJOPNM3EuMoXU+ROfuICFC3RLi9gRq7GQo5wlphndt1+RmyGp
SR3Xid7m46gDnc909pV2D/K1LaJCa/GwYXL/KcX6KvnKSRRMMJ8HL2qvQMOgxObqmtNZVgX12zHG
4UotbK+2DQUAfCP/znLCNtUBnxa8llmShgzkLrcunlrl3rFZ8pE0isNNUXrtyNLhQCdZAy0Q93li
xnKoaslYneEdQG+f/vxexj47SsqM3n+0DFfZNUFxCnQaUT2G4fMEs/Ai66hIxSs1YrVHXSJNfPDe
KaLSyvDMpkjCsY321wSO6BR8In35HFvC2tygIlP8RLI2hXYqmvsyLp8lsTApbv+HrwPLx56+LIoV
W6FKbwKknV/kpSUZhQHda6oWSgS3h6jeMFRwArcWRLhzPLB3xTYVnHdGCcfpda1S9H1Zvg41sGtM
e+ATvbV2aP0jSOWJkf5ottN4NTBUQCKL/Zz1b7JIqxCq7S+O7YNI5V/NHN97B2Tosef6gvSjLTMC
jWSiul3aL7fQnJptR6PSynGCoYfWYa/xeSF276hX58qaCQatiKjxfusALhYi3nVShma2dYx0FVDu
kSxXv9rMVZvJGJkhhyd+TqFtaVYOYC9XN/sgP2w7VdqT3zpjOTwtB507g5EZd+ec9svhGKIJOtVr
ON8Enu0xP53V5AfohksWUH1EVvMmL/MpCLYR2SlVEDhjtR42k9omTja6q5CU+K7i1rrJqzADiQxD
Mn8Hw54yLx89pJbRW+/TajWcnXgj/o6E+LJpNrwcP4G0FVlWTRNAF2SkGL14e6NKya9RdBkfJ45I
kkxPdgkFdLPtKdAtXlVvkbJhlUY+WWFO950wuVNqAh0sanJzdAhPoKguXJO0csIEz/0bXDsDpG2w
zNTfFI0hxuq5ccobUdqlPzR7nWFK5HaO0SjSUXVIOMyQPJU1kWgPM0QkF+OkVKMnL+d81w63169Z
7v6EnXWQj5fj/5g9ixLoTPFlkmAUn66BEE5AcAGuVGAJ9422jrsATY2OZcuj35PqQdyzqjOB7gDH
A2/iGcN9tzRFdeEeC7OzpzthnSCtr1Z5d19ucx0X+7Sldo8DDBr6OGdp2HctOWpjHAPVc6ZpQ5Rk
UQJb8zZgQ5Op7Ck5YLTStmfiWinSn1N2sHjKvdRr0uB4T3VNnzQ2ThU1FqdkuSzAGfnX7/NYdzYX
1i9Evk2OJzQMFkoLw5EGa6Lyd1YCP36FvAE08yiftjY3f6Rec7zg2vyn0cMkNVAQXZNICILwe3oF
FCDjKBdO9L/kkv6o0jqRLxdrYQqFagluMBZpQ/bXi4IYIBEX6lEsqDMJG2CjU93MafpsK78k1TJr
8S91nA3vB11BW7A5RFbYMTx/fZcRBji1fJOcGEVa04tHMlGWm8qHL/Z0wkiB3xqQlsExrSzTmLzE
ZQy6CS5mkLA+/pBnjH1uZApFHqGf6srz2aObdal8Jku3JS/1+GjgikwxGO+ynvEX/zO6GscxVOEL
YjmM6dqFNLIlMo2zz6Xa8m5TXD4VOxt+x3/0V6jLZrInkC+2PqWuDUqoeKBFWSVxmwYtYMlv/ZdP
rpH32m6tsBEWnz9896YHUVSXuRoXGbTJAlfHEP69bshoIbggXvb0eFA2MrWf0BpMCN8fkz560A+l
zKtGKxywd2nWN7dQfgTV6kXQ+2rgb+WiFGH9gkgXAL/r5BA1E30oIsXVxweeNzgLe/b5WyHMcIHF
kMuhCRsyXq/p564Sexx2UOyiZx/U4kCpc7esPkcZtZwo+cRvz41bhNwL1DANQSv7luQ3sBs048Fm
mr4c6ycsB75UHh996zlE3bW2AwQosytOFHL8grOWkgebDPdG1v2jG5jKeVwCthULloKnb4xxeTxE
XgEg4j8vg+7szFMsQ9LNWN4F+PI8qUyb8T/5CGpgpKEf0PEFG3n91M+yUJWD5oxSKOO3Hj+XJeme
EOEoWGB0DxC7sXxNCmq2UGn333oPxJjDTtAz96bw3AESjCXbG6gGXiIKpjo8WKw2BbfR03CGPstH
3YyvKbNkCTwQmf1CHN04FHM21S/TQyzuNopAZr+MD0JR3jlw54Riqr2dJ174au1yIHZUjASHreQb
BEksPEG5P2EQJcj0xmMtJ1N+VxFFiv0d/botn9r1WufHxDfvTX/DZGgHlhMezRqdR/AVmeU2Zloe
b1KnF/F9BKpAN8DL9Cm5zw5jNW1NZ1u0rcp5uWKVFtQSr9wti9Jr6eP6Z3fMRsUNFL5+oU1Tzqo0
X6C/5ITzt6pDZeLSn2/tUg3toeQrRAQ9pZTkDfSrUEXXpanrvOqE8hOBTU7ezSPJf8C/jhpfSYSW
kNVudouuFBq8I4KUp9/beyywLagosyEwe2EvA1eTKOhF3mJASgRqCj/0KlUqqZmhC4oZ3Ma1Mfkq
3XPzCROeytfIkRcRlrada48zyonQoZ7gV0y+kANtSBbPy4qozXimYmLOp9m+rlKn3NTfkEWY/1OJ
OJlY32XMMQcA+ltTfMbTxH9dA/FQJzdQOLMJUW7LhQjjtLiBqqQIuGYrJTgiluWdIfFXTnrBGTkH
he/K9Ov8th/CE/QZm/do+EmdvFKrv8uBV0zbV9CbXfWf4xbjzIZHv4u24C0xC3xSJik3ANq0Ppq5
V9Sw4ADrPTpBhVo57h0WQGenJc6uYPRVrrKQe+zx8aaUn/AgOtAxnVC8kcr2Rvvo25yzbfLyWM3f
oNlvFSi5/cszDw0Qe/Ouupxa3cMWbK/nZ4ry5QWYmhoDHd6EnFJFfU+6DTQfl9/pAbSdk/JgTnSJ
kKLwhzyri+kKNnBsZDZ8ZV297z/IZNbw4ER98WA8sCO01ZSf21z/IwxqqsaivsORQlLKOROtmMrY
s+PjPQZrnzgAjmJwiKJzWJ5B6C2jYZScNEZynoGF1OVo/Drt7+98tY+Z6Oa68awIt34l3eeKXe61
fyej7UERg+3qx7JRu5vmGXD9DCSAbuwJ76v96BXCZzfzgiarPIB4l7TZ9JJpD+W+0pDZJHbOvuu7
bYGmxeFqljYQs7zNo+IOaXhjbuI0wnVG8hCM2cZbgRuI+CEdZVGVX6LCh8otOSkCrz1ZgexrZtnw
22d+FYWhZRx5FefPpGH4ohOF3BPo3YF1EvmFD2c2wPX4PZ3rj303GE1G8EDBvZbv/yXtNnylKrRs
Oc8TxXfRUmkDCc/wtcpKwkH8FEuQ5RLsN/tp+n6fcx9X+ShemsTn8H/CEBu+BCHBSCd0sIba4pIu
DJA589m04XuxVx/m/V09iRu250cRMzNzB1/M45KG7LK2zh9l/1zX5qrwj1YTphRcGwIU/sGL1oJk
tocolKv3F/uTusw0uaSaa6PNNmRv18UGSV6iLA6H//qTjrkSCAETxr/nDy8HSajhQJyl+xSzJFp3
Zs00B0VJJBGsAebqJGFQxtbfUBR0a8vH7RAuOzpw14mBiQbbHMwUjFtx/Rz07TAvTE9zR+u0272w
bRbjjSu3UNyahsEwAIBI+R+/a4aoZ44mv4Cju4hcC0Zdc73rnp5utDg+VRqqQME88oiav6uUDy5v
/IBLFJke/B4nFDHvJPTHlDuagNCZuB8Y6EnTaNlu8uqUbVXc50VIv08J95HRjjYA67m5Os1alN5s
fcyFEpa1NLrQVxx4wCMe/+KEycaLOOuK3DZu/cSzuSFPiIe6xAEaUZk/dOssWx7vYGG8j9LSY8CY
vwolZAkt693RxwRhJv7IzTLkImzWpM4fVuSWXXw2TAbBulCtQd8rEVudQC1+uT2OQc6QYUaG+hqs
inVkvF8/rA589ZSVNYALnI/c5cO+pgBkOf/3crpwPmN9ALtNq9uTi4dVkxlfPxKGO1DbJRKHEqxo
DIMRN80D24sr+nPJXDN7nKgbkPwZLj7yFmeFiw0ZEeXwodnFOq0Ljur5t97D88MBUb27dCni01v3
yIawM8esa5a4LebUUe/7Eu+E8iQGeugTtkBTkK6RN8EApgL/suMSaQR5mJnApiZotDEEWRVzxHrp
parU4MtzdLSMxPLCQX2O5M2JKl+DlfAqtvQ5TPZ8wt692aYNqeTLPRYNilAmcbKQwris0UY6yqqg
RBXDTVxRN5DHPKT22Ltft8BpL83AkaHlUHlgHDk9EzXh+W5wD9sE++xVtS4gL8Le9+GEqByjD/7c
QpQNM2QqDpD2sNnZ9R0VzyJ5Yg/FK/MVGB8OWcWLgpWOTcnI2K9pa1mspkJmXk4FQY3E0NuBAUwF
9yFkxKDCAAVbnkV9piyfiueUqQutKSoQu5F0GYYVj6H+7zciWhJVV6VZPlwWq1UiyyNR+XS748KO
NC6GPJ0F4E0NWFrnpkV1MYj1xsHEN4M+7lSVMMldmtq19F1r3EOvR87Rx9hEJF4iXCeAQxvqZuM8
i3PFNDvDERNYsTVe4kjfYjJ9oFcSWU2U1hgbqLRxhB7rVrDLjaEd/M124zQykm5XVu7dGePW0rj0
WorKL0k6uzNQDj8AgoYk+EFtiL1/NCMnEx91tyZyWVuzxbE8o7Psiiziber6dZqX6u/vdyQa+Fou
/hiWhJ13HJ9bWiFPI5ivgXtqNPFnd7NdCEE9dfJS981oy+OTyf6FBr9JCkdPHnufF1RjdRSJO0w6
y9XpKpY3aEljNYoIpVlgAM3icvW4Gz/yHD+hjRgXWfF/6z+YIWk/ADG1nCSyVrnoPNCQ4plmEuJC
rNg2tg5hmU6k3Yww62YOy1wlAGnTTwALPVbIyWb/NKHs52PVRLuL6AfnZoibhohS+xVUor/INFgS
p6RZ8b7MD1PHqUAe4y0thmK1DIIatjizW0pqOzLiJtdvtTMlYDtGE/rB0XfLKR2lqezawJQtcxsf
lIIKW5NFVrMaBxXuq65Z8QLZh9AKcqWQ24h56lqY7SoOqdYJ9QLPjwmyNlO3l/lcadB+NT+b5/BP
n7UHTBo7CC/vQ836KI8Y+AFULUxRPYo0tsWHmpzbicvUAaILNMunAZliN2a+FzoPN5p5NGQ/pDr6
/pz2Bhvn7wAGvMh0bcuJxwdL2iYo29HvjB5oEiVv+7ehwZpJ1ziLIa2YtATYZAmKA7mxE6GirPSg
vivTCB1LHUY5rtsghKf3LOxotx5NAj828nacCZZk8L+Bo158M0iyZsV3EIBmcRwIRE6akr2Ls1BI
l6OiCzkXrj4y5GlWzKAw9LsDx/XwLpbXiGsLVglc69mjd9rbjcf6KQE29DWMSmyAm4+g6SUshIxK
JcSB5+03lsJ2RY7+um/YeYF+GPwPYRMYhWKVjYfgSZOcBRp7BPylgcTUNlRkwSQKv/8ch1CNlpzT
hHvDelm1o4ynY4EnPuzxHxp1L8D3QO6pyO/ORZ8+WwdtqYOWY/jfrEhMwgtMZ/o3fYuFJzFXNftJ
n/tzaaRtoVxGEE9MP1tcAIgQcdicpEHzoRM6a9ftQobiVD6R3jte2uX/HJ5xhxzqmUmo22yAldR3
leAcUfTPuMdnRpH/Xi3o6q8QBTahBY61HmwPxrGwSG1tJaZ5ZJbL5S5kX38tZWJd9z/TCUXMUaQo
5TCXc9tHlogxfb7YuDlDNZCzNUP5753qppa0vUN4CueVC5R2LQChyq+P+daDoPAZ6VHy3VnoxE6T
c7lHTHZ4bhz3tHaQpOvw24ET9t/QPdQ74bVynaGCzG/Rm15pkAu6PeKIE0rrJEgECEKzK7i1diMi
rEUawt740UHRn6JyM3oLDucY1TSgFTaWq8ljLFc2tpgobh1Efhr/1/+IaLtG3D+jgAMGCdbmbbCa
ZGvfRWozN3tkhWnCeJi68Cwej2KDwlrzJmTk8Magewbw8HJoNb3fdVoqe1C9n/z3m6v9fa6RQHfg
CITpDg76FRGAesKE7jp7QtAbobRjlgAR6xfXXARj0XMJZOBN5YV6PN1F8V7vwQyT5Eaz1CqtAACk
2ro4l2AOA4a4NsuoaiJ860TIJl/q7UUkzoWOF4T5AFwHe/8I/KzD5SF1WLczTTZgIj0SkR1DApX6
DdSsXNQgVXDgqBCEATgLLwnN/L7J33wUuwB9l9cFIIWw5y8wGftD3x61iJGI0x3IJ4s347HwjFF4
tLrZ6F1wLfXKWF8d60giTotHYZTvBHNSmEQUJ8GEZJSPZUIeC3CGjDeRiUGSCC6SjoFYSpYQdsTB
Vyb0bQFlLF0e1rt5aWlTxk/KJXtcGhW9peJ1+W0qlhFUz6kbcpvdq06NFSRKsRo8B+Ive4oHxdR0
U2+sZt4W0p/kch0oU8+lPcBI5IMupX873zphyhoZ7/JH/1wcbGyIe2YctyTvxvEiKFeMRuTW0dqS
/Kr5uGT4Jr54vtvphq0KAFuYIhYscBzTZsz7BtSMQeRP1UcHzayRww2Jlm4mizippJG4yuFVSuSJ
q7n22kCyz5IgnWjyfs85ukb+oR42rZhzFYK+s035xSKu5YVkU59N59rjn4Jzn5L4wb60gMyNm2r0
hwWMIThVfxvPsGcbSN03NobNGe0PubPWOY60WuIS6enCWS0b65lXZryu5D/AzSaHe14aL73/cmxM
/PhGYchn2lIqF11DtQaOrdRHGtGy/uv/Ay5mYxNNNZttrSkvfaCKe3IJPqmwNMlamCH46ji9BHWT
mNRvATySoRffhbiejAchYlO9A9C6NPz+GS+Md+b+NDNFTogx7+FzGuXYTXcBis7jR73swJCtYRCE
TwMI67sPwCBZG5yJl1EwhvxQtdJpsgouEAskj4M/r06q351iLfo0Bcsbb/ec12peErZlS1biioEX
lo+40qUx68yuWfSAeWus5/PSSRFw0VNTLQ/ogcPTBTyzasQZhXr0MtmOc8i9PkC9ojlBQ+fz8/lR
gKwS2TWWyffsOCcaodaIjixMBVXreUyIsAuriZ5KvJ0NyJVVJLtwtgz1FzhuhLQ3DqsqkWxxpTqo
CbFKJUeTeL5GRXOU865TLSdMZ9CVgP+65ONjw7x1C89JoO9nQlMgPK4kDghXplBgOQd0yHjKnx1e
iY+0D19CrFMIg26s7tLxzoUHIELKjHVaEzGuekGEBSN6HA033A5g14//b+kJMIHGxKKrdgVk3SMt
DNQ4XWBG/uGxq1W9nQczYgQKR1zQebEhN359AB8HbukgiMplqKnLSjavodkMp92r6i4ln4obCg+m
eGnPYCJGwk/CKYBIlkN8LBwaqOvGAFOTIhBm5cnuUInWWRqNrnArCLeVZX18AJj0NjjkLEhYk22Y
mHP8f3Wsq7bJf/AYwa6rqG1ypT8h8z0+qjfl1CaMSb0xz2CNHsBs5ds4PFtImxrfsX72qkM+dxxd
iD1natWZ8KsiLEGzuP5pVsPyXF/0x9ZSlItjwKm5M46LgAm+Nd32T/7+bLZ+z3+taCFW7H9pztvF
V2zjP7liy39iGpirMbszdw9n1VJ2ozBHflcbgOXlk/Msctr/B006y6mZXlz64eeqVPGT/Cwv4AzG
TOLoKFLaJj/ZdL4VyiFUWACYCpp2N89gdlN5PxtFSA7uBw/k9a1ppTNeytjocP/Wp8T92Czh+JP7
+MIk9FRb8PxpxMAQBc2oh/SvnXrAzZMrIZ196IpP2hKKs6V6aVOeDxU4nI/85GgZyKU26ObFD7mM
xXjOZOvi7MYalpNTSxYSwbCRTRDqTAbZ0ykICOMRhZZ+jZqkxT3D+jvv+b8cxaD3mZmjMZA1Wl7N
+FPsBvhhz/DGx6g9lg+cearbLiFVuAQ3ppr5+H8GVbBWTLTT/3ey7+AZ5LrG4vTURk6mprvj1IFi
l0q7kY6AewfFXv6bKS8+0QIh/KUwuN4a9IEB98elqn6FCZiYGA16K9V2vNFjpKsGSvzz5N6S3TP7
CBRyG97drFMEHw+KHC9V4EmzkNiY/zcXSM7HV4ltpJNLOLab+uRQfY4DoEvpuLBDeHi6Vj5mkMab
rHMYbjJRqriOcyVu07RH9CA5+gfIUv/WolmBI9E/IcXzmVcJzwrHUecI6QvbmKYJAsmeHQFN4NM8
yw6mkhESFZsdrnfW/M8QWEa1BKIncwUbr5lWHhcnX7OlcnPBMEm2RSgjnmyRBWT+/Ec4gaRNt5G5
VPVXru3DVO5D9FrtpqMSz3NGtY+/6Ar9qy33KqJPHndFw1pBeFQBDYcBPQ9+nbErbAGIQ94x0T5z
btvzewjzGcYBefMQlzsQy22AukNzapEMc3IDILu2wYi1XEMM4zhow4bUVi47e7C6BO+LZ6rEKEe3
u5bCgJkhrLyFLvB1xYL6uz323Crhs/cie4qbeKIqn+82FijQQ8lAJQ/c1mGqo3fPp7pMAvTcD58a
7BydxwAzHkobmty23s7fJ/WsS8UTGzp7nwiCz8KsdgIS/ExK82/8KLjvLpKLzJ64nW/jlRLLPI+G
HdZiZQoRD+FxSD/RJrjmkNzuQXAMrpT2oMLTzVdy/tfnaf4MMEbDPMBerJy+kI0+7fKBROg0Nalt
1NQOQQ1MIj2nvHt/BgPCO6mGTaeD/z8y1TELtuBLO4GXRz25qZKqbLUIhgGYsCrxrv+ojb2F05TI
A7EM9GlqfXEdC9ChZ0I+LYIDzdHjPT7jhaNzUPyyTWbrvjcGfR0/xwnW5xNvu++2M990kG8RY+g0
JvaVIM5eZhWlknL50TPO1CMBzhDecE0qt5nFyq6rlVox9GnCtAiEaH/5tth7fQRGReEjvzOE89Kk
pEXqGEsnF9QuxYGF2Z3E3jCan+jrjOooSfKi9NQEIi+IbKuQPPoOgJfJPaRiaPcwUZFOtCGAHE3z
EvR8wgj13O2QpJfP5osMSlvZjeLblAKhY1LcBVeWd6RxoM9CXQQKYhME7QF7QQv2Wzabjh4EgIca
SZ0VTz+HfBFW9fwEyzeV0Ud6C9lL2xRuhAmT+IyDtKetxSo3Ys90KBQfUQPSqn+j2xxq/mTES438
eHO84FewGTBQdCI9gJmWxpgyXbz8qI3HJkFz3ar1RCD1s1r7oo+dGGC9G+45mCVzK6OD/ml2MeQW
25U1JYsSD6JRZA5X86VlA9eEUXiAssnhDzOgGoCo2BV1i67v1WNZ9ys5jsRhZLWtLXbka/KWmres
8t5zJ/prpUk1QpKKRhBPzXA8Z+kv5Msc4c/0rsKcAPLq7QrnEsFuF+uU5mctGXW4mI81DbfRigXN
Sea7AkCABQIMKLlAJy2+88Rt26dlfNjiCWBDqo7IjDTYTQALX271BvrS1uzB/0CB56JMbrDvs7P+
0RcTep3ASFw+yoOzcpjSpvig3q4rVBaCOcrMBKqVkw39S218beCnbj7jpwUJmQWiSIjxA7kH+Ogi
36pm+JtGgn9DFBpzpCgHo642Z1lMDzpeMUbxc/QLayajX48Pd0WdWpU9IksSkgjN6q/tUXH+64Dk
5ie/8h/DLtAx70wMsPo1PU7m0y0QKQR25814wpMo0hwVKm7xaN9E/2OBGV8vY6L8DrWo1L9rYwsV
eEW1udDcHvvxEyFfYTJfsJu6hh1AeKuzYwgR4jBJuyemXehc8X1sPPNgwWAV/DnQPYc018aFldml
DXiiFva4YbiHZ8ik+DtMt6JW9YHEo8Rh8hv90q1YA1IFpRapcl6hWKtnxW0Us/IIcxgll7mr/+Ct
ApsNd8nSY6MZMFUkRmZsWoWk5mtUs9oj+dbshrtYg1C4torii4/vZKEmXw2WbEpXbeBs7HHEkQlU
hE7oRxLsaiqFoazVwSIeeJIlWm+Ks7IDrH7n1y3VLdaktxMlT+pzOKCtldOC0rQ/5zgtaWF7fyXt
QVTZZhoHMMQqUf8uadhXqflz2rwf/dntMQX125I1BNgLPOJYap4rNN8ynPowtCIgPsVVtzqqE8yH
/6Ml+k821L2/450WdnOweU8UIhHFjgBFfpZ37maMbuLcwq7qolWHjMOXITt0bwsvmzgb4+EsSpe0
HCdBya4GcWkWVq4tf72yNAHzWZaBr3795HFEVox/7Mmb0O1TjjcImHejk5OuN+9UyISvAvDcrUXs
K9x2ioR0xEeiLZi/T4kgETLmfMItCZ2Ku3AzoQMSxwxt6XCsIkNkK2lZhO6TWeR7iCLIdpWopYbC
mRQ30MSwCtGSh1HLl0Ur+UwTINHrzbPp4e4ygjEmp3EpqxO9/LeVDsw8AC4guQaDXHroFR9Dem5d
FwjNQCEr375RTfSQ00e5FgUVbUHuNzK72k9TpObD4e9wRJWZ1djqBrOKeZ5MwCSbfsstxFCQ3HeN
6ArTKVRNvI0HoHOO6LI7IuvOVPePH3P+9XvCblDIfr2iZNRnEHULP12F1TIZzZBaUVI3TAGsbDGG
S2bc2sy07XvSyGFXx1zQ+qtDlIhqpqzPZochTDsPNCvxb2cs1g0muK+yWJCLlgzjk2jGWMdIFYOT
0nVAm3q3Vy7C+9RkoNjGBMBASTYnUyCqUtRTrAGMP44Ga6hRTOyhGY1iBnAy3LPlJ6ByBfZxXPZb
GX7pMLY/YxJGcoLBIsy9iD8sm1yZ69wRcau8RVfwDe+6j9Btvs9WB836ubIMSQy0vHBJlGjhAn96
FlvnU9NTHsRIGoxtezXaGt+gHOJqO5bqiGK4d8BJmtw+3Ll+jRrizhTL5VYRzJELYvCiPWe+93Ze
yvK570wiQsww/irQeF8bMUsrs8IYCfbz+U9+00nCi0TCkKB1yOKBwsSLurDIHmkGaRzFUAICQKM/
czex7Fw5/AtMcEF+5Ctcgz1fEAc0/xMyEMG6xE2cQj89YR+aGijNsdmrpYn8Vbi9ks/fD8qean54
a8ahLnB+6sggYL0iuDYlM5LZbF8d1SZonFM5wJV+I0T1hcM1jFc6BcDBSfcKenDt8aVY1rDlHZVw
GjnFCLuW+i5GCJuYKqAiTv6QqGQ7XApGPosUfvT95olDqNpJjQrBhqFZuACS2npqhyakLaRHdZGN
HUGFGrSl3o/ApVwPUTtaAFlbtEnyO7614QuDZpurenAIkFZm4jWi78d8v9Uf6B9gNjbCQC1gwFjq
mm7Fnsk4qJAY/WHFJBWCZhmJsg3cXSsfX4u/HgQplJQ2WdvHdIzIDjrNSeRDTU+pJErQ/7qOt5rs
kyUxqb5X3xc1WNhNiUv6L6L5fL/91WNL3zo8KYKJM/VIWqdT6b07bx1bw8rBjCp20TiaZb5or2hw
0pBKci82KaUxkKDXeUYB+G8r+RmiG7aIBjlTxp6TVa09YYz0WlTuik8J58w8zjUO776Yky7j0/S6
+/662EEg6eUX5d7emADThIjJacK2FR15HNnNryw0CT3WNH+idUxr28Sij9cG6HgrmMRnEh/gZgQu
g8MswkcSFyhLUpHUxM1+gCwg8QbGLgqMgLbcixDkHELYpulNfxqz+FDA9ICwCDymX8x1zvZ8W9M8
kLlBf+2/EXMJzNQkEEl+jvFFoVwrm8CcYGJ+2FAXEvddIMvpAp2KATd00z8By/CBkM+aZJ1i7rBH
R2MhvF7fvgmbu4dPgvHGHnTvnkhWKrcEWufjLhCD8TX4aLZMsupyrznn3CtPoxH9QFfe9XfURf2a
nd5AUdbbEnaI26dlW5X73+Dx1kLEo6T+/89H3CaaLTiGfTrpfj+UKsIkykUwOjVGHzhH+bMp5jDE
jLyNFJtEEXx/MXqzsHyflVZTxNRVUfICxui9GQtksELXstMba+xTMG7NBQz/lcsgagRky3+7vtZq
aaWUh1kYmr3RhDLdaWTxsGllgXW2Dx3N0qqU60/CDQtArxCKKl/jD4L8/YCEI2n8ZhHHWqjv70gW
fQSnrQUtiNlULbPmW1H5x/0E3OtBHyTTHIXH4MLxyvw0dD+QtDrkUrcQcFitbp6/BvDKH50Yhc1T
puJ//JTjZVraFby0XWkNnWDfAEFKA7ZG6ulih+sSRnEZYoLIbvLZJry0Hf8ucgnKbTl/m2LBCdQa
XIXDHNflS00e24uMNywLGO2MPBdO/aYVv/JX7eMU34jv7K7vDmUQk/HN8trfLG93nFAwu8TtLp/g
88O6ndShn/Q7JF7ZJdNYfgiB66GONo59xWcbuuuoQRJkX10KQLr8xZqkFNahzw6lBgBBVqm3jKrF
29WMOiQDHAW3Bgv2e4SQv4oxFIkYXJG23PLaS5IY+lt4OY32i47HUcDN67n+xwAxRs9v1ZpYzT6z
eumvDnmApu3wpJZ1aSUeMaGHM+EsoyYGYQcFzIIv1pJ8x5HPDAQtxKYs+t3oSlP4trbvURKBOjAp
sWLy9iTFyjbwQTRk2n5jT8qjMteF7oA56zvqChI7aMbX4xqLDvxynzlTvnxY1d0WC1SYnoR9MbeI
cZmwa+KScuX9jYhY+9gw5/rCtkU8GmJtyXl+z7Q6nHIdZf6uGqPqOs4SWfTcK1V3LUEsoh7tcMyU
/gKX2hwnvndFOcUTRp7oCy/zvEnw3BzwMDjC/abzaibr01Wdo1ab0fDxfjCTjcKMUjzv/N1k+NBe
B/USgeFv/eqlspBlE6bFaewsvWm9/b/DGzyVhmZ1fLmOA6XDE9ozD7Q/iRuK6R/kFFwBt2TPc47Z
cQkklqCG6T9UTpNCKyjL2FUhqY49YGYxcpXuZaNOjZok9UN1xrFYvkIs29jeFJFR12aL6I+p0DzS
AojiIGEObmsYnygUEf+bsNMnLuGGAnfFOBaF77a8g+MS+Iql+/0kj5rxLDCwbw8uJqt9e4xkpLGd
ibCeUqXJSW3yWsY6tv4j8Vvyrf39keB0m4IeFj3Y6PJ0Bf1tvgh0CznpiHDxTmspwzvaeKqjWEf+
dTD/FErHfm+n5pxqOHgs/BrMnjnTfB2JLkYnD8zC0QJRnMmt4wyBQh7E21JOF+jLRO0BuvnaJtV9
EzrGAvWdYmaOWHbvYP4Y+9Twa34KM0BfBTGCyJhph0mUu4CmHX7TRQ6qK2FNa6t3cRf5Kh/h+UsM
hdjYajJvcQUB4BQHD3Z6ZWAEMRsKbEZeg2+OcLgwqWUXp8SK0UjtsagHrrgLbl64YAbKLYXK/x/e
DKU90oS9XYFGvW2UEjt0/k+XrKrQHzKVwFvB4VD+SYTHQQmFxlsgZzIzJDb/P06bitRkEH+X3AvM
jLIoAWyFGr3kxv3wQw+YfxEL3f/t2ZtLjeTEzDab3STDdgn8Lo8+z7I8O8tR6UTZ06SrQ57NKwmz
hRmFA/xcv3TUa7cB0x0Wq95hLZFA+t+UcC0xUeMH/yxOHJoILH1t5YU69PcWUgnaGE48/IaR+mTC
c82JgOV35YYuG2d084wGaSaY/li7oyW6g5eYSDu5xsMPaF7Cfw48Xh9OqQJv/YObXfBKzazQSMTw
kU8kyMvWs2gJ03ABR8wRwXhmhDOEQjGg1Hrv2ZZthS/db9SmwUnegjxAyXWXN5KpJfsP+faRTJS5
tp9LCQKRmoSR4mAaCc2d7hYGcRupwzB3fN7iMFM4UwPSpEJgoZZIdG6glJ7eAtwRlyDAdXAtYUCc
Wj7v/cYll1b2Gs0EXIMTdOVo9zPXErMfw2s44++apj1AIy8LNRI+1vkyboV4ynSwS6wsT429wBmp
OlELVv/O0P518Jn8M9t2uUryM31B2NS2iVoAKhjhtTGbjkre5OYgLw1jfGB6pQzx7vum9Wb1qYl6
RnVM8tjGbGzOLxcxDA+z/qGiRyvTmVuobsEtrUTCaeYP/f79gwK0siVJbgeEcC6iSziRbeNp5S79
j9X8tgl6hKeCE2mkOyFVvdktNL96M5uySWP5Mc72X0mt391Sq/1hx88D3nOaXQGBoA/b9PYDKc7i
9Yo4SKbeJORm/NeHLl8CsSE2TEumSkn0TZUnMK8z6EricAC9MZfUNMJ0IX4WHx0VXrjaUbJxRRyy
4sAdrm2ZwbzF9hGyevkgP/vPVni0Y+SItsdKGFxqtHTD36tagYSLIy7aiHu87TUaPsUmJ7n/vU2X
r27klH78b7ek+zuhU7vkZ0iNy+1HgAy1mVn+8e4kdzOXZEbqi6Ao1n1i5Vop1v6v9O9NQhe5x09D
fAtdUjwPahAt+OZu1dWmHaxsc5OGb6B0CbKzKpxknPfLymYmUGGaoBdlsMKhmQr0CM0OE5Yn1/Ww
GB4du97RxlJasQfLOHrSkkEm2DsMyItiV1SDBzwicaZsa450VOdKeiXnJSydjz4dIZRbZYIsTFo9
ycMhPLKR+YymkU6f0idfWT7c6SqwJicQIzkOnS7wclxOzBGZ5ozMzKjX8PzzsqHj+8rvm1sKQ56P
SFTrh6CIaoJPANHgmcBnW8x4KngLl9j7YzylbCI3aYn92DMeQpZF71FnZXRjhGvPqLM5dKhJNR/L
S4ZAJkkVbcj8IkhibYdba7ctax5SXWwaPFwvYFPDE5iH9NT/Atuxi2K6JhOqpsmsmX1qGGDjxWlO
Kt6tCJsPZdVRWEI9IRgNq2/0yryIsNCRoa9XGssixwP1xyXo4LpJOKiRYDhD7Eoo/p7ohEMNK9Sc
WeElMt+eCSVo9hE4kTqY+PO8chMsyJUD8OOCjF8RpoU7qbTWAfMZi3hppt6mJlbmRKSaj5AWgt9+
i+uqybfDq89SFN8aq4uuz2XVvIW93S2NuxEDiCvqtRIZW05OgeMH9F727/ehfD4TivnxL2F2nI9I
1jlF1g5j4maqR5ocyr5GdPhHa+/rINMKqSsuEiG1HvP1XUYFVvZGbBMEy+J/DfEWQnJktXagCQy2
6doeuP3RTb1otiBOAra44BXypODczR+sSlF5tbGww1NcgSSnW6CYfR960WyMf8ZrM7OAB6U6SOOv
kONEy4AMR18V/Xf3+LHW6A0+k7Xtt66cr48CZM5RMKxUvKdggYuIrtEDhOJw3phN/RuMamzfaMpU
Dw5PPwOIVVMtBgSiFQPUb+e4Irdm2tch2WSoCs9/xpM7q4MJcPWDcS1OKYQG3dtpAYfqHmoh7Gsn
3Zoyz6nlKl23FUwh3I/9xe/S9lgqarsXyKBkU2o9vOrcDAZZZ4qfhwvg7/QVtGphOSW+MYFQfST+
6qYEOpQI7ds9eN7ogZrUNFBIIzq8KHKUYFBTIuB8NymEIy33I5ClfIPB9Mm0uI51Pa6+L79X2Jcm
N+dUYBLkXqdY9hb4FdmM3lfdBhTnAT/C8sUi0dRQcaOqg50RtnDpqIfVNuEUeJ0FIPRdmR4ofgRC
X7Ml42KVHMMlE+3kMUsfvi9FGqxHYMVZgGAN2LImO+8eNfAMBM3+k8wN5PQyJ2h6OF5sFTuNelSh
Gg7Tm5LFCJlhCX3IXnuenD6sBfslN2WEMe39BwRpHddJFczBS3vjauAAfthj8T4qPO6IIte6fAil
l/w8xGGOu1LyTRmkLiV3+FRjb3RXRDu9eJu7Fp/Ya9s3/Yr6E4xhOpde/tz5hInQTMHHGfOiZfNR
JllCJv1hdSBc7g+nqzqrYx0M/HjxJRPmr7Dy/lq0mRboA/lXuSIij9lnFZZHdKEMw/GR5Es6YIU5
jzmA0VDPkY0wdVpTrS18abhNtMstsE3MNX6TGYBh+ROnp+U7oQDda6suOxRaq73/AUXvmbWUi1jM
hu+681MA/d6VCmFYqGJhzRjhUjlfv0J2toVw82ampAMVUeqe0iPQiUrpZJotC3HE+Z0JHZ1aLwkU
4w+aiAGDvY4Lqm6quGzW+2vNU6gm7uvnAziNxbD+UTet+hrgq86d5/SCecljsW+ALmg3VPSSRdv0
zbSLZE4hxCowjom+dAo35ipmDsW8bdOj99AX1VB68yMdbVvTV3lKuqAMTOQ/3ObKR4tZeIdxsKPd
6EgK/TUz/PJQqQmWoYh56vNsJ6TLc08dad02SqDGuVb0CG3648PicyuA7cZwTesiYeiEixbN5jzh
k4NyvkJUR0/A/RnPLmsVIVd/yGsR7H/kSCHVslGYIJ8uX9w1oa+tBQtNQPruzm7v4n6C61ipvRyc
N1nkeXgUZRUD4zpfiheAxP5kpNdVoklUpi69u3naGPwuyjbWY2SNwrMBLiydJD80KX8StqF8aN0y
LSFu2DckD77IU24lbSc6uCRmnl5HuVg3/taTsXaXIeKANm3YiJk7EcBEeEatGgHqfyysHYu48/2T
EqLvy2T+VJk4afie8VWyho8ERxM1tvnZwYngUFW4gUMiw+5vbIbRHC1Kgfm2AEGv9Zt1XOtb8Pb1
mNfFmZKMsRrbOjkWBVbgiVpe1vNvclQm7TlPlYbEtRr6BY3PuEsR5U7SaoDM/I2rMHZF2Mtu2A6T
iEMmj3elzAdSNhTR2a3j2ZPp/TCh43I/x8TkSHsYRMb139Q/+GkVrMK2oqud7aMDa1AzoWiPbvwW
GxmZviFwmV+Q0XCj0VtXjDET9iacholJai/HExAuyFi3XV/sDq3wj7yLyjeNxTPNfC6UT9m3cS/D
FIefv9ZCK5KJflaJ4fcHK8WzLm+NCFN9V0hkiP/fMckRU/E2HRAZErWoMoS9GIJxGknEk9nNSHlw
+6LgFmZmiySe0GRPkGsSTzFgtNwM+35tzkt29u7rnVzQC79CFnTssZp++rlIboagwNFoL3nxOOFT
acxKA6MMhmalfX+vFAjgbGajRGOobQ+XXJPEI2/20g1j8QAyRqLwNMpDjDF6uL9P6+Dh6VMPIRn1
Socgcy6A72wPzIL66Irz0TbIcqSOkCpeqB99ow235O9yvQEXfGXYsTvEoZlVb2YGUAQNpuZOCOlS
PCXyarBxCCPDs/vYJ6dgvWyxrF+738BfpqwWpp++ed9ZxOV/3/gg/8jSgj8icVsYqJ50jZk4DmPT
yBVsFqKrgfYmN7B2Ts3mOjYBBwgT9MQbXy7wyHrlwfXlRwWCGToMghqPjvpEyQ4+IcKGYtHjFrEA
PSo+tjGnw3a/mXCh10ixqhVoXdry28o55qSvdQ/ieo0K9tSUraK8s5uQlOjOZ8VZ+CKyttEsy6rd
Vy5r/I+afnCEFc+PEi9+LYF58YIUTnfqojx0zW4TrK99ocewaqRcH1KUgAOFYJqrhpZA1v4PKsIA
T+Lcdoc2OFnHkzGEp5+3LMnsOQWEAtS3JaySvT3ZBaAHr+OnvvtwVxVKg1gIH99554d2g6sPhYo3
HA/MT7Vf+JyGw8wt/lJm+SM/dv6KLBllHpqwYkJs8t9ad0zw5wC1R3tEcnvCydcEPT/7CFFJgUW1
kGtV8UzZEiO0jM+8YXmgnqFx5oX72SzT+F7MPqZifT/lowZiVv0cCNRFHJ6y0VTnZOPPD74okDrs
MzSv+khWuFWsGpYKm5/Wluzezb8IbVL8iRjHBnTy46xoQ5eygT51q4Dlw/FL59rSlXMTacDq2dH6
y55luXWDWd0qjQ2LXpXFbUZlSABtXYfrol6KyVgi3jW7nyOW7Z9JmL2t2kStW0luK8XWsYl719FC
w5H4pr7w/LzRcqNu8vn0TfeDH90EaUjtFkCAYqwd8H2+7EMh9/LVz2JpeQnOqK0TYbNi8k99Rkru
5NbbPJ1T2ehw4CJb/3znk0xLPjpp8bX9NH9Z4ZH8oFcXhZp5t3Ns8KiAgheN1fxhG5oahyB6LhC+
oEbWkPmqjdm4vxmz7jGBXO4JPuHTJrLkijDeEQLs6p5f+i5MjZgczqTLUk7OKLwnZlC7ceMbTIvC
YfQDsykiOb5RAXdG8tPRks1lysNMUK0OGxBzVFXa1hEJTaA+/S6Yko7TOERB4pc7X16ftv8zPXQ2
QGc19lisd1KR2s2gILduTHjKpObfqH+TPEynsAydJr8BNqQSlpiHprvd2mh0ML5EZgTbegCDiQLS
A7IQ8loVkAxCxyB95wdYpC1gR1FTw5Hxi8yngi8ZvP4mt6s56BEgl/ZjKzmIZIWXlKANXKtqMEJo
l5xk1hhb8tW2m1WW5ZvZSFnuEi4TNRDJeBFHUh+vwJzGaQbtZbE1broynGqQy60DeUPlypL+sxle
HK4TbyUf0wmoYogYTmHGxjWhr6zXmpmdd2sgxVS5v7yEpuyh/+E6/WsL5iI/2kmDuTxnft6zSOrL
HBmlqFnQFAkw+KacP2+++XAX2KBQvFA6CgHZz7v/kSED4FKqLvcJOLScmWtLZ2ZBlshcJml/jThd
8Y1avPIrOF8sZfGy7MQwS6MO8lDzkBIUM2/7pbstjHeUhHemkpu7hDke+IAl0ruOI9bXFhn69l77
5ETKISLlmaG+za97w0u+pP7bGpNaOtIkzKQ4V/Atq7XVIfvPYg/PG6W4ymIaJRWyB4SNZt/2ZjpE
7vD7H51sx1r39hnKXbO2YdCt1q21GakdMDmQvYxtJK8iyWb9bCpoIT0u89d6oA+Qzh9OVP9brSaU
iCYq63gcVAyO6m03UjWP1igNYdYGUkgAdHamvmHS7jCyjHsIrW+YnW+5aGK3pkf/4gDP9h5Tw9On
p7+esy1+7iOP2ow2cR/b+3uvT0nHYdlVrTTXCfkUd7T+yH+YiTmzE+jfU95x6Wc9t+5GbKCsoQAS
wazzCvUVScn/MGHOyqrmX+oyrK4up2mRMlz6fYtl0ItKCmUPDJMagqFw00H8EMxNItlwN/eoA8NX
0AqhEvgnrpoPDcGO2W6Ozw0F+jMumoaeQ2wknwlygX8uvM2AaJO2DDRtjSFW5BLLhD55j3bUs7MA
l1b4WkIQL1i236JnUAWCf+Y1eFFHjQ5Yy125b2RZ6JQICA3jBIDFKJpNKAcXEg3uabzqq/rQBCZP
W3kGGcUXHR2BAVPP9roqa/iVlgPlQ3qqYB5F+2QeYXtt4KVSIP+dUNheX4730J3AdQlNYnEVurh+
BfYSlU/Cc0D8nAKAkPE2mtFfSxuHh/bNozxNjxf3Qc3XA4VtIHgu+eRF3n8RJijc8t5eaT9GfPON
htZvask1Ecw2jPa1Yew8gMqIFwW15jbhsS1+4x0n/obKs2pDkWbAdwmMPrqcd51J2zf6H6dc3zH+
2QplsgcIH1j2I0ZdusNBXTpZVLK5Qiy55ItkO/y1ksRRiz+Kp29MFS/VNU6ZXA/bggefLko1CjPQ
kWunfkEUkmZ0iCQFkZRof/e6lawpoX30xn5vKGV2hCnEeQPOfhkmiMiZMwIswPn6WRdzr9mzznIB
4N8wq1H/KGYKCwVlZWWnikdAeS7R8uYG4Knjs+zPqqncI0vwOkUAEQXAZBX9INWAOFfq5s7sDcVg
HjzZS6NdXfyK6zgl5SYyCjfztiFIq5Bvpy5J5KPet2zog/XPfaFdqbbxoF6AKFSCxU+8At2+L4Ir
ihovjh+mVbIaTIoaFO57TAxvkNcG159s4eRpW7Yy+F0dpthuSO5wgk6IFiu9B0PQEreiWt2J6g3G
jEQNSoknl5KAH+Zm7T6Qtrzu3fFXv5TOO55QDun1APn9SKwf8HtAxC9GS64EMpZ6y7ZpL71nt4Mk
yEO2jbF/vQ5EHDtDBS5F6eGDVwPBkk+ekDMBpY2XFdZyJfnSwjdZIKJE7zhfNdsZvYyon1qKvx4E
QI+HekPX+99W3XV5XgwAowivp3Ykx2CnW/3lZFCNo1Pu/XfRpCD2MmhvJ6sfeU9vlKdXUo/zNxIM
4YXD+ElAuIKlyO4Nb43UFXc2yVWHQudfxisJzTx8NWXD9I9dFnEswIexHprkMYTxgNADLJnN0lmP
LGImZjAOx1yZbzUZjHf4C977Zug5dp93S+g5oPeWbM1wWwUSRb+peifM/zcmVsqunj2EKULMXAFh
gzBkJhyv+8dD/u8mx8t554pkz+I4B5cUM/v+02QieVNYLPSjiTc0L0ODUAvVLi8xEhlCUVe4nG4O
OAD0B3AJKzQ0Bl1P0Hu7M8s1HmsLuaSDRe9+tW0FQ38f4bWhbEWtb250iJUiMsmJU4wRN1mFszX1
tO7z7ahno0/cYeR6Qzy7xFIAvo0bGDVBJUKBeEFpiPYORx9XNt1sCPgw14xPiL1IRBTocgrgrjsX
VPH1LxtW0VGn0s7p0EO/UyfEoLlAIx1QkV4n/zVqCHf/517np855TtjAXJhlTZqiUDTpkGFQiGW8
ugCXPYj4hvE+/3c4UpAQMTt5SG3qEYWICiM1mhkrtzI41cmJEkB/UQISrgQvsA43TnqfgGsvuXxn
tTVzTbCkfkKTMYC7ClGyb42pzl69s7BJ6ncSsqbXaI3z/IuimB1yAa+cUDytR3+oe1tzne399oHv
knxDnsMr75OuiJ71w1Vp6TnPqKUBgzmmjSb797RQVaiF28s4LuPABjFmCtTzTOOihmspROz2t9hq
y7Z1CUytqhllesBix2VnlIXcmNSVlSgrqxGl8Zrlp/641tnzs0beK0UjnmWr7cejoFAfd6AxTcxg
m3jF2UMolM7LIctsZg9d5zub+7snE/ZCgQT2azt0O0bt39mjRO0OqLq9Zg/vvaDm4QIux8qb9sjY
TkycScjCin0ReI93nbx4hBNR5y9/knHgAMDIYZW6NZ6KCWoj0i4VGwjUNbduYUQCy8QlflDDuqrv
PPfWbaqgfwhD+wLK8dmKQAneywYXIcB7daVUY03AN+Fp4Q3VxUhilExCgnOV4064WaNVZNSBFX6J
bbMvo7N/OW/JL/0Mlituy4f7MMc9LqW7cLCKZCaCHpmhEv0HwrBHYRWfxRPAZecXtcqqRwnnQhdJ
pGWvWBhgNAqLfZ7SgS06ZqqjEQI7i1dByGdrMVE0gi3nIxvp7KYrnaN2qBQw4tLr1zzXb5l+alQI
M03BFVfv6rWZZgy45i5/mTUUSLTCOA7TEA30hgoZPYr4hfGgR/RPOohmCvst5KPXcLDRzAz4pgOC
kT6zr8txiZ0hQQZIS4AJy8wb7ykW/GdSh3cL5GcCTBDUamizP0gqRfH67lL2tqTV0DSYqqbGgg2n
mlaGvBu4zTOp8SVWgf3bsDcykvfq9L21ToQjUIA/5uO66xI4z5I+ao3NoGQzPfaboLS4+jXXWmsf
pMJHc0KuXR98ss8YxePrlzht14GBmwo+6COeTZbbzeELxkBJnbpbJMpUFSkyhO81T3CkkFlcyoG+
HTM2pUfYf5BFBrwQumUWEAuTGD1mGEHGwLtxVDJyQsO/Z9a+UcZa5WseRRtrMMGXz9+bWmsLc7Vz
xZdiEmY3+rk3RwvRjvOOBjMdZ6a6B++r2FM5LgaD7j87GQ02rGO8ZaH2d02vrzkFMPyoJklSw9NH
PvWDDxW6/zKtKwArlc0E/SrpY+96Onl2ysjIauZN0R3z/tVnh6rlYo2PTBKUAu0GOYncxhQfTDVv
gKpzCSDaI1/YhQ0BXwNpm1M9zfHrVNsuSTHW2Ouk7Wap2ZTYCoqtOP20a9rAim/9dCfuRea/+9I2
vRkOmBtfAsa01y4Zz6+xM3HnGhC5bVf3ciZkSREjPSmbPdCZEQZLdGyQNyILy0SCzbu0vhrst51z
Hc4NYbCgoGu+jNcPoZJmsGAb6fHQ+XFFn2QL8H5eQ6cf5JP1I+qjvc19TEFNU732t7Sisd72MX1d
BTVtLF4lF/FYGQE8PBKO5wWGGpMIdOqTQ3PfXyNTGqI9m6EQaylcm/a9GqJNLo59AZU62YHEv4aJ
v62ZW0iQiEfgsLJXmegZqvF4v2jIzor6QGgrMSSDzhv4YqUAWctR5njtUStjCp+CVlUl4RhMFS1f
2TLANTujJoztJGSAhnjId0/oGbYmrjy3eDyTGMDJV/7Yxb5YJP0EtD/kmfukRjJJB6uI9hgokZui
E9WYd4dAtEBuXkNpmjbWCSxSOytB0GtzbXqj+fX70QQkg5NqYC0n1MANw6W9FV3PPxMi2lQPLPyU
5Rdp1fsGyLw2pV5QCtFwBO4jT6xlLjIOtX5ZVOkKlk0uh5AEFEZYtMVNZhc4C6I+/LLaq/DbYoPY
OcfnemIDWGkBVhMojNHcczMrSbUi5VidoTizSwzo5Cts8LkEiyowVp3S5bkgcEFzw3OUa9WTSLGA
fZ9z3Jj6cUFkJ6m9OGGXEmlMp7ej49FpsugKnCDYbyttTpMVZsjJtSfLYFqh85/+/LCu0KFemNm8
KuiIFmziWzIwQTtEu6hUzj8l0+AdGMr3e97zecN2VM2pvgKBnWc69h41x0faGijiFygMsZvAguDR
1HIpHZMCfaJa0IeuvLLf5UahgiQE1nFH2VIjy2hCi1dhmtCROQQZPntI213/npDFMztX17T3G+Vm
92oHiWmm36BQEXaS4v5wlxkA8SpLrxpFwm1giSQlMYOy9Wd7S9JAfSnORHWNOASljN+unqm+VUX6
0BC6KTHrN113ACP7d8nInFxdjYbb1jWyYQQxzaDT9PZl/FGnnkO0Ru0s6g6wZU77uMjLiCe9Wbtv
fgNCA5eP7HIx9/MghKjo+28xq96dMXGfqW4x+Q9e1YD3aTWXkSSxZXebspQ2EVRqEBdYFGoPimiD
1Sx3WCJn5H5/GSb5mLzkyHER4rTJ6fSsO0JcK6JBW9DDXwX3F9rqhzNcsrSh2tgFXC5jaM/ECdFd
fJlbw2mkGR6jUHDVz+VSb8HA0R9SaiXtXD5v39zfiAztkMpPqelURjlbAjacJx9I1qwuZ2MnVuM/
dCbMZfquLgh0MqdrrM4p2dpcxNtkwlfLHUtujHRaueNW3pxiIXncqyweQY1txlJN7SrjIIfHS1+D
Lde4sMQ4YsDF3pieEL9eJkHNGw1/ZHWDZ8kOHfOhcbG8CiJy94z1Mww8oH6zm1e5uZEm5VDSzAMj
0uLEEwPda2eFvvVJM1PkVoa91i+gRXvUF4o1Y8SD9wjR2rj4HXG8YUYnyYMQULzj6kfOaDhRvimW
K8fM/1Q2nrk6G2Ayc3Lhqt0Qd2jagccxoRFw/A/OqwkC68a6DTo72eMkEWgNiHYvlxb10ktLk7Ua
P2TaeBHjxlqJIedR7xofOq0HHQBA/v/wFNhRGUoLs3hReSiJqhY9X4WY3LyKfJBmFvXKI5UjPbp3
tz+c0/OkJ5vjKofnxUWSzbFjlAurh3lhWuN33ZfwsvIT/kjcaa0CmZMBiJgZMoNE8DEfcnlnIhWo
FR1A/h5KJxmScA8KKkheejDDA707quui6ODSLyUlZKt4O1ShPK8Gt3K2pMuWRLjHx3xFXDKtgXCg
zmhGA3CqRq37aLeww/lG7//s0cxjdlY2ijl6Tks02i51TnFU7lSle4AiPEQPKQvvnS0z8mpE3rhi
zuwWreAlYMEmf+cuEAmlTVp+k6VRROQ5SBbbMNv9WnhdfoKBIOb3GlF/TnGOIkeBQ98iK+51su2a
91MG3PeAbecIt+PDfz+ZlmvAHdbkapy957BGO8mypiS4enuHxi86R5G6opCpJGS7zBev1hxy/Tvg
2pINfRwUN4M8EEFAN37yvqjBoQn/hx2+zOFIutLiiyPv5JOU+HuvGu51NT4NJCtAwpMO+cVijHaS
l0vK7LmW6Vr/iwBzEC7kZ+MFjV3ATEFVblmwv4opr4yXAuIijlqOR0BLJ82EC2zhA0ePjkIy0xJO
ji5IIWbzljocQwdTrg20xKtT+oD/q7yXxjK3LonAVMGJBWG2dX1IVfsl5OgVbHZ/JVQO3h8noJby
71P3rjliTevElmKSRkusXw9+6ZBT71Kx6fff8L/tyCfRkfwRCLWScVmKMnDzTGoDGZm7+BZIa6ga
wMNYfXun9BNoko//6XEB+arRbcs4A7bPgxpEMAM3D7A6ZKIEjtnaa68UgbCkIyoefCYJXkF0EIJE
vM5Rk59QbU5Pvb+8zbdzaomph2zhGI3Zspjk4Q6p2BqBUIMBsFLq6MH8NT406dpnxpWhlUO6zeO3
kIZ/foBgjoMrwY+Uol9FzEMjb6ihwJ9nED00ak2JEZQFuSnPYSOLZIaIn+1KGcUQUXkpqHWTdCIK
8AoeycQVGHTk08nvppSx0Rhube7Gj3d4iiWY3ZMScu/gSqQ9V/nPQ48oNNUYBj4G3yxVfl90m3GF
f6//mwoKR/oOzHK6R5hYqfPoLYbQxmSWieo1rdCFANZ+BA/Fuj793Hlfe3EDFVX2PC9jZnxwl/WM
MfsWUTxMf1F/uQ1ujCNYcPAeyTqG/hef8Ikgf1zorYRtwadUd4AXheKbXE9hKqUbIJ3QJoUM/vXb
VnZuLSHvzss+7CO8hk9khntYE/Pqhdv2xIKRPNyFOY00fvOMACBDu4/ipSrKxuNhKAqVaNUZBpHC
ywTZPlBEWaoPBt7icck9ZP6aQWNBrpTUk5657A8xj0kW1Vs9aKTTM0V7Hz8ZnEDfX9+67zVCP8xk
dU9nk9AwKdBzG5hru7c8lEVLMugo7V9eC8/ZZ9ucq8G+lOxUugFhg2jh5xVofseOtkNNmZplepyF
AwMgAf4jBp9LW05k5ovOUvdFsPrV4dSVkYg9vC4L8q2HgIGFBLN60Xm4XjEf1VDRRp3UwOwa58IT
+OyIUmaAgHV2K55YEMQcJYXS15pGvGBWi8Q5CiSdSg+W0biuoAekxbHA6NgT/UFb5YG5FeIU4BLb
XOUw1G3uX5AYMRdttHI6WsR4FUZBt9eZ4jwYyyIOcyy1qkxZB6DAZJpHMifR1KS/9SGlnAB7RXs4
G3YzGVSTiEHAK5SejVlKf3fO8MgrOGFD9zbVHtUVgSkzWllOHthR0i0g/99taqPX/KIP9Gs7v182
xj5h4EaCrULVhx006RuKaltMDHfSaNTAabrIpfKIJDbRTiV2zRW7fRpKS1EnG8Sjl9NxNvtFDGQr
+6gyWhnMXBCHiYO506kjZbdAj6YnVJP4sBWmvTVD31dIbkDXE7lM6lSiMjitXqO2AtPqowYW8yjh
zkoELkqCCWWKvyWN32LBGP1L/dlFg4lbmoBr6t/hGSH/lRCHjrAV0h8+W1kZc3RqOSm8dcLk9rXY
+L+VhQ3AbdwTYYZ+n6YbbPpuuh4HF/Ygrz+eX0Ff561sAzqVE+r0THeCiPeQq5BBgvIxUQ0jMScf
0g67mbaASr+c8vwOUTY8H2W4L1J2DC4Enm3qjiwLlvSl0puiyNfzHSYgfelPUyVAHl7ZBMQ42cM5
q5ZL6h+0bN06Vp5Qz8wasNZmRb2JvbuCGb/o9udHUlLQc0UX/bdSjfAXe/oueB9QvOhpgnjM3sC8
6BM74nno+mhJVIQ0kuJpdVxPuuhZsujFHHj/RJeZhVaTamR4A/QBhL6gbl9v1UryAzpjpar7fAm4
ZBnWuxMxQHH6ymx4nFJVHJSq2Khl+bE+j2HgIXpHo9OUkvqxLezHSIuEAVxDsJouWFBkLKshAPJ2
ypFcdBqtlc7P2P7o2C/vFHgUWA2bQn/1P+xXbl17X49/QiridKXSOPfGBf4TLx+IktA3Ufz5JW6n
Gp3uaW+gflCU2azM2Bmn2Eul0vG2uLym+Cac6/dbs3/tLKoCWnDDdJKNLlIc3XndGlMJVR528NQZ
jvLEacUYsuClQiionubvHQvAmmBBVqeihtyiwEnGvX/Bv29L+Y2UO8z07Gq+0lasUb/SrNZrqC/o
N5Ghd/0rG84WNMb4TDKo4bq8ucKX/omAO1mkStRdQKwqdnmN3vv65mbTGmPFCVZdGFdGD8M8iOLs
ALXul5elXs4NnG7zPpDoKHo0Tm55YcDs3y1G5I6wLlTaNgNsHXQmnbtg9p8OIWVgKEFVABMwAQ5b
hKTNg83YFLJXgwc0x98vPw9/0iAQo9LNRuC4QVog1csKocOAUYtfsGBRea0qP+EMH1lA7te/L79Z
9EeAKdHfDY1TsLl70nUeAsHR7xCK5w4vREtKUCobyumA6dy4rrAaBlbu+EdRH6VDeajG8OOA95iz
OZ+v6oO6eAPovmmBeODcpjwKQpSaui0anKFSTDC2Tf1w0BL4ENDRV//vmkizCHhvGHIpP9khegIm
+jqrPQcTueqkKhAF3OndemxeBJLYSgcCCQpLIDe6VgOwwPJuQ/De+HP/ioEWCIhg90jTR6Wrkcso
3CCq3wxyXGZYOP7LWfJJ8VYA4JC8koYr3mldaXmf3yXWOLTc/nfRO1LJQNo9PykWvjmZ0vcmWi6K
O1bIM4rdK+ZtQuG1mfwvWCMVXrugChU6rwVy+/T7sRCAf+q+WW37vxNON213MKZHGEpP1Wup+ndh
2jy5Va0Ju8Kt0UBFZRFFfbbfQp07JTB0vAj8bV+HvPbCthPPVNc+Iz46u2zYuq427VotuKEIAJwV
2mTFDDxWjNo67b/TQG4xogEe+dehu64UmDbX1CTmFQ8Yd6ljFlmXsYBkDuiAxtUTjF8cqX1VsbHL
yOcM79hHud1yxwmOlWZw2v8cI0DTk+BLHPLFHAkQPT+8+PUqHhZNqiu2MoPWfIBZ1l4Rh/UsDJg1
58Dhp77YsvUnfhlI63wQhblFsKnNDAVTLyyP1poq0Uq6/JrmQ9NZI+bXwXhpRHqrqAa92+228HEW
xEvy6JrRWrI453bleLZdFkt7w1+pTXQ+G0tV6TgQiwt9q2nFtfTGTJNzZ9XWSVLPrlJ/WGeYuGm4
LWF+nVgRMtTBGMcg52I/BnWUdTbl4izbIc4d0eQXNYzr/YI0BQCiGZ50o5npf3lGGoDZ8ihi8v12
cwS0b9e+itF+RmImzqcPIU8ynIXHgNzFFXxesRODQAiozJFdN9wK2lq9sMQhsG74uwOdIqufXIKX
f730oXUCQB44z0qWF8/LKox5yrPkGnMYmijYt1fq4MlKYxw5qQnZfGyhG3Wd1lCwnyV/hfQwjGaT
yQZT3gw3eNOsNtieWOs08ciezbk/1JnIpHmfmCFsSzfRMoFY1xyr0wRJGrK2+329zV1TTdM0tOw2
+evNUAeYnfriy6+8kjFM1cBnwOLzJbFOB47nxtyUl4vVtQ8DVJft5aVLKLtFZBKe7Gk7DiLxpD/L
m9AYsr6+hNCcS05wwvEcDAw1vWW0x/+kASYZGb5K0cdAJ01dOlwSDqJqyr3aCKNDCG+H6czCtbK6
zDGnUzxlnYPWEhgRUs5OO+UOGinGhTXIZJW8yOrTOvS5RVCewx3DeiMY/Si5r6R1hw2wmcO8W4rK
2HQ7nNMEcN0fV/nV4VOPf7CK0VRfoKT+VODlBUNdqhRCaDFMHI2hpo1WNx5PxyE0zrsyld6+68WY
pU2bVT5EnEupF2AwUExzqSP/wm1H4/7D2EkHZiQ6S6jJ/Dr18koEUEkIVT05S6Ml9s4aSVm7dJ2V
BbpPQHpfMeylnbx6AOzy+YYnMIjW51tbdKVdsEYHZVhHGnnXNtauK+FRxFuaVZMcFPTf6YQ1getR
21HKvRj1CD60ptmdZERXd/n5qautyaIRRVs+aU68OWdMD3Gd2N+5BF+/ONnoR4CsRSZ5D0qFiOcw
x+QM0ceUx7Iv+cHC67Qck7HPOxd5ZZFznrEuM4J08Q3Q84MTm51wplNCuQAPqAKJhewwwbtBkUF0
ZRzl9GrRRBf5I59rxA95HDUnzhQvQMnBsMliRR6JXnpJ7FDD0huFfZRqsRPtpNHyOwFnxAp6qppm
ZqYtr1euqly/ieKHznacTm+ca9hIDE8tNPq4+cWrLJBCsPEVF21hSosqbbupDhgi8m3JkN0Kyl9r
vOzPgKrlt5VD0V3+3tUGnYs1jCHO/rGvrLFHMScEf8b+kHoiICg0GxNW+zIyzMdE/btNZxAcpKhD
cgqxd83wCMNoR2Rf1G3LzVC8u0dTtROKAHeuhborfBOev6Hlr0hIEP68BqOu300IHng+jZQ9AJvL
0JHYCGjqfdOYd4SbBrzdWGDzYwZBxSdes6sHhDdozM/8tl5JFNl5oNwypgnd+pTmCsIIElZKQHYC
KsZvXLhdhInsuFRi/YZ8Nd3aoZm1HLPWv1DnDU/b2v4ijRUZCfQiTIud00pX07ic9H0hK7hQxITG
o9TLXli5UuKQYpgataGqMPWcTBCathcwDnMg4DfvnGTsjSSDOg0bGTpVsm3Gv15jEAyLSJzmui18
cvRAY0xANYrNlYgH47w4iKUxMwXWMI9Fw8CWFAycteNrwVsOO20YS4L1MeWgpc6ugNyCF3wsqYbv
1+3gtmbN4kS05oRmm3ni5IdG/M9+zl7RVsiqWPe/0DPR7ZGp3qrpCNgX9qGVLzzyqbKf+l7TBJq0
Gwg9+teWu6nlvpUBjCfnL0iEaBIwc9oEBXULwLuU54f9Px/vRc8PFvNZXl9N2sjQV3AeqyNDYMgH
DWJi4wcd+4U57xTh/eufEF3brgniH7bpo92W3hy3bVMKy3lww4N/kRmeMxcaQCawCyBSe2tPMuf0
qTr8YQVTKUkpP/s7aoeBAbEoA9M5AJRuf8SVl4S4LlBOOYLxp/Nc9gworaj8UbdzeN6IWwC/ii4+
w9UMPeLk3sAdaITjKo/yYAtFqFtoXUyNn2OcBhsjjQCvsspxDhxWPAiEgN9UWbqHnP2IS4Yqn483
41Cig6Q4b5vigLYKQC9UDFvy0+00XCFPDnJ6wVMmeknYu28SWqOLdGsyMUco0Zj26QZ8KH32Ac4J
GfiZ/+e0wmSLUv3mHzJHuJR4427WKQM8yGx49z/hdUpm2C1yPxBIIT8VpxEiYj9o7ZoBl0WW1Mvz
o/7xuGbPWPVvJ8P0Sm2y4jMotg2CnrN45687LbTspvT18XDcLyWpgh2F5/ixBbYitbEMwEgAvsV6
2lKch5lwD86Q4lSW/MwiO+2wKCRfP0jKSq5PV7bscdf44qicI7y4UAEQOG9f0vlVjcPrMt6vMwmw
6TIs5RMzeGUUUHl3UtATv5i8yoNR0tPEXHyxAhRFgalRSUzrGXLTCulgIevdUgUI+KQvHbZs4lO1
BCKzH9lz9Sad10j3A16mbnTWbH+fY+1QU3gV5MMylluMhEJvrjsGzPDc1Remh3Sg2bT1dTs7FqOP
fSCLrkFxEtPkukAGQYjgU57JFBXEX8VizjJocjZ/ebc+Frl3jES9tVk4lp448S5TVR1lIuyBBD6n
tKmAZp6tA7Jtew0JoS4ADN1PIMHJMvQFMRjB+icCKhnS27wEOdoskqv/MiU4gOE0QpTip2ZZVSpf
JUDxFeGoqpRhOPSZeOOaqWMUjG0yVjlkCxWVj/jGEDBpQY3h4Hv0tOaKgd0lgFh13ZJ+Uh0gx03o
BTJB3DAFRDpdpVnfisTOdpk0/lECnhlvvO9r8DEA+pB1WD1aaUH8QCfg0LHthu6KtReN5M3k0f0Q
lWFTvvIbGCjuiVc07WYGZqMnM4Ja5IS2yl9VpgH9YbmzopRcY7Lrqsb35L+4gGHXEimSWRhD7m5u
9VNSwek/JeYe9x7ltWOypXzz3oDkbNLj8cFwyNrccBoi/jBAnwdw/vCyV9AB/d0K9Pwl1YlWrwu+
BZIvx00Vu1vE1Tn8drkmu60QjlyFo1ALZbIddHmMSOWLIhxZ1woyabH3ejX6afOtES3pB8AnxDwU
YdtPWS1vERyF3qGR74j+lePONPsMdzMicgqGRPicipeQOB+84/tTR8Qo36ndMomYMSin0u4l/Wiz
YmMJk6tdEN9x631Ttg5e5TWLu+YHZefK7cCHIGCMTfygXHpkK6GxOoEssA3RUzhqE7k23gObPVSc
HT2Ne7MNYS/ABPa+1vnqEpiPi/lg8Xn8APHprkNp6r/nbS/IoAORPtu456PRLBi8L6P35cbT3sB1
sKoA8R90LOwR4E3VTEDrSsrJoyAEe25z7JjWhjBAHE+3Z2kKlpSEDsOP/ny1qjyCZiLLG2twl2JO
yjKFzCrhK7dHn61ubNI9Tvfc4LtK5gcED/Xp99kmhw/wf4DScK0QmkuvfgvHYnlqJZ7OQbb4Q+RG
nFfofQ2qVjJyImXU+4fyeSU3m70KA3GSb5OD1nxf1YH6VqjFzOSdhxfiJRlv3kCWjdjlDlbwvijs
Bh3KVQdJs/64p1qJcNqV4f4pQufmrSjlLUNMtiCbNFqbhVbGZ8TQg6jtISIAYngu/MEkTwOnMgaU
MKJYUIFzoVGXqyCWfQTbdYSFQveuSCNLjvE5Ilix2/OoIopnEOpkc3jwCMoSWSzwxzWGUCBsF63c
rxdSW+D3JYF2DgFG5JKkShd5ypOvZioBlOBRKO5DAM0BMT42kHpUFgHD/MrNEYa+fi4mGcCTJWel
bfdlVybnXv9ovLI4MtssuQLZTv0Ed1HUnzg88LCOOF156qWE4ZiWY/AxBcJ7ZVO5Txyy4b4k8X0i
Aogro8VP+XcCiLRlSLmrndMYYlhXtaEe8lDJzzO8uaruWaNENIpB4h288YSvrrcK4+IJqLN3tcmE
Mr/nciuZCGFR9D7cVrCjT3IgguPDwMNEbYUWey6anmXL7RJgvHeNOJXf5TuTTcpEtw/YrRSurHTf
/XgI5G69tX0qqUVaWEPGcmvSB0jMSGQFJI3GrOG06Lugw4l4LXQUIm7G5ZCfmJOQVdyY4vB3aWbw
ReIconOAQD+2lBeupBBkOqqzyBycGKcLFrod7fXeHowG0dc/POi4SM822gli31Xg5kiqafK2OXHo
NYseO8ImDW9gUEsmnsu0NtHwjZXONVk+fqBuzuz052ok3trixaNlKXV9yDjIu8Jb7+cXcTfgwRwh
rwpCsSF6JjmW4x5hnlqJXoT47eSnx0kreUImrF6C1oKoPVS4mNmuuolIDWXbThKsQMX16X90dWuL
fbr11bQ+30pFwAcsyO7QZSWQAWD/qpylUccOqOL5y8pUDOH/+96RAwkeoIxH4gqCGvV9hTZJI3CX
kPVwZ/em3Yukj+VnGM/6OrEYkpl8gqRDL0J0vY6UyTncqO0bTOsRwhX4WlT9XLBmdisk6SDQTW02
oqWWLOBrRKuIPN64UtzrvrD+MBuF8Uzf0IL1DSfL1sl6hpSlCch4Tkfylfj0nIHF49yREYuyCAkm
Tbo9xAkLnhmkvL5ZR/5fQUwmTktjXqOlgEVC3eE2fNisTJVExEhjvI5RUfLswMuIfJUS+GZmUg7U
Hb1FLSSRpEM5iNdsBAJWUYmyeL5xMzgZGO45E53fuv73kPrJTQRFuaQ1APPf/n8c1cU5GrTHxtXr
asaM2EwV6kcQ8WOqLcZpHP3g6XmeEJDKJtJtNvhk6crig+RWohDnIxjR12owcz8trlYlHw0NVNUW
46E2yvsUkhAuhRU9hYWbuBjEnZgadXVID6JFxVy5NJZ0jVEwU0K+ztyc8MP54ZdoO9MeD4s+DBoT
W4EkLd0bQ0OneUOf8UEWYPsdsv6XhLhcPRAos1fLyOaWIwiGy7l27H5KaClemOxZLHSO1DQAFozM
wXCVWtKi5z6PvnLHkutWhrzR0hxaH/I0TX/e+s5VRV+Fwf+rzcncW6DOqiEZ3bALITRhnrRZnoni
z1tMDMpvTUa1w+opF6nw016dhPFbU6hchqIB5GzeZ0xafROcKSVRw9FNcrKKMM4KUk4aykST58MK
BC8bM1AxgRGiizNu/bkMWQqtkfDziIKwONKTRaSo7ekwo/dJBTBLafOl8XVAIaVaiQ10SpPRbqZ7
TferIuxJzpkkRA85nWEEhgRa5bZuQxp6ol3QMLx7V1aXqHq+wEmmSvN2i3uNW5yKQV0TZCtFAIo0
4weY4woPg4wPl35wzrEmlkQAHZVfj4mI+JgrCBa+7QWgfkfb9vpxIQOzv9W5Bi//AcBXtClkmael
I75tI57ZwTmfZprlv0r/2wjibXq5NPu1M8LSrR4SjEWCasqJaPwf5lCipNUoV4BxnKgM8oKtQKBD
Gg/2lvG6fq7IRJRrDSdhxDIwGZU6DSN3pxjt7K6VxfwT/WQiMLmQuaZoJ/bdLEL2TV2nLpaJjclR
Ld3/PdIcTCLuw+GJ0DQIV72UGgjF4HPNCvMdwrHK5y9hoevuaQSuGmCPo2i3RXpVvR1e+84M+Ev7
iGImSf31TOJlBGPbiTwYkCJyptzFezDIGeFMKZIJhsnlhFdZor8c6SFEkS7iQdguTPxtHC6ocgVu
B1+yJOiSHcvkopHtDJRmktlYkwERj1w29Zkp1wduxVJVfwygNgd8YtaRMkeU70dI5+q68WeCkmHa
IFnyCeld5+PPj5E8UzVgGo7AA1vzLQfvzReyYNktjR5oBqSxeXAH26Kt1OgXBGWCdQ393NMR8zfB
F4WEpLCkruyMiXTwygsK/imxUcJLAycV+driNmbO5dKcxZT1Fs8/bYzjI8yDgJgTIioMnrzSecCV
fp4og/mWbsKXmms6xuAo0TjDd7bjP495CRmJOruUUzUBwxQHr/z+c1RaLyDCMSKNSDoK5SRUqw4l
qRLGsRzGrNzPyfQXIgwflOX260Sd2wEBj/gl6iQShpsv2GdxdzjtbTc67F9N62yttPqfw2BR8JFR
1vhgJ/+i0zKHOs7iG193empC/QBanyB/Qrk84z42xvwLW4Nip/41IgfYLMVC+Tu+05Q9FxZPQ1Qi
6xmHpeZjCe+nqivLAeI8RK0f2NNUUic4XZOVBC/8mwdPhGrJXpt1chubA3jOgzhgQMue/D7VXNRk
upJkdBU//ceoeoi1JY7xdaadYqlDFKFt1/R+x4EXWw6I0DeC3koFDc0g9wQhIS/kFc9l2/0FP97H
3A7o4wwCbPdlqpsnL5nRIxfXXIzOoau8Ug5FkjjfxWTuxMOoLg1C6647O7Cgi+UD/dhwfeKT1BhG
lkN4ZjCnXnquWPaBPOip5GkA5wPRNLeSI4GM4gbEDHHwwMfvoEmcK9GYFAuuisRYlfpBh3jX31rf
KSrJ+48JImcp4W3WhUnCYTBrWUr/hUs/MwRH/ivRHusvNexL9b5uzGhSzop7Yu+3HBgVyiloN9Fw
zYwH0TfVWRhKtSoW3izra6FzpsIAylukPVxhwAC/ij2NphxFQ5uTxb2KIN2+1rR/dmFPeMr5fnQh
21ojDdf3cmxpXNIl2G4MU9B0C9ouy9U8wtmipq1PQqo0hwmN4F5nE6Gf5QF3eFhlF7DBDdoJM/fh
G+pft2JvUnXiQrOFzjO5stgmr0u+qQYLLB7WkmX3W5b3qSXStCf2mmEtKFOx4xfHufjT9GxANFtR
AyPpaHHL+KbJqcj0HpitP0IpA23WrbSFlW+bmT+B1bK0wVsQmg1PlpKmfeI/aW2Qb4ALL9gVHL11
LDWsnsaisVE80hBxzvna3XNPOZ2M5uY3gb/S8CyLXl0/QwSQCMfzLV1yKRHSAGXB2I0dt4KKPjE2
NYoQuhZnTRG7g2sEZCO/rk2ZQ2GSR/BDQQehzWza75/EVWCgwd9CPI+DZ0Loikts5a7FvILXWhmD
6/OOVT/dAChqfRDp1/ougFl4pYGDirBOb4f0Dh8yEN2fXH45YDOEx1sZRTGI88e7jQK3RL5T7SJG
C7NJgccRDwiOnC/feN6uzTjWU+BYDsCL/fwfpssQby1xzRwTLljjKvsAKX91Kk7t2DWAbjCTNpVQ
8cBRvjJ3NrXjMOUv+mABkFGQClNFmcVcbvXnaDFPbDrJpbsPAVcDb2piitrX8fGcWKAWY2kqtC6U
z8GdwZjeMUwGB45Lwj+mDapd+s8/Bm0ER9y6Swp525Gw2fgubCNOEPmJwKwr9HcYD3j5GOKPPNva
dhCzyfPWodTnlV3yG1jcFKf6WwvcT5jrvi8B/AijZpLfRif4u0+HnPsKnydh+7EQSxsHGNB7N7J9
eMldGhgYo8D9JgkoXE8CbeiWEr2QgCnCU0xWLBeJH3q7aBSnN+I14w8eTnL2Ct4ZMPoNI25PrTBN
XJvFTWMD6rNVX1C7ByKvYrQ7bN6lqDxzA6C4JQETMZREX+3UBR3eczXD+5ecDSB5C7fhLsd9v66+
tdqzNyP40iYG6s6BSk6091+0HwCAZFB24emYz6yvx5ppBu1rBVm4+Fqafft339rP9D0DiCAF1S4s
T9WfjLy/97xRbHQbTB4xXYlVVbyw1AGg0iBc5jGNDiF8vvJyv0Akw0S+su79jMa//9UdGWRPVVhC
86Unj7QxhDvP1o/qyGbeUgj/8RClS8Gu4HDQYh2M6hUqqgGSVyJDpwUTiUkaG5CgTjKHt5wmhlil
ZIEX44A0qskmnbTY0DqwhIJSa+f6au2z1vhjE9us57A6b0vkaufx/KBRrwaL1zN6IciLMarqLMN8
BQvQ3wQMedGw0djJhpwE+557ou91EhPn3SyZ6bSYus5s8kkAffFS3LZV9jxiFknJTurQXbRgEisE
6Lacn46/ufThitwpGra0UkcKbMx/dNZAl7tv6ohdn1z2f8RnNBOipzzCa7E99QbvUYCmiqEACKSb
RJslbS0bpBbh4JWHrdHtbIoSDlxXB3K5CdoJz85kHiwAI5Kp5uFeHol1jc1L2qtFdlBTzOX8ne7c
tarRwphUlZgJ5Q1Q2/VWPJJLWhQvLkLDH3MkISIdnWg0SjYrLVRZkCUL4StsPTgWFBKrq3Q1PWLK
0Sqg1Y0039pTuShWNmmk+rkVBK8mxTRNXzYgxqQL65v99cFqjjQp8h7KYI3Gcmcs8kPx55t7qjtJ
cBoK4ZcmYhtLW9gKZ1t8LTzb7K8bh2swULw+FRsLgKgMPf5G7wzgHsFVvUVh8f1CkYqNKvOoqK3w
iNV8SEssHxNVM6Gp9UXfkUPxL29DaTz9dUj2xWkqtGbn94SzI7AE2+ugO33wxbmbPG5Vtq4KDd7a
+m8Ul0HtDuE29sssb+LeMY0qNpWy30Jx92zv5hojrNPqKIWtHmoa15D1pEpEAOhR5Two0P0gbfwn
KnYN9TMEkfx0oEGcTtHmD5X0EMBQUeYnEDh5jDY/XqtJAujKA3J/LKx/+EUByuckdyqUIIIx/Q9j
L90ZsGxGSu7qzPSRL5kcsrzCErvbEcHNDwRKwez68D+IJaGS7zWmt38XY9vJHv/l7a7A3bpuvS1Z
Exm8fu4yYr8Bj6ND9Ub+6hMiwdlWMRXGZCTpL5csoElTmMEBR655i1vfPMOdqBrwvb8w91QMe3z0
g8jX+X4TpRmnt/MP/tiuqosBhso59WRr/2xOQsqpcZ1rYLM8QoO1VDiByHC+Jz6CHHN1v4Ohrdbw
UmfpVv5V4MtUmpRC+2v4q0EVtp9vt5gaXQQCqLsFk4JaOAMUDzfqrKTR4jOi9IdfDIWQeH25yQ4Y
qWpPSXEb5HykZkp2AY3iB+/3pRtf9cnT4vHDf8/qkNz6BBf2Qw14iqtzn/3PEqvPCo5Dg6iJYnwd
Wzh9PpiHqorjteeov8LKpIyk3VMJu/BAUlmWt3kZsfg9P3ZqrhNMCGC6G6JVrHNbVpYPPb/NfkA9
uLabX1KWq+tXON9+4LgbL+5TWj6wqtrfRV4qokCyXLpsT6rRmz7MReafn2JMXxGtR/LbX0mrKR8U
Kr8drI+dI8DHJBMRWMFAZcCqv8iT+k8hB1TRkdB9XZX1/EphW4Jhk2kbhLWGl3OERHqGbIzDwlAP
kd94pm/bX2HSIOiiRA7YS00w4UBz7gurPzv/ymfChrChHKvsVpOzc0IxGviYlLADB0o+UNH07Y9P
fGIeVBMkYl+z5aDvzoqx8dTXj6azyR/48JN2E1Jj0NNB+P9fZs/UL84sVZuY2OazaGpKeLERmgcZ
bVa268+RzGukR450SonOCFM+yb5FEOGlh+tCED6ALVgYmHtLi/3d4sFvxDOsm4i5Wf1kZVNfIHct
eVCBBw/mNknljtrQoNEy1I0klkm51qkj+/HboTmRCjrN6tT+hSoBqA3z6bEUlvPdvlQmob0+MY9Q
7MP1vmcrLYYeMVLKnsZPhUMzKQ5YvKGjnmXenl1/3S18mqcddxQhEujS59Z/wDL2Vu12v2rOdKpk
Ypm88GpLCkdLxy604oHdAKOQhotEmGhpRKc76EYtSF/UCYiGuT6v8kZJcA7FUURKZlcbD16xOqYH
R+71GkgjuFadmdXz9PQPpAXgRziWJiKSQUDl7AYmZZ8XHRNAy0qRrmGQyy62/7wGwB/GN2Cgo5BF
obUH6B5oDbR/jSParBvvk6RP9x3R+iN77gTWyDXQTpkAcxRePbajtyEt2uQHq5VeC1u1mRc5qafW
aVYYUYoq7cT0BhroYTloGXU8T/cymUC+BfAyLFOwYfOuyQ8wvOAE8YhC4RCDW9Yx55fXFIBALDnT
vwO/8x98hkQpU2OjwzvoAb3WLflE2zcL61oTJjumPmLcllEwJDaoMHQieV5LKbpj6tI98n9r4SaG
yQFO+0J8lBqZdRrk0aOHQIiokkOZoK9FnHPiZIlOiUCsyjmdhGpztILYQCz8ADi46IC11LIlF4ka
D5OUwUl4jrWYx/QoHoZxs6dp3DHQW6a/XL48imklcDdNkZSk/go025FnMestuxEiaklur2+gK55E
BPWGhXGjXVOqr/1CnY8NW2xTvngMKXTISEvYXkw2Ffmf7N6gg3qrftyfUD/CYjb/f8tPHFVsYPVY
6wVwBsIMygLQ0+hd28RFeQAG3mkTZAxxLha2xGPYS0hkTh6oazkd18W3c7RgFVzKMzbZx7TioOjW
RzONAZ4DswPd5h6Dw/VF7jjO/CofworndC+VdOTro4YWQUrWezBmm2TVCStL9+hQcqJif+cOBGn7
IsLBiWZlut3uB0/Wz9ZIJhltE+OVHTXO1P5wdLWIcWOmgIpV7kx0YKF6JTh2auCtLHLcZTdWT2ha
xVjW0BnVucsoOtoD6TeeFtibggpEi9wbCxKnFojAxpvYpxPmbyn0XdHWmBJPKBKaam4RDnuJwTm+
DdmT1kS2OEfmkYFPvuECzGM6djaUcFp1rjguWhrZ1hdyI9Kirz4zjE2otySRft5W2QBkxi1yuKXm
FWmEvDv1e20acIHHeXGuXak8y79efLWEIwhAmQcxUgjngoUspHWNwK0qBvat3peBBPZNnS7ZFVjR
McRn7wwA6qVAXFUlLm1jiFEha0svbfp3V6Q9t6vmKSR1x4CtjaTS/0iISHw1QiZw72qEI6ivXAnh
yQsnzx+HklVdRuObtv2IgfqoV1KMT6Ecxbsz+CVEkQqDeY0ZzCj3oEsI/kzTdX+i4xVauEF3TP+s
TANuGjao2AGds1tUlIdJ0gR4wkIbdLFg01isN0C28muGEYGj9dRm6zEI6WleNSXsgMV80b/k+7k+
ivHfiDW1VjoVw75HcCP1T4GKT8UnCDfsShSSosVxQ1a3mUsIlcnTiSWYGeHLYN7K2nt43U8qbWwv
wb2O3YWAc8QvNgtX88TajOcCdE1RvPjy35rqfj/P5hMRHnuFSARQ59D1lBI1B/qDJ8S/9isk3C1o
Td92Ciginifys+4/5dSDmBqCbGA7rmLq9fGwiGBBC5m6dwqxYPvMBElwNoRSFZEtlX/6Alc7Uged
QvB9s4IYHKfwV+cO6ihdNlqOKjTSgh1GQXOhxDyHngXL3Vr6OUcb5W0HqCqtqlvVujOAYUjU3Oz5
s3Z0zEytbGEdrSS8CqbeZseXD8y30LBf5alB+wUb376NbnS2gUPpD60UJsVTo//D73e6FEqSjqr3
YTfKKvK7f0RCI262+imHFYp1M6naLHcoypG2RsCMMyAAGAIcBpXr7MMbGMJfqivLEE9rP9q/AOTL
/VaUcPJOAtz0ID/a9So2odA1KU5oO4TFMyjgbQmwiFG8mks+UDTWHNM9dAKfSdEOfbySrrSxyIid
KVNya2DuGHoHMRHCIP+hmh5fbiREhDQNKC/XDfQnWmP5J8RFhMxALgbSalGeL0dDoyvvhJ7PF7GA
QdaRPnDg9B//46hwFRmEWhYM2gJKH5cjICW9au+q4g6VZrpsnpqPaSIhmeF2aPz7os/4C5c9vpo7
yOsakEqkw77Do36n52S+ee5iCZYgC4amnA3PaFOQMm4AaJR4k+kKQx0Q6r/M+J766CMihou0nUn+
PdyLJTksI0oUoLEHqw3ZBuM40OdVdR++DHIS6MHgCpUDubJ7cYlrHvgdlg2TJE0Ti+Ma6c6ucOUO
u1dKA0CUUvuEjjKNnnaDB1GNr60/q84muJK1hs5Hy4xHpy8bkfqH3woCr4QwpLXy9uxEKcLgd3BY
919UijyDhrPCiQcTmxGvIm6ock+YxX3pfi6i7gXiX8CVES++iKFZa20mzeST8ZLvitSBuupzTWIx
KoJUZUxkprVpRjsGPI983ejHyRm1BDl9F930+/JBsWPBTqDFvprj4k3kG0/hb/FNgN0CyxQTh5Zi
qkh1fjn9rUDBHw5KrzOz31DPxnWXfqQyFDc/doBkKsJ84kXdezr+C1p+JsDR1XbVeVQGjmpw08lz
qKDaAtd52H2ZhQndkP4Kp3CllMI0O2T+e+76OL6+Pxu+zrCi1jqsdGd02m6NzARCJgWL1EHi4bh3
biKcI094lqqGbslv+1PBQhTnfibBqhs8UqcDUEKwidxwQMH1LxV9Cz6b5hu/+vFb5XkpheC3DIGo
edsOkPBGsPr/0b/qODMWIkrPS6AW0azPM3WmHtyY+bsts9tx0WciAuGJTkApDQCAWSXI3cyvtsvs
i7RBgRzcPVstfRDpBofDqweEcQz4HTLXhxRHPmhFc5E4IYglT9tKhZkycfke17SSLeuidC0b8oha
MEpHGw9OK8zxByh7m5qH9h6HlVJwLFfdfFzR60bPl70b00zO8iB88yEd5SiEr306y6Vk2h8ZUcyw
Vy8oZrvTUZzU6OB42J1xM9qxxCeHe6uZsk+Vz/SsfERXbDSOe0m3gLQXwkf6rhJcxeelt8FI9KaG
5trp7YjIDiGYZ3zWaIZim49ZNrheFtLh27KyLERPXi7SeLSDxRiHF1+JqIg1VODpA1eJYMAl4F8n
DBIJR05nuGL54RaG7ke2F+U7qTl7amLwnFDByf/rHd42awFupU/8HF+KzuklwrqsDJwdb/QBVpFp
nJ0xS4p68GO6cA3lfZMVeP3oAApZKCTfDL9lYVtN2LdLF/jp4kimjuZ09I78hMwAyeRtvQFZEJZG
4i9gkbUMob2oEZWvaULUyWn5eARdRlOjhjOCFTHqO+pbU/DFkg/OMc7p83AEI+9K2AyDVfkkox8Y
1fE/sRwGR2SilyTrLRtV3nrzFTuhuhQt7I0RqUXXfyrNNBU7OvKAYT/1uPUNY0yDy3py1grVtaa0
THVQvAZmXL7XQuaQy3+SD26MCbAWxZivQ5tp6pnBwO4hNouGvUlsSjbWSIcscLy8VtTQAT4xQdt9
fLC4+rCoWB2jUnTCDdjm/k/x6V1FcbnOJkcEmaLYitncRvrYJnx3Ofj8HIt/QVuKZ8aIfCQOi2rZ
likN1f/Q5wiS7ZInWs5Uwy9JT21G3dFogy4BK8G9LQ2vagzoKaQiPfRv1Imus1BT+TiIMlVAroYe
OO/df+eG+F3gpgCrTyvcl/qdK2zle2Ku+AOVrr6fsqGjb9Nh6eiCeqD6RIB9Pdu/E0KRw3ZL9Mqo
NufrNcnGjLmLmJTZ4B1HPmGVkFrCgd4i4p2qUDi1X4hn9svJ6ZqYzoUKSq5A104fngwEbZ1MkVrU
BqvkZnWOPeb6ON2ITVeJpHQcjGVNQeI+jyvWjWSl1pKDkTSIHK6sUHgKlx7myCGa0y1vmiVJYqwq
6rgspgn0IhlWPgu1Tjoy/z8zlYF6k2LntQA6lU3u9KcgdRbxMljol3D+Px/1dw4MzfZ8tM0wfRhh
V2Drm6RrvR4wGO+yRSB7IXF2FiNHW5D87VnMubs4E12jzlj33OBDAoAFFvdoSBtKPYRu0tZ7knWq
ZW5Q3I4jnvposZsuQWeZwn48rg2mr6zxhbX2rnrwdZW0FyTosUJ3GapgwkK6aEu/k20cqxVd6l/q
1m8/L4Un/6T1gNy5hkoE+45nFWEKGROAAM/KQBXjYUimIxk03DtfhSZ0gyqm4coLV9La4vitIxoc
3UFVPbNqbT9aQBS1F/xKPMzqAda986JmwN5DLErM4ieN5EdRKJSMaV+qB/paZPPmaXWOvUhqAnG4
YxoOBF67DBB1W25vbXZ8vMjBxoJkQcMZiPxctPuxPIA7UkjO2aBM+t1EjDRDTYgXEM7doplep02x
Kg0LbDgHCe+2FqrIvv0YATzt7zWw8tXZ2MQJ8AiZyOx3aofU4cKCZQhzlZqw5sVATz0jRaj5FhqJ
yiGLLCS7btaJpur6RANdSpeBWOsg4Mk7cB/X3DoXSydLaagE+UBK26Yg25fVoDaXcTum1aUSN2YO
QBZR6TSp3u/qNE+0KloN96Y4wul1EIBCwt8OFgPSUZ/LaAnHgdzdNSvRBAIJ1Ri/rO1Dn85oMeWE
4xUjro4dob/K/XKjsi9IsquypU0wpc+RUXSxRMVQFGKmFzdY5rRA1RUvDCLL0J8iBFocevnNRLtL
dFH+i1ddpDHEHjcqs+3a+zADNpyswUHiwt1MDblHUvp8/mVMpFS8JZlvLGCT6d6QJtJzMMx5Ocfl
tL7QjnDtvNwPA+OgnhpjG8NScE7nxOChLG1vBxMI8o1PkAwXtQwAl7g5WOANGthl5fmosfgCf6ls
ixONNZBYmisarETc8miC7Wf1+mLV3c73tgIklHX6qz3jXnTYpkSdMIS9NLvkAt05qtXWDcwTzoqT
DAGCyjFbQ332SdMNKa+qlaoOKqdMD1iqouWbDvWCV4IKM3Y1U1rMHG7D4MxAyrb4iJ5kJzRzSRe+
GBgUw3UGzL6V8Ayj6ENsIuAGedvfG8xzFy0z0TCfhEb3HvNfELiUZanaFpLsjH/glA9u+cVQsb8n
1UMqkMJlSEqiuYSNI3dz4J2elchTMcobdL8/hHM5ywqX1RVAQrvCUaaRTLVst/7+wctyboyW3S5j
jZpiu7VFEqHtx0+0gSHqP+fhefQrli5R/fkxt1kpPNVtGJZKfDfEHIGFWup4ewvTHEC1mFwxPcr3
wXUzjMIdEqif8601oNTY9zIERzY2bcQgHKnhIFwt7r2ilFc4wMfhNJJ7aNMZaG/lA7Tl2Fu6zpeB
//T71H9TvQcZ5fMlbAkJpp+VfDouO1iOI6WCI9GwmREySTf1KcgMWjBiZisRBJzx3Dj1kFyJQCC2
/uqgoy8D+ak3jYQrt6supQmLYR/p5qiht3zKLEKvuaWjbGfmjl4YhKohJsbe51G3qN7q+SMnmgIu
wbmkD04Ed5xhwAjKIJI7MbQsYu79ifM9vWsiSUS0NWwDVaprA+bFdthlOIuKEzzd/hFiMpTmNO8E
/6LZnFx282tXgaKCYU2kXZO1lY3WUYy+xC5HxRt6sC0fpl4EBt1P7fkZm2W1m6oM/DXk6xGoSok1
9jJSmU8cJUscysjYlEGswJ8KvLNaU3whRG7DRZkGODP1IUdQU59NuFfxOxB/2+ObNYALc+XYeYI2
Ul405FlLb8+yzsojX/4qCB6f8O0fBcUZI+JDeXFgL1FduH6Fd/L4/wUFfjqxMt+r9KjSBEmL8rBl
SE5Fs11V3kqHHAQCjopN64ix5q8Mu7MWj5V+4LiN3whaoitKj1ZMgJ8eEZM+7wNW39JJHOpGV3BW
J5tm5VThfDFnqMW4xL5C5DqIsd16Rf2XmgbQxeCTlGTxdnXTeLK3vUw1QLslYsEE5Yeq409nu3Gp
iBSqaiNVsvjyFZgzlrOhegMKUvO1toBMPy09016Ozv0H5VURBUboj8HlACv33u8t3jlWGopzROug
m+GfcPwbzzcEcoGNIq07fGy7iSTwrW5VFHGcAMmCMG0/jBsOwcemDK+Y7mi79i351cU5tKFUJiXO
lD1VOKdsg9JhBWqi84TetBPPBuqTtwfBFV6lCH3wgWoPdCvbIBOmMjJJM7A1K9TsawyLnka7jMPa
ReP3qEgoHsMabMJ0bJA/2zFI+K8tPauNbX9Wy/C+ucAv2usZWN7cWDPctHbz0ifEG+Oq434xYuKW
3Sw4h/hySnBXPt43ibmcrzOsaKG/W0zF1xa0l8DrSxp9xH2sNYA0sq8G4Z4LdWOsDceKT+1o+4rR
Bqc7+NX6IwLVJU49XNGS1fnx7CAY0ZNjSwoZDVUejJTiNTrkHYfcRYnZNKH3193KGcU9inuBY5uJ
kYUgjI9E+fUSwRNrx1hVd+vG9nVkrZZB0sOWkZ+b8O0o5d9TBESpTMAAgagMsOd6GtfsqIvmAbWT
qRe1D7e7docMW28q0EXy0jJaw3zmjEA5nNuX4EE5frWGU00fsD6SHcs1SIo/+skgj0Rki4BnT+Iq
rqzCtInPsrp5AM/ysHMPJYXOvFd4X4QNfi7I1sQ8A+Y1hytACIG8DhFJXyiBeOqvp0+GMoyJy6fS
7w2hIyrpZkgic0bIHkndKIhwjrWQwwxsE1uRXs74abwSoGRdFPMKN1VV5uGuOZzZyqwAS2YNeYPM
2NWkKRbkJ4twVGfVGVd8A8m16C6nA2SVEdKgD0S6bJ+hrNtTqG68bH2Mg7/1Uh0gdR/c5tkUHmK3
VQKbI4/B2tAwhU+r8HwFvF3sbLpsAj5GvbpJvi7k+b/azcP/C7qzkslkP1sO8tVJNT6YRfh0CpXD
9EOBqSL/9Deh3lIBNP7rl1U/0BAej94Ho4F2S9Z8vNSDV4++Wt6c9+impWGVM0Sv/wOEhmk08gwD
hPj5KVwjC2YD4pd5NW3mLj6+ZwdZS8Wibpbm48q2Tm32oR+STeS9rlFqUnxp4dZQhcxAMfNdtJni
xcu61qA0UFas7M/Iyzfy+xcyuOw7lnE5e/RuLCwIBpLcIE7TeDOAwgstbzXxUkIR3lCd7W0YUcdf
L+4Ok1J8s8fvzMiyMhIES37GCJ1aFDSD0SA0pkHVy7VhQF6AXcfirCmfcFqW2N4xLHsWOvnUYv+W
1UDsnElltekmNcEid0FP7uM8zkpMy400QCCD9AVJc9uwyuDIXa1XINdzNL6KBpwyLVB/fnJgiVk4
yJ0vteTUmm7kjaFSKRd7Z2x1rwXSw/5RZMB69FhvW/evjC4bnf0TosegzYsOcWDkcrmfbsR0zvIo
9DKxMOE1Nbv1rFRhJyJ1FsPWwfA1J4VbUKmevJZWhQPXOvH86Tr0P7qd0NQow4bFVd1OA5tqLxcK
GJgbV4rgqDzwIGGmstcGOSdzBbHsUiJaVsKBkrwmvnLHtZ9XAFIrxCXi5XrI8ixDxPaFQewClBJX
IqYptza+BN+XuOtgBAwbmAgRWLVrE5KlBtfNxLJXqVGyiWRoqGIXP0JR0ILpkuVkqfrdsDOkEjMt
Yu6chPDOQgV+k4/nn2827Gaa6Q42urszwR99a8etBFdR9FMAzZhBFvEzsZW+WpMP1RSHLOMlcWzn
wqE1Z+fx066biwF/cRrwA9n8/JykDvHj26VQhaiquerxSUzEBbl/XToyL7VC0pc0F7MIG5QNuPCu
tEPeejsCIH2kCd5kBRxzYAdPLp774FCRmalWcJgMPU8Jhzgg0r+p9RRX9cNldgBIeySLSjKLZFKr
ddLdQLYtj4LKr6NQ60Y6qo1qn8iMVl23FSvmd91jRWbIYcLZ0t90DjpVxDi6wzhyPBdCzHmoAUNQ
DhqAs3x3f1xNZwFCSDTdgqbj66/OsFggAkWmFL55anq3jR7NS4DBlROCY73MVPPxTDDvG8tnMeys
3154PBF0R8e2lDm9IdMxlS0U1NsUv5dhrdBAdkcdzbh+q38cFikyqaP9KpJdRx++iP4bozqykNqF
YF4DqNCQhJ0CLBfNtz2jqlHluxvQm1eKb//zvssip2uVWKIGca3lbHIN2Disyqqwr1p/+4ndPFsR
UHZQx4Yf/KFH6SyEvbouesmXss/j8F2vd/EBuxRfvcCYEuGG/Goz2YWIBGr4hogAS5xeGpPP0qlp
CrRNOylayz81PJCpaaUep+5zxfO3GK99kSp0gYJrTPtFvHkTx5mvNwnyUHY16iQ6B6c0cHN0Z2q+
BZPeFiEFBzrT8koxxjsxF8tMesuKcmmraqZ87q4+j2H93iNm9OO8yE1s6AAJ8AtS5aiw9EcmP8J5
kZgcgeacgC+U0z/cuX5rp4MPfPrC5k3l0Xg7F4nMEJ0yufEBTLHGcEavuvD2KC456XgB6nVMslw4
5rTvdtszDdDtORQunLV4EJK3YPv/RRC9LloIeYi/gTVv+G3+1188kHXhwhkcbVmzEtjEkp3FZKUF
L3J1EH3SGKuZSs19sqpQTATCNu9bAcqfOpKXBeA/ZvydfgIr/+/sJ6tdrjBbwaVC6To36xO/9Js/
RDpuJO5GGosg9fNo4IxgS51vDUOiC3+ypZv6WYDh/68HbzRczK+IXUMkaa5tbCuT2b7cizVfmF6P
U1ze+w0bYaGybt516uzVwiwiPCh3HxjQPhtIPaU9Y9RI7QKrT7b01ZZKgTeU+cPfdl/l3q0nvhJH
J4eH1g3+N4tvfvSbh9KPSRUa5yvJXoD42IcuKa0ohGfoY/uSdOHGYJHM5rpgHlLik6RDfUPgt+e2
vO41cIMFAbS2Q4w4id+KA1Kta7WCi3b1c1tUTpBNfSFL7Rc80KsTm6MiryQ4ZSsYJ9Sk53i0+I6u
KUAKQtQ1OAF+q1u/iavo+xS6WxBJZlFh6OAcwTjwzHAr09UAhaku8crRgywXci7li04TOCN/FSBs
ELi/UxVPwPc76GgR4NlPCZxbKy55unQc5p5bDdH++j5xgrMJBU6qxdDyUAfb9PZnfPWkv8emk2PT
A2nAASD9vBqJow/pjW2YRm5BNe/qvrMl9NLzMCt8e9SCw2J/m/dW1gexj+FKR40C5t34wp7U8LGA
3MKkXWewSwkdoDClSAWRQjRcXUbjHaku1uSDbl8ey3Nuc2zAvX8Yrw7tbvPP7En5tGf2cESsxj//
u55/ExkpmhaaYeGCSpxQNYRH1h79PcAF4MWLJxljyc5H33FU9m/7LD+akFwHHtB0WCF2OAdULe6O
prFJ+u7ZXUoR0svLMYMoI5rLVcpnc4bSaTGEfbCel80dBJWXj3Uu2paJFm7/7AXnDxUFKB9htoTa
0R9R0YKRfkasi9H6lz6oj0CRhEweXI5uQ2cdYFEC43XIad98QuVdqFH96UkYrIm0cVCDd726anqV
uXyPXAOM+Xn7cK68nL2RhmlONroWOTb77HnoRYOwTpGIpkseT0XJ97Ja2QXDMMsbb1Cfve/ai5ao
YUTTtu9ChLeMTiyA72OL7j909W/UGpHdXBABRdvr5m+Cn1ZjDBV4a1Eu0pJLGT/l/mG4X9UxX+WE
bB92f0DQoeZjtrS2n+u2at6HMlOS2Ews5Pf3/eTr/+N+QWel3Wikt8KzMxaJmdA1wQ1hsw8tZHCl
eTj2T2TlmDFJPt4CSKNipJpegBMyb/02YyBK2Nz+98/PvIUQ2k1NHqaN3rHODX5uUa1vatF4JHEB
lesph7UOk2wcGzhWwqxUR9OVRj84IQxPbTMGtFUg0iF9y1Z6EAZBcnSj4sr1GAipjIs1WgcH17Hr
Bo6SOf/byruh8KWR11WHGIOHxlvrwmndHKg/UbcuhefvegrASlOWKYpQamr86MLV+o7Ix/MoDoyj
8WH9SpFGwifpEs7e/ebwGQHjTjolHEED/K+ywifCRNYdknHJ7Sd6fIEQk3iuGlEYKax9Al8JhYxZ
tog+9WYVv9F91mb0eMxRaKiOfbi2Xs7zcvMlYWVl/VA+38WyxTfD2PfG/PJBlgYCWZaacX3h7Kmm
67wvcAGD1fxykBV/LjqadneUsC4UgmDWU6ThOSHUGHWhdivxyyUYVITowvnC2CVBphvHnyKIhu33
YELPGJXzsgMO8flA7PAh5YwxEKQ4QgA41PWPsdzPmdGCID8KMq0JRe+MfQjM89YCtOEtbNbxe3Th
hcQL1wNHkl9lFYwHOwjt64Ri2yO8CINGD+8HTOdNRRmEu2ij6Frm9rMPBRFwwTt7we7SjyVOc39F
1yb4+gsuaHKA5wgxOLVux2BhIXDcPTz3PD8Jb+hCB10daR+XrAY6u80us4JQ7DqKesEkK2w9BiBN
dwvHfQQU8aBXPuLioRbfzePYlDYDEtZjCZZRYOUbg3Xx5JbZt0PFeeqjka7UrWoHOYleA8jDwoUx
AEuG9B6IsAykWG76v/vU9IEOcsPRDZt8DE11hf1HnEFT0vObO517NBFzFaxI82dIN3lCBFCIdb8Y
pHW0vlNWGsZR/5cE5xBF1ZkzlsZVL+3itbSluBX9teEFOBWdLwYHb5rFRi6pHmOGlzUAmyxYy0f3
HvkqBTewL79lcuTuGThltTIrJyTOs/LQ6cBQJj3+fi3FQy0TNbvQ+ZolQgA5DsblGqq77SowvTFt
K8c1+GUrqF9QuTOGsdCjShDi/0s91N9mKN0qJtt+nmdMGT4DbgqNjNTkbVyXvsMD0mz0Ih7WoYr5
hX7n6T54C5kB0eX8KWMFDl24Vrc8D/cF/V+zTLs85OiQRpiK/E4oST8T40kAel8BDBnD3jLoS8/A
pWFrSCmmR4kRmkm1oxfs3esLnQLY2OzFaWVZ9UNv0wyzMJCUbz34en+ncTh4ulCTVdykn4CD0dmS
9pMmjg3N4YMpOqtHt8Hj4/ZuoEbmZs6Zmd4Y4Tee3QTzjoiAoiM48Mfb3KTC7EEjXeC5U1z4Spyh
+C90Wz+IAlhAXo40TNwR7TCsB5wH5cgdThwdczOo2BJoINcSgwMAIS1+qne7HQba+ctPpwrN41ro
MH1yXvhpyF7k2R3JnqrkgtWKOlK2K6VwNcIcC82zaBDcgW0S5+LH8CXeFMgKVlIW5E0yszQmuhSL
XRcF1ogwry+spEM7PxrcGen/7Wu6RWcrmUXzfi99aWL00yB9byHNQ6GTO9yeqk6t/QTplE9DNTVR
/OMRwgS+Y8J5l+OruCJrriG4POeVixxZDbsGH6+jolzTyxiDdjCBw6dkeIrN8bhOl8fnBCzEp3wI
7MTSWscCx/CUxdGU3WqAXpAOEeUBtQiKvn54f6pF8jPyRbrct0iFjFh4TYCKMWAoByaigj5aEC0N
HEag3qOHFpbza3zgAGISuUQ5Q2DuJ95s+ROEgd+w1LB+vP65/hLuUvTOnXjXOsIajTHUAKb8LDwP
tc+l5OMbEh9UVBhg4m8mu6NvmgScyQ1NMzdQ3ZvnoK2d9JuWJD0CUbS/bOx3EOL1mtalmOfzgQ3h
kmDGOhiliw49IoeIZ9ERrNmlsCBllbLD1kv+r9Q+h/yiSg5RsICXF8Z/lgOyD1mmRlIqV0iUQB22
HGuA6jVxPiZXh6hSzMwMoljyaYie2aDrWDwm9NbvZe8579w3+G4h2P9zMC0z/RzLV2fdAIjNq33V
1Up39+zcjDDtM4BCbLNCPMZfpVBSK8L2ylVmpwOTt0Ud3eSd/R8onUx/TgRRp8uEH/At9zX36Ox1
1IWm8LawJJU2fqYvRbOK8dde+ksqtj4uqoLP/4O30YrdV5bM352y19+PqUW3X/uVJCqU7TUQYeMD
fuqStll9zAVdIHXrQ5Oo30ryvnH8stC6Tl9ckYBsqKEJ7lAk80zE2ht4b4S6WRCHXAbPKm2UCd3x
i+Y9o3QTtIYWD8pCbPfbsBMqKtqU+bTc2XVHntfNLUPdKnLVqEfk9eBpDHGVsvoEF+w8+Cg0aUq/
kbHUOrlx+cYx9WtmJv1kGUtwVdhrc/bmVmY3iZAVCW1q83aWTQFXIW0sgsk6ibdz16DGOY1kOl9z
SNrXoSemay+VYY6GLwP5BuEm/Uf3DjtLq4LINv4mUCCDYV1ARqacFqZsE7pj5dyY3N0YnkYbbbiy
AfwD2Hl++fkm1j+BYO9AmV+D3Iwkw/zibxMMpJetoVUkh7xbwI+R+xsYVzdLpt2kj0dhfyEz2AwH
XezB2irBZ9SJJofxGSyLXSf1NgSCSZwr/kyKqzWGfvUFNykhbUuevhPFG8gBwKANTL8JfHM3rsW1
HgTZmlXLjvl8LpXXwcEYbQt13HQCIZy0q9FtMMt8YrbZJn08KdrAQ7pqcPIgd9bX4bbMga1Hq6W0
Q8sufWCl2IV3SKeaTjT3DbPKf6eQcXl/bUk8v1CrqWsi5ybkU3Q1AOrhorXPyhK5zu5eBO5+rG/Q
8N6rsHGsVx26BoZztPHXF0oTio0PE/uUMSYKE8pUrL7BEkbWFl096JbdW07s2FxOiWqYIXYvIaUg
IjuzZ8ZERXqJeqBwtnMLhNBEikKUrAbGKvLU1lkG9ODDujsWQxGT6X/4J0T0fV1ygBU+7UkOzJ2X
E3PMoBzu4pj+aADnejn5IGtvNIIaoqiiSMINy0EJ7uMG8xam7BsLlcJe+WfxQy7sru3RHVIE7Dxn
33dzhbv5yYlfzdAQTzZYBHGRbH0lNYQP54SCEU4yEBSLeMSmQ5MtVEP8+muswSCwoz8yzntJtTij
GYbOszwp3CAWpyS9UJ1qWaKHfEfZF6xhi8C59ifv0C3BV5uh33S3TNMRIfGuCNWhiC6TOCgseACi
/MpHMULkJJIkgRi3Hqsqjs1iW3MiPAmSMQ27Gctp8GONqggioopR0tKKBBLpDBsR6YXGa4KttTp2
/h4fRkXV/q80m4HflDlJ8CwykFnOQYyBoHfAirSWj2Kg/n1zHiU/NVXe3OCbpub8+L84pr5KMgM7
gw4ZcI4sQh5xybT5gWpOt497Yphir0nA7LRVp4M3HP+SWcEQnYgQCkrkK62DwcVkU+O64y2M1/lM
Rf9iZc6U0cdV1RNua4XYpu9shzC8sApA64qVIUhMzvtaqDOHCL00AIZ8dwzwsoo794Sbl8HHEUax
5VnjAbulO0at0oWVHX8xzrARqeKKBo4t5FlmKk1jO510Z16a976u/Sal4c+FZdOoxOtcAT34ApRJ
ymcQJsL0aUkwSQ7vh0ZHwilLfMRCkYRNKhRbnyXrNu6v0UaFlWGCXVy4BZ4T+mJs+4SbFOaJU5AZ
KANcVEeWy6h1SMFyX5yvulatrcqXjyZq+7T6XBLbzcLcWiVxq05EZGllHSzUI1BmVFjxHC5OS0VG
Uw2TKYVUvkGNcD+89rNUBKbOfmWozwaiQ3cTRFyNvjgUZW+5F/vS3RB5ctu2/mka7+zyej8mWxXc
+rHu3nca9CfXChparGEZOiocYqosCsLIgjQX2dmtZrFgNqTOxkXGZSpGRfKK/4WD1rUHWLDVr1Aj
JLibBCxXs4AKxW/K4/MK99q+WI/MHu91vuc6d2qACwygXcsJpLTrXnGIcnHV7RYX8rBrM8b+IWZe
VUbkwzs10FD+qeVh+6uo5srutOaDA/XAWhK6lW5WQphN36Lw+jeo6WDxm9TJJvO1JosvX89SSLGL
AYAtKZc5AyARzMyij1X2m/4HXtnr/Sn9z2A9ZmWhaVZhLVX8BlG1a1b6F2QtzoIoN1U8BjT8NDQW
qmLQQ0idhKuVjZRPe3ZNo7r5pmzLanTDdKZWmNuIYa7gYm6R1FKOZj0/DnV+tNQhy+owZyD2bEcT
DJKEjtM9uV58mjn1fBBZu4btMfNOuz+wXXzsGMA7i7ipIS6CReP38B9hA3ID0wn4L+pKsa+9pu9j
grYVqLCQzdymd8Xtllby3qhDohA6Gc+DMo9LxaCt2D2z8uz3r23VjxBiZD+ZDg2wg7t0bWNGBDMT
nVo8OPgtAVnN7nF7T4EykXgVcPPl/8hkM4kF+cCq2pmN0BAMxJpIQ/y4asHfexXSlR3ia4veGWhv
J3meBBausfNIPCiyW76JjyaCcWsol96/vgndH+ggREt9gWPduB8Q9In4jFUUGA/v4F3h7waH626B
txtTRP/vx37AiNWM+jdiUKkucPfpna25SBl0e9joj7AnzkZd109L0kqz2CbcBtyxjiY4WyoREloy
uupOw5ToIORPzifQVp+a4sSKD2THCJu5j3QyOfE43H2jzSDWR0y0rwIhSjyWLn8azSquvucYbKuN
tlErispmEk7AYxnQD3/+h0aNe3J5Q3ufwwo2l7EImUQgsiFMT0KHfmyZg/Qs/3+7vyYv5c627nfN
oXipv0e2cynaJfueL9usvXLqVeLaGuEnH8mUE+6MSTCkPtCUAlVZoPBdt+nwfF8o9t0Ygo8IKvJj
XTmZCMz4FozeeYRdPpHZ6vKYSsuYzqSh0oMq6XRWgAnWtZpjTXDUlej2kffFgFzWtSSHm6oejqOg
xuyPIHrfIqTlnHEs1Yy00Hnwue+n2xg29OpoaUpyp0F6DtDpcLYeoRHr1laXy4AiyOlAoYelu5Ow
vhfmk3tmlMRoYxaUdHSNgiQ4o18EOLO0l9deYFOZKEEFHiE1XCp/MhviDEhK27qiW1jyOVh01SZ9
CxtZaYyFWcBJzj3kfTJcLd4gkCKxgpagrEIXRC7vCH3oShxXd56H/xKwBibpIs1S8/UVDPiw3lMo
QCgNxZWxYljpzWvdTWZrCeoHPzW9dUYNKlR0I9vhxPg6TMcJvDWPlpNUXf87JZdR8XzH12mIeIoC
zB/eLYF4DJ5H3Z2LwY8GqGWwA4Ma3PP4EjlBCX8BLVj1U1kSfzV33sLpiDOueLF2vfpPGFUsa/PP
JtbI6alq6OZ0XiZEhtTzWgIJDsvUPb0GWPE8qrAcugUrAts/nJS+u529vnpXs71kaftjiijcVxz1
ii2JBrBkYU8gBImI1pXb8yndzm/SCqGAqPUegyQ4hyLDr84nx139i18rToir3nHXXzuOuMbd/ZIV
vbf2mZyxAdEJg95Me7dm0UoFP1sFvNoSuY9rzuUvemKmZ0tNlJ8T62NAEE4J1AEJmPqymSVr9BHB
J9D53QTKWa1Lx4dnA3Cw/4cplXOxwdaGTvMu/4FXUIMIF4a7qbx2h51Fk5I0jMAGVrZ1m4sTo0Pq
7zPyaHGTMEw4RZ4ui819eOvXp2aEg4FfVLtrL5o93TWMUAEwa386WJXTFV8IcLcjcUyxXgw/sYut
nhHqkQs2fSAhIGeNnBwQA8JmfEN4TdYGPAC+PiW3edVmAvOyc/WC9d+zP56FgSXtaAD9+Sr4Tcfs
yyyPIvqqQwB2WRjji64Mv1BATYkmPevVUAkx/a6kUEYMHfgY/5OIG7CxUYHNcpdiPavDv0sxvfLb
8TkxGPQLLgOQTG/fQjIYsq2aE6ezsQdJVSpHdXj9Wjkfv6Po/vXT/xrwLDCQEZrqcSnQME/348KI
kO3n0JZg1m0DLHDF9k3bfAvuBMIHH7YuoQgt45IB0muO3loqhnaQgyGlQDNcaCVi5pp1nfOqXrSj
U3F+z7fMsQbcs536rPCrZyFVyrF1Uh2O8s5ERP4Zi896TuId7V3vFIdgPpkvjE36odwu0N9e54oe
RX9eEBf6GcWV/mb/1KcmhcA4Ydige9SeFg09s7xHLWcm+MZWcRCHABp9ReVBfo7pzYHpa5+SXR/9
hIzqq0JdvX9Tv7RL3S0QnIj6rhTehA2n5LNBu3gletGY4b0Ze1lJrXCBZcEgRuLNo8+O322QUf1t
1jdv65uZuXgxMWHwtbJfZ2OaNS//gYqePUmLHO+q42PM+Eu+sv/og9quL8wSlAL59OK3sGOSHuo5
XDz3I5/C9ywjbFm1/00/ORODC4lwAwHvF+/Hh2Qeqdcc4Kfo89SxpFtiIh/znHlknbxkTb1/vTAb
qhrY2JLu8K/f6nhSNvguV7t7eaYsoeNAHuQrNSj4f9uzHj3qhwSsDvQu0Q6UjbvPUC6C4FHDqc1p
s7QR/WHUbCnq4FknziXglzx1GJ6+3S/zZAM6EHyoIldugqzy9bByy6YDRIPJKAgj/rz/Ybx8TRo5
qZyT6Gcc0vEVJlVg70nedgF1QNSuBFymikab063x9mopM0cpdtiGKCtsbP3Nq/Jt30psGEUuzjNn
m53/04veNkDBgIR7isiuht9yMfapwfaz0QiRcJrSQQyoUm4byTWgk6aOe/bc2WP6AnRLzU2YLeWL
6qTumB6BjZJB5TasRtJwJNzWmuEtkxhRFcQkd6ZcbJMBx9E1tb3taOjh5Rc8nBz3VUnMw0ASTuf4
ysOY2RItlCkPnsn3I8n0521iG1++JnVCM/5ClPJHt7FZUZT7q1kxMjZ0icBo2PrfCzB45RyblDiU
TVioyON6nNp/wOOsCJ7W7nrob+HDUNWfdPAGqYrinQaCtebAw19+XZ0th11LXTolw8pIkoLb9S5F
td5cuYaM9dqDD6pcX+bmp5s6PFAy/uRL45GoW8WOz4vTZN+PUn9ZvqXnNt55t+59KmZTGBsBvCdI
DMwZbNfPu7+yaX/FJHRa17rCs+7/kjcE2eUK8Ie/ICxsxEO9FCQNotoUF/dDBvulPBhrO6UgFMW5
e10bzSlZWw8Z0UQ40ZOgws0SH3FP7v94wBVigoLPIgntTntJUSPGzV84bYgy1LJ0Jb/hbH1pTsUH
4Rj5NIsAiFMtgfEQO0DSu/YJjbbPXb5xcshFHlioS/TDx6OBrTiUUaM/LB6fzE+TGWgF73/8Rnp3
KMzPw9Hl6OSkW+nrnNOujkyNxOfbAz0/w+U3oTIdHYiDCIG5tQCyKeRJQmtCBSx8xYZUQhzw9mBc
lmAT5CuSaVTdNX0DxPhaj+a1Cxol/DmVsu8S955ZkSpZs+Ie9po07f3br/lwAyy/fsI7jz0ERy8S
RcC0u/tfxrcop8CTD077eBM/CfL6ybwTrx8I5ElTmNneQ+bMujPfEFFkzxSi5b+6N5J4aioAwexX
HvNbScYUIT/3tWb3FpIEQ9UPOHL+LT8oRgtunwzWosph86SyP/fmPc6Jdwf4yOHpomXFk/Cm7bbK
UBwtBUo9PeMwt4U4JUVx4FSwE49d+7RDmo27VyCEN+jD7GOYErqTWmF0CX1on5mr170oCrTHtMMG
Fgz2RGj3KvgV800QF4Rr2gWSUt/txJBJPVVciGHOZLn9GxWgVY7vEomyBtZL2C+Qkr01nkp4eOQd
PDwCy+jsWPtiPfAWIYu7q0wQHVvKqhRjZAYTMeFlQm0DFKcKrtlane9+DhzW5P0hcKCywJPq3kEn
CpvnFhIWiLcuAbzn+xsbonPm1PlXXN7CAOn4Yj9lnvddr4mEdfv5TWMDJ9SSC4SXb/q6uw/liv9h
sEO+u8/z13OodWbRutxgBfDhpjD2P+6aTToT1uGcLxx3WaqBEgBVX5HEEy3KC5hw3HEQfUr8hA3m
z2F4yY/agoElGLyuRyUhThujjsu/pxWWeMPUNlGkOoB7WLpgmoU3vqQNWusKNFTnjxLzndDopEq0
cxSefHBFSM9MS7T0cfLztaVPV8zYfYbNugpwVmb5lVC26is47bMG2pkxgl1fc2mdmBiOKE9QwjRO
6x6E7DZ6P/e4x02ixTAKFNGHP6tD1rXZpYCod8B8qHRkrkLnbB+RxGPk4GwdItXfEE0nGh5xS+Az
XpZRUQllNqJhcNky+0K4XEMxNm01Te96PRMTPL523VBdzx9Rm4tQ5KBINz0MLeIRf/QZ9TeC2Yqb
HDlNM1mxn7WnF6wtdTejB7QdHsgyVi+6qax/FiFqJeQvUf7UJldn701jQc7bljxY0M1PeSGd3HpD
PnHmkXcKvxw8TOANRinCNZrg3G7usL9tyOfZd3JacKVlC8iF0qLHpdg1kKC+fd76irvO5CJxc77K
tJ3h9dnFOB0P9fuaRSiR5ZBPTPhiJuCYXTwmWA9ytSQY89wSrN+WBs9htJEzNUdWkP2jYih13xEU
R2uCgEEYxVa7lh7NcnQ/5j2BYkbXxoQMV2kmm8JdYIeLB1AkuUU4ufymgxqAF2MdnFylr7C4fS7Q
7O12co5cDIsrMPbZF2EubUghSBl7Ld5D9EM8zJSRCjFS9jk/BH8GxjvmP1+dM4MzWifReo8i899A
XrXe+ZjZ/07DoCxSMmxw7Wu0RCMfm1PewujCFNEkyS351kUaLnV0pE+W+b5MqdQeiAVDqOJtGkK4
GbkE4+dW0+yPXIrzNlKed6bLDZEWZbp/XFg2EL+snL+8z1FJ4wwmGT8WUGF30Z21ryUqAOJpBvHh
UerZaxl7xZelJhX+TvZAQubjM1qrXhtIuQ20e0htKI7kfrbDTMo4uguhweJZf953LPguqoWZ+q/S
7uHnhXppbHprZed7vwl88p8aaKr1fDaKBnRrWLUq3DkPneytIaRrzOD0zV2jqOzpTArRyOap2Gt3
+Bg7sdx9epgC8gbmzOzWCZHa4ZUpuNgPPaXdn7VvlS4N7g/vpCRrS4ixjJgWMe0aema9shYWdna7
rwlzQ90YLFPWqpoAr31YCltpCwefw0qEfTMLiRXWc0tqS3SjdWePZna4ZVv+st5al/5da5tXUScx
PcQ1zqDazvEN0pYYZdsLbIemHRa08CAHPwEZlsIih2Yl/PunyHUg2CGgNI17nrEJWC6nLamuiKPh
LaJ+jVDr1qPyLWxTs8MAqxT59JIKYILqDOzaBYO/YaMf5pc6N3/ZSBPH7uWz8ueJl0rl+UUhxZ0S
b1R1GAMQh2fbxotK7jDRJHkF+ebxMkt2+HnjfGI97lbLBA47pPQtMOdnNYke9TiIno4xOQrJJ+gw
2so4Exkh6C8G63pFSlEb3Mnhwwfo50hVZ3k90Bzc8qNA4Rgi0g81rZLZHqMAsIBEIRXOACkETKrN
ctjE1qaoRvnB4QrJ0gMHbArDS6D3irPKBsF4LWGwdi/8UrxxE7dNoQOxwrQ1lvZ96QPEzZKGG1ap
fwtztAOzUmKfddMgg+/zngnBdkQMeA+UjK7V0QtBiL3fPmndaQcVJ/DWOjErohuy2oNDL6EO7Jc9
2JlECwuu+Knhc14xlh+b58k3yiqkDYm59oPQ9K+ufCcTTDo9Swba25PG0HLo9A8Jzj2bGNXJnbyy
2G26knzsuDBTDt4YDgTj1JNMm4Fs5wJr88pAgSw8xHi/0D2UaERjMshKtq8cTjVdWkrpedn5eDHZ
utBOljOKRItRDvNJkeVv5ymEqCivaE4FQ4/cN4Q6XAt+LOv6e28A1/wAA7KXzn5IFjHPJ/u+YQ/q
RCAxU9ovIKyKCHYbquD2JduTKEVIPoYMUpHXUqo1kJU+T1b89sgF7eFTtpeI+1cLYZ6E9pV/1Bmx
Y58Ng1xJu8LAn31wfl7sMVJkrLbnsj33kGB0eMwkdrSosH9LdxImSLbDEUoMxGBw7SJYXJyirg3x
gloAfI34Cy38g2S/5/RcbT1AwKrn7MeXleu8qE/pETuDmCgj/1cpnP3FpD+Ya/VvGpmdcwpua5hf
auJAPQfutgiVvhFNNnpJy7BG7x/aNMh9u8XSZbXipU54TpgLDyiiqHwFxLmiM7Yzl4CUQT7diukV
s5nYuNhJuNN4PTUdceUHwZydkqUDy8d+8L/0Vkn7YmokEXSPEGqQqPIRBtORxkH8+k+4xOe8MNxf
wvIOrTEsIAmYZ86CWp0GtxHkx906utAp6c1rYmnAzer0nwS/jOJhxSpJa2vMpQE70i0TNMRnoUuU
jBMOtWSSaHLR4O14lLMCEA8NapS2zKnOLSaod9pNvYhNp9zVlLkhpIkNUrYgRgr7Qrzrintn8rUz
DMfS1fKeXjzx8WwTlSCHeEEBBrOv+9EfKaDk2sz6YRy7qONZyqdW6lrsIb4TwwHqC0Rxn9F5k0uM
iCdfXPVfacKBYIqAY8yYoiCUorNTSKJJi5VzpbsXQh6k4+dBgcLywXmYeJ8/uQHzyKuhOB9d8DmC
FjZNQhEUhXL68Ywa8rItF6SLGW3gxQrkv37Pi0OWIAocXBzupBMR3QTapbrwG6zEP8GDnBmE1NqS
s2XEU8KgUWvh4KrrEP/4u9UhEnWXVMJ+YcOY2uAmXWwxGdoZK1pdZUWdl31M9+ljSZfMjJ6PCeGb
XUu93GsbSH2BwsqA5Qc6PSJmq0zGi4Ne+z2mzA2Jr2bnsrvXRCLA01XL7Y2rMjWUl3oE7uuenEXQ
50ybmHo3ER1YHXGbyO1RZ72+K85msmgoY+enQ6GDa/m60B2y/ulTCRqwZHCW8Ff/eI2vknNj7NpG
RLoDF3oaZm8l3LlyZxoUwlQRdlnrMoNCyiMJ/H+ZgJB5zFDylf9s4ln/IuirV0+2vxFdHjCa6UOX
E4rgzJB4pgFq+4qfZ15gskjFspsLnGfb4XVF47FEKISNJuvUUS9wCWvyLkAENuazQewnYGpNvfC2
mwitF5OhGWNr2KC9rFitr/Msi2WfZD31OTXySiizkP/550Y+zqLwW1MiYviGrm8CgCb20tAspNtv
yEEG6aQj7uDjGHaUHO7NwuTr5o85/bzjQxRGFz1ZQP1NmsHoeGWdqXG2tdNnWwQK0hh6DBU6Yi4R
d3pXXlcUYBkaRHZj0HgVRqnBgt8pjpkktSQmgfwdMeUYRZdooEVoRV+k4ofArjD4lVGygq+6xNyh
rs/XbkCLj2rkbgsWqzd6sWnCsR58zZrMAxsQ+WAajQQ9+8zZMiqQKKIgss6lDwEqj/fULB0UAvYo
nhu6EDpqgPlDFBmk1681/ulktKUMdruKo5VYM1XEPdiNg1JBZgirNHM1DEP8S7Zh/3DI6VJWDJxs
lhJVtsg0fb+LVu8f6vQvvO/5KwSCyAJryehO2J2AaaJLhXVrWwWoktyCeP6jvWcDwHOYXVhqClvu
ue8B/3pK7JI+9r9TFiHvJZeZnxDkUIo54iYg3tFE0Sm9Op6/b85Kakxg4No6sJWVBWy5qWJSu7Vp
KP9XzQ7AxykoRbF5cmrx7tpui9hNfwbRe42n2EhePLjO28skuXQVGWdJeq9NjZ0LW1p64QqvXFfP
TvEFkr3FMfDDUsY4rVWDl8FlgchN/7qLVU9iYF5tN8qnZoXjoNWK45OTXKsjVqKqw6NbMVFrGwYb
yIsj+ALEccOaugiv8ftEjarg83sZD10KYzJOmkqqYF3F3S2i1CNVlG0gJPixw+d+BQH1BUAzUy4b
JsfEsiPgusJSDgBHitb9oj+Gt+gOcNNhZr3zX0VmT4hB0Mx1OdhuDNT0vMiDoUgOcRt2IyjaZ38O
tdgSf4o9NKwC5n05kGAuddFyRoK+GLX4s248rPgvNhbn1Tzw9ALEwKhkthD2E0LvjsKBeGTAGkHf
6TBtQGb3axbcUx7uSa7DYghzK+hVfM4Hd0BoGdalMJQhLUdkQHWKCMA4/xeV0sjZEFqdTxMtxHbL
Op57miVG/8/350M3vDhV1ZvvWhtBWNzPu9DmbkNT/uxgsIMnWKdyd5w2QSgSmMnwv6T0OVUB2UZ3
+vmQfvfqK+EFfTNMCHmxFuPHbjF2u0dRxnSOBVVg1eHl5++uDwJjMVDmGTD9jEO5e0un+tyzJzMa
IZv4nJjTfXvx95UBXffWykQdLKZdtaL3rBL6PLshPqCdBUlm69CdQaql89wzEp2voY3oM3EmmUeN
+S7C7hKizyT77nWEG9NO64bI5pgOTD77IMwO6PlnQIXlQMcDHWBzVjfa6pwNy8O3fOiq7EuD0WLJ
LdpVhZnahUuCT3ndfHAy4bbTCcT2EcoQAjoh+YREO2Tm258cp9ABa0ekAlV9oNpoOWB+ePTqC2/x
SB7i/eX++orQB7NKU/T24RWO5ykIVeuUUprUho/dRKF9JVBkGaZphucoa1smEentB3IcjTLD0u7s
VEfjjR1Tvw1xz+Fz3BXYwnoz0nqQqDavvrVYsCXtBBBuOfcTjeay+4MVqDGxi0iufAVPAq8tbpa9
tZQkCxasMIBOGikqV90LYjb4skDTS3L6dIiQiCw3CmTC6aTDTAfzbhSq0PYRjDuqXp1vl2AZ94OE
aOZyATWRpBq0ot/D6IXLN1AxMGU7WaQS9SE7O9S3BPJcWUzMR+PAOF+R8CBdtZj6wmv7iO3dgBhs
Kyxs5XTnPRdfGdAkpY0nYb0Cix7Z5FmGBHy/3foEmxqQw+cU34Ne0I7e4ZDpcnvwUannMiBXKc3R
DKpaUyo40nPJ6X4abVVYQ22rjpzFh3upbCNj5GbQUqqMvwEK7Mqpn0skpvPwJpY/TDxbExPhgWOQ
PDYu7NQnBbaajmG2CfhULWBAwXXUr3d5Ab5atsBioY+jJSmudItfjw3a9+RRbc/Bd1Rr1P1WHJRQ
Ih65NMsiwpOZ0FhkUNJbW418vR9Oi+WTIBaXA3Wg7CUi7v/WEe+aFZHSNG3az7D0onnZdyG8woNv
+nCWLDDv6hhwOf81MjlV99z/bPgT9UeN39/vnIJXcgRNGb08vcGGGXjlGr2QncDPCdJ4tvCvLXNG
/XWByjuw8XY+xfpXT/Ft5dS6VlYEDDwDur7s1mVwdaVd2MrbHdoRQ4AkucQmF8SS3zOtQHoGo+Wc
qa5kAzJIEm4bawEvwisRKOapvIz2PCzJCvWRSjqFcVcNXkDFgekNPocnp5x1d/Daa5nNLVJzQZJl
Ms8/XLopMNgkY+DjYRzGH5795vttB+7dTj5iP9Z1vGRRFQGsCg52u1Q1sAEu99E57k49YlCPaKfN
e1rBDcg+8hr3BtznZNp3zkB2y7hPhsG5yhQFE8DQC5FIJuzC3m3IzIU7XGKZDML+y2+B7T4IVJbF
GYDALD47fSfHhksTk+ud89VhGMjaWwRngBHAh/y9PTqgHI+9TyMk5s+yVaxo3xLJN0uswe0gyFBr
G2IcW6GYQE+Qw81RSv6mXrj+Ttw/ZyaLszZebgeXVo0E6rVNQrvleNTG7sIQH5yKr2OfUNT3z41p
000DJOCKPid6TKJDi4fYqTSsBB3sssX1PDU+D5eU9qVIM3Fq8S4+riuksI1GhW+/aMq776xWjPPd
3oVqU/KVzsxJ4MV9Nc7fg6f1l8pOKR2iTHwHgIR153wdTM14nMKbnfMooGkFVObLjkr6YTWQGwSu
defrov1t1tiU4n8U66R1FGNjdnM6G12+zPJQQoqapES6gBVGm1US13BSu3Pg99ew5jH0GAttLgh9
WoT2d6K945CBW75QmLbA17FdWOLQDEmpUHUZYVf7p5TWUrSRk2YADQiOiCWeLNNSrIysQvbAZ1rO
H4mYmNM3r/8+Lcrrk3Dgtf8y87xtNcACXg2xRemRQkoelpl7ZO+Y0SLJ5O7VS3O0Qlx3sRkT0Ezb
zWxrTVsrOXFRXfWXi+nYuCr8iL/mSmNX/bN8GQFYvSMEzAvjLWC3r5c6OSXJn3KXgx/ugcKZLjyh
k8v+nIKThbWw/EY4T0T2tUVXI8MxRBnvbOE/3tqM0fE76LOphHAPUi5g9/jA2Ny/vPw0SicSVycm
PMgcbtXNzNXYl3YGcRUq/0rrvZP3jeRLuXD1GygirAMwrSWIt7f4x0XEY7kN2pxDDCkRfiWkB0Z/
hOjSUDmYGkypL/q8bTZS4pj3QkQh7fpSL7bcnXcPT6FAQNmOACl25aXTn3JSnTOBZTie4Y7ayrHu
ZXeP00c0JcCNcjaV4/GIq1qPUcBOUFdyKOisI8LBvPfH+PjtwdtYfqiBjCe7D6R0wk5bqv+7PmHm
BXeG3vzNZrs2QMigp+0R7qIdct64wLnOX0U2sQJmgIjr5fctjIsk8TGHQpgBK6MjMeOoSgHIDYUK
jMhQA3gBa/ZYiUGHjbPGwDKb6sIWFLg6zjn2n8wtVcI4cqJaBQ1jTXkam0W5bLgHcw/ZKyTejSqZ
ypMznh2vYP/5tczZM5NwPIgAsQe10BQpoVpW5EiQGEis1Iz2w5yruDwJ3K5DWh8MAPgMM1uTa9qu
QYhwIEqnY7VQLKgdS/cRgd3lz88WghThcipeVcB0MoT6Qq2OJgtvGas5Y4lGc43qpAN36uNFHABx
nNYHgo3H61GFcQC+BH3ySFtPWAkjzg/2dJsoizFm0EhcJIs49bNaeiooJ7Yo/Nw4T2SDtx8Bek5L
SXjf6lZioQpO4zK+PZB4Tk2zYyu2OJOk8jMIDEMBImuWplt4R5NMQ2yIAEd0hVEzcVAJmnj2xqs6
UNvqYMIZChYQA8TrfLPagiLJyyD34Ad5DSYsWuI+BitJuUPGoRxeLmLuM8QZGiyT7VOUerXkiadB
hqwGAteaEmPTfAnvRPcttkncyzDCUG3ylXqQSSSmgrDV1dFR/wPPYFWkB4gXFO7Yh1MZPyvOeC5C
T2eXMNmnLmr+WAyAMqUIqbNLw7WEoyYDmuURVQeHcVTi6MoK/SYHZZdqwW+8LhsDccncPCGFIhbT
eV1JSjrXnyWzCFLZ8QdVT3HH8K9r1atzrIlbOU1RMN7B/+EyW9qrM8gup+KRi9pTxm+wgbt+EMLd
/shoRZLXKtraea2NERul028BQ5adZCzem5XEDJoHPC5qVcuqSeQysX0Typb8Kk4/YXkRz+i3owBx
xTQlN1ffLfEcSSGpWOKV7gbtjPYS0Ua+q9vk/vNkMZQhUWPbii4IeCqzScFskxOVEV2hFcl56l46
BtjZotFsCzcHpa5cJmIPBCNX5XKO3BaEWmms0nWz65Cl4ip/6hNaoKfd+T3ExLr1LSrUxhK8TvQi
7IRmWEmRqL2X7+O8Dj2rfg3z+SxpyeLc/qrlf1owbZPnG21EnGlJeM9rfUxzpiVQfbphFu32PCfS
J68aTTYihjooEVC/URY6nS7fGlH4VBiQfYBTosFl+WNiBX++B+3i/gMvhMVvVp//C/CEHvisO77X
/sssWy/kDhSIzMS+Bn9A6FQQ09e+Io4UcZc2BT2SRG2sTLhKVmpeNL/hkFh8fBqQjWzEwHfU4JBL
xeBXcLp8A0N4HCrhmq1iXfFGtHMaqhwGaDOPVSQ7PPByoNDJomsB9YUyYmUdyebypHbrqzM/sp5s
15Qg9HOPL42nk7ECKu8slV/SQ+pye1VUhqS4oobPo0Yb3e+Yr6OtihMwzyK8kbWs4p3G9R19SXJu
8EBTebJTsE/ldp5nRKIaffn4oiX2xGblPfho62GfAW6fUd1yL0g9uk97h858+0/PFsKLP5kClQGn
jMyWAlXmoDTfkLYX9A+946Er+xk0YbuyKa1PnUKCcDwAYo2chPJZWm5o+eA6f5kSoXzsGHEO35rL
TiuG02LOKQG/D8V5P4UeGgBnA8JjkecxwkM6iauEYsbJvigJR+PQ9PpRQNd0tvmyCdUHDQiinLbK
RS9p7ueVFZ85g7hp9tYXj3qAtMedCiwTr2oSBgUleEAchh/eiKXIh9ER3H31g9vRclVLXPwO+ArP
ypvJVrxunQVV/R6UF07ySGlk/081gYxZe/vxdOrBYdKLrrmw+avpiqAV9EGbNKixQL4ok6ueU4Ly
Fonwm0TOvOKPiqYLnUUWgcm8mySGVR4XSOuhDfUOFrxrCkaZsGYKm/KqxMD7wMIaf3NsXKerY2mh
VdZD6G4Mf3AKo7nONLNVbwhhKZbURIfnJYwV6zEVOMsxcIVrW9loKzvMaN1I9bT/vmCvxaYxNfHw
vxqrmzV/EuAGp/y+DqxG3yHAYSFHcVvbnMId9zkNy+NjFiL01v3YYeHoVuPgMN1pGOAmc+DzxGZ8
dUrdxaELcyrBIXhf+h3pToWtcEPueIUJuvQh9Nhs204JMuyZLOFGxDoHC02+1ISDyKDaiTRX8zHC
O1dCkrro4iI3bZEdBm5BIeo+T27H/5y6tmQAfxt4yZfiHhKFW3IQlOSdhJHWERyjIJ7f1NFWdi4N
NyWKP9Bb7Fn+iCabMMkqS4QmoMbDvMSA32+W6hp6Jf6+dwHhPbcIfA2o/RIHPYzST+P89L04VKfU
5Clggyj6SX93pnKtNZ+j/CbpX8XmN1ob8HG2gfBabQi63OAoVU0eeMpmqI0k5i9Pw533gxiwObph
0f23Yuh621asPm296X2RWwXGrW8YiBY6xEbF0DY1mOwAxd+xT95UB6Pnrb2V1Ky9Z+qnqCS91rtA
G/3ePpgixaYgv1oA8CZsYyHiER+DWb0xk2yl9rPELYxLDcyN6MK5rMGuEoS+CeQPV6gY42cbqIla
jVpPJPG7cnk6Gw7fESyz5tYmv+Pb8wVyT9VNYJGYWwTdOphKdThnHRpuzYooaYGaEBvMHxAR+dDA
OHwLsVfEcTHO+Z9/Ixh5DAndUXlwkUSI4h/GIH9SOXOGOsIPTd160QBAMwDNiUhU45Y73FlCTKRI
mlrGEvXZo2iS9YMt4PZorcMlsBAhVQMQt+c6ayo/8cwMURReoufz/Wb/gFzyLvIfVmSMvsoiTcoh
cXM7fGPkchy7JGGVPIGibqeUfgtWDqC0yLkOxNOwukk/30UmL3ZewbM4ZCNrmBJ2vmLNUlvBOzKo
2uYMYNWYN3jcbmhGDNRrmVS7gMo5pMBCjEDTJz4Bll3VWTrEAz011GLBpgndz3fJG6szYJX/AwqT
ZJlWa3NAROTmSUXNjYZAH2Z8MrE2Xyi4Iazk3heqvcQZJ7UcQtn1wDaqCGSjI0P9xNuY4Km4vdEA
v2AH2Bom2BtnzZ41fl3a1qhJfA5Pkd9kLetk5GVqg3FKhCIJbhzBng9mGcxaRCGT8KRVaJ0oYNYg
h4DGa5z3h3m0A7juJjzXPLhUa1Xi8FdT6xHl39O7wVVQ/pXRhNiQfWLopJuwFP0FRhQq0W8OrILC
82qrxymJPmyDYbeGbXVEbMUHP+FyiLzQKMHI8C5qnLF3IBfTLHff3BpdnwIXNt2AWbMrXZu1KpC+
6FMtbC6zha1kL4fdwDfeNSsCFmjVU7kIqFsU+esg7RQ7KOexT086C2kcI+Xb66L68jcGl1ZVp9Dh
skN0BoFfayx5Ac9CAyVR5pLS3OzfOO5qxmHP8jnyYJIEyUP06KfxRnOyXdKQzF+cSM13d/wo1TJq
dhdJla+H27/NftbguqJP8bdklwCMmp/M6u0oGbEpQuKk06oZYwpezrZgw1/OLRzxGWIUuE30KqkV
ckeRJQyFXtrIlQw3KK4PFxib3tsk31s5kLjchXGr2L9Hge37YYMLeg3w8USli8Lr5pquimvtABf6
KVrcVUJScZ8OALN8/W2TnBm8Zt/2zlPuHEHN22LMW05FMhIXPQV0Hwg9oJDZP8/Cbq6llL97NyQP
L/Y46bkQeO+CRSea/BjwvBtU3yLjTeGeIVoL19rPn2n88VTTAExRRLGbYLRIn3NPcSiuRdfd/I90
bIleMj+FkfJ5/jzNQBYPI0ZJAVBPhauQt7Rn4440ia5OC3puhMlVaU1LCX79hTnpKUHGnhkw2vAj
d2rftg9V4307PaJ4duC4DvZyd/DGkdB0ldmRZn4SGdT07msuLbR8JhJcqP9CS1l4tafIhfydLeDw
l9DYYDVd0fj5HMyeyzmjYR7ubmKtTa5iDnuHKY/QP9vGjajh7qX+S6I1KhyoSXNXApHwWr7cOIlP
11TAWJXmM3jfH0tkWQaNHRqZNOv1RQVW+EMSJFSnCNAWcWu2vAVIeWabokHJzB/6rmGCYx+AQykj
KkNSDFPPQwi/WR1X44CIntz2f5icdp6HQve9OnSAdf2TqL/2+ARLytskd70ogKbaQBUX7dsDDa4e
oDveliYiesX+EFmuVNMJq80YftjYw5knMYu94VbKaiAoXS9XdcfFSWv8KJ72G3SeBNzs5y9T2Jsk
Q0SBmTw9EBYh7dsL6SI4+Psns3FUl26TA2ErNLYEkIDMWeAWFp8a/rliWxXoL2YZDQZ7emphALAK
nDnzQPdWFg9be3RMmngUthBY82P0A1DNIlNpPnX2Rz15Qym7wmNv3n+cerHSciFnX8sKN6Mjyyp4
C/lqMixueMUczKLQqtfOgiXjx/gA4fpkdLO9f2rAajlwgJ8ahyiNBxxo6bMOKwlSOZU/rqjPmpI/
r1Lx1/Sw3fe0w+DsgVEMGfDKFND4CIbdeOP1gDmVaoIc6NA+Ji/BsYayVEBEqvSvNc3vSoQ1LTwF
EJRK3SWX++LSElMHIpYDsofh3/s12jdsh7FnBGMjUybiUlldsstXumGmo3WtAv/voAv1bNGeYSXY
StMziUJ9RGU8yQjHTUQJ34PNOEdkQ8IjvWaedV3k2GtW23YZnQtbofTMJdnPLR6zvsmzRegq2D6P
dtylj1ZPjXJyxkogBcwpsh+RMRExihDE8LQ+Y49ZdJ7ifuBCBFJ+GAe5+MJMmCvDqt/PuvS2eRRc
afDsFHvw+SvCE2t84kYvg7ekxAk4UBwN6n4G9m8Sr6q9T7mPxdKJ5FBZfL92u5tHYbEBB5B4cZib
IL1qgBzvrUNq/5oapV+qGyuLzqm9/Fty6ee4UYDOHUQEMh6iZl+/ZK054L3w1GNqReZdElo3IdOO
9bcqhWleucW5lynUB6u3EFAJxSGZ9yF03Z7amagAkTuS7cg1YWUEIMWhr9FazcxSML54fsxqTDeK
rYQvnyNzp+glB0fPRKFsfgBRYZhRV+it7TPy0x2IOvAsc/4lHZbIr4+ptUZyG6ccb1jGc1bk9Kx+
FFmoXUeIbqzsmsgue7h38Fi8/jDzyFMBydoYyMibcqHyCYZ4yjvN3t8ir8ZNWxQdzxzJBBpXl/0J
1oX7SaaWRO6F+yIVR43Y1uZ7iHasBrV/mgVc7EZdsNQEu9KxoG89K1CYDV9udN3ehtu2VxCocEtD
+1oVbhjbThD0ueNbQUpS8dF7ni3AFpaJO1u+IOdf0ZyW+yuNUrBnyzK2ns70ZaKqzdUMp4p0JAv0
Refi+QQAE2GN3e2hc3X8phcsePHDVOs1AvhF/7vijhXOkFglpL7tpII3P0SEADz6NK0jV8Vlc6m4
+36MXxyn8sKJaEAO11+P/LWD18mgl+iyc3Zqfi3I34s/ClAzSEsnk3cgPRPhJEEIAO8Vqup3FZ0h
W9dFcOcbtg8Dd2LD2roGTcCi0/hYiCVyQ3+QgWAb43QK4Tai+3Yu7QBvDCD/bjSMA1wIAGczhCVI
ZgsoMuISZgRuzpGqvggDM9Sn8/L5H63NBolsM+Kmu0B3h5iuCIMzOfVYkI6WhA5hoEXc0xmjrvt/
8RIldUpTIcRalYJJa0oCkfgAgeCAAL9240tFaLCWeD/zk1V9j/4HYZui5MbnDl6kF5ABjrmpHC1m
ds5/tm+lzrGyzxWfzZ+jQQElWfC0A5Ci5KPl3KjgcGph9jqOb3Kn6vZOgCTSJuJYArH9sxIJnvAD
ZgT5BjXRLlWP6r/e0q67nzGXMgF/X4CFR2XokpVEpGgp4YfhPBO57TtRWUQbYxAHA0kRIolUT6Id
QIsNav9tk+/jbia0kC5kTQzr8NChPwxVFVAXu6bc9/WXJopHx4VYeMmgTquck25hpzaIph77VQdW
FW/D06AYU9ztD/n0rb91k1WrI8eS8aicDhWONwRd0RzGEx3n+9JZOcaGQOtjBPL8FGpafyj/WmdX
sfT0JEtbCiKVUTYdi2QDdEac1GvAEmnS2QFMEfSixGypIwbIBwgXknylesvp/4xUqg/WufHUwj0w
e4gmjwKNAUajdrnW9bY2TFhb0mz9Tar2XiOe/eqEDNj5yN/5K8f5+4EdbOwIa65KuDUTau10H8ja
b2457tyn4oLEArx91zr4xtxczrEHrg7W/FJ0umNtbzInJA5g2E11UthnTN7DLYxVWNT6QfkW1JKJ
8FZq5PM/MEKl4nLzu0C0BL2vwDDv2stXhAe3zMA8J5gUVDKyWze14LClRdh9L53WE3LjVhmfdAOF
6/3xxom+CHcv0WG6CxvL0v1LdOgJg7oO6QfYeTeTvlqxH+2ZQ+p7lhECgEnba80kpyPSznzQ2PHI
qydk7wE0EAmCkp6HNhmTkGd1lKCjQknQASAKdYp+moIDK3YSI1weUA6lUcWWIyBNywF0DmXD52Gt
1livdkBnzbeQPlJ+ew8kjuM2qJh4XFpy/KCdM2nGDyCmP5AEvnTIB8Spjd9gIE7I5+JykznLvmbZ
JZQO9x92CrObqYpcIZaEk6g5ZtknUWUqj5/CDnKbUWkskXWpo3o5A8TWY3xe8KlumrMTooqWFzxr
OpwzMF6+3g1qb/5HPdOwU8qeZg72Xb4W1AZDL2K1cSU5nYLQskcuTLQwEAZyRAQhB1A3uBq9UQ/O
oLmnp38GJdbH4RiM0W1t8zdt8sLu7gdPtjcKiECso2AARO/oOyTdIh/HWsal85zv0MpMv6Q2iur2
4Z+onU3flu5PB56/bLtt9g3LTOOJOWoczPc5LLYZREOfl8AF+qvrsN3CSeDp2rjycpXe6H8rphe7
iz7WCeJkGdMoxm3xhWn9e+fcZzw2sCPY2eoPCYFL5a5R0eXFbjJ1YYAQhICmagHPV1CGCpADqYHn
Nav6S6DNid/W2bdM79riFoacawtvhKP9ErXUFbTr1WOys5C8/H87LLCUqjMFcGEho6C81wYKsA/2
x2dIAcXPRGVGc5zw/sFVmptbsQrmbi6Z38TgoAMkbcKscnOf3TDvQO7C8/7Y1b1jmmKIzpZPwiKk
rwswNUjNBo/a3BpYMYcMgfJTiECErMZegCZ7PWUp9JA/FDC4RJ/Dm17jSqrrrGkgGHuNtZzLtkWO
R6ofJJACsJkM36EeXMULphQMH2T2vUZG3cRKFFNgTspPIA7gars2VMvUVK46XnUKdtkOhaFXsIUO
FnqDx7cfopuO30r2vUafaFMMG1E9XwziI8WRmoCg30kDh5fCeeEWgMY49jjXB+D3ojnFWyDoFsVz
leMDhes2nGwH2ZR/qIIZStYLQJxmA+ZSn1otF7XDpgKi172TPsDMjTR8wNqqERMeMQiPIZaX1Tdr
WiijUItkVW54hjZ8XImUSYyzvPFP/L6owOJ3luvCqKfOgLe9LT8ggb+wItYOAIvxhmRju1G9zZ44
+kMNLolM0dPWlr9ovQv+a2w3jHzRMdi9pKhYr319SCI3gXmgFMce/rsxacFY223YXc7FZsW2xFCP
VR9JP5wBatlm3/ZPYLvypKanUHEQH4IYq4YswmXLc6K0f+jNccxgsoT0oqRuj9+n+G4AzsIVey86
Dj4hHVZ2QB8XjKHy6tkYskoPFKzcpS5RcZjkod+E1hlDyGrmjVEzst/nirgdnsKilYT3dtvDQaUp
kcfonGMvzzWMiy95ae3oUlVIbz7owsx0Sli1JAua0G1LeMMjwtCf2nLBB5HvrGyKmH6nMdQ6AZjW
Dh1/zcShueEWCioKTNnqNftTl/B7IN7rcxQEYZb6XPpiFMSXU9Wjd+7Uqg7mj7pUqBQ2S8GiYp2L
wA6uUeJmARhsDQw3IEFjDx/EwAFfDtt5hHvrSLiVL+c2/BJkEUH7tsn/zqGN65r8YtfH0/j7gN2e
4B8VIHokNzI0sh0yXj9fU/M1jSweo4ZAa5VSfv30tZksjr3MO44dPnaOgrGdOgpatLpq77iKqqh2
nZUFFFhFhbO+63dSYsISDqI/z3ez8rSVlHQa+grUoz9Da/rFxUMfDNjv/9RIHxwZmyNTSYAxdsrA
vADb0vCbcdsFQseoz7xDxQbAh2T/629w3Bc0tCHy0DVPXXwFXOhGZTBwx21WpbJtL9ph1YrRkjfj
QgGuiesK/LlzfIawu2T0EQa3FsJPSZt4Gq0UnR/FwXuyaHoYuCR1zYlqmHXGVrYnzTbjGCTH18qj
NLdQutWQSQ3FXtNebfrNh2FgE7C1OjU8VlLAFvr9Cg5lsFqVFSerJvMZoA8dzDXMOpSj0ZtDvhKX
lFEQipHBHJ2o4+KE7upWA4PTwdpxhpc/Q+w+GseMFR1iVlTiX36ibDuu54vcOe9iD7fTo1Fad7+T
qEf7f3FmLosKBrrmxqfriFEVYjemxkKnPr3ZZcqa0TYXRZ0AQZVrn4sQKxqCJLL8HD8yWjSn4wmp
9xMHoEZEZ0S+VIYCZgyVPfNOd3Wl2tGrHUmOrgH7aM3J7mxj/8m4/kOLWi/8mOTiKVvpoRy+70pq
THWNbtHzXeZrpeyVsbTqchtvb2Y+NzwB79zsRcQYrbH8lXmZ8ZFOL90Pd0R1yNihi8SOCBau4Jkm
Izs22HFFHMwpokeqwslToLJCIbvFSDC8fWZp/TfVn1iDMIOHEuWbjpkCe8rU+YtOtzh6uZbUzwRO
f7IOG85j8uy2bY946bwKHhuKq8rtLnku8gG3gfweVBCGwUG8I/XT9mCmHmH9I7tS4RjvM90U5zWa
/AlfBfPc3cfYl2jaGc17pTltAdlQbaPfC/5laYDBzSkl5a9W30wxw84vEPox3TlqNgbYsQwl6RCb
1ONEIFWAsnr1gshA7tvVfiN47cbBg5vZMCR4cqevFLQe3BY5tStB7XF1MZmW0oeH1DaQ+y/iOMRv
TCkFJ4rzg//a8CkU3a/sCTWLWWIXpL0aTF8JQ65N8E2Vb/w98Nq9PBXou96ntUyZOOgdJR8H4E4w
NPxaVwwcAGbPGIoHi28mSS7Rue6KHgHr3TqiMzeeLeLZ1hDrCj8tKtPrqWaQu91mDzh9BoEBHUA4
QKFfI9qxc1AiwDBJaiRqCZIvGhcrw+Zmzq6OFp45NQ2JQ7rL8m5ANNdnFI9le0gxvRQpA87nAasD
pbWF6Nyo5OkjbJ0KM930sPvRf9L3bBh+iNwreC7D2hPCgjJYC/+YMeul99tGAQbHqw1WbbIfHHAr
7D4HPtfOHhnJC5lt64tFiDweIcvD2HKxOHnaFpdW5qHbBo3sk+BKiyElunBn+62sOA2lgIk8lxbX
UsXcGLQEPaUlaacJWI11t3jgA9LXfZ3PmvtulH0amOAiWKkn0F1fLV6AAcGIA4iv1BtKF1O0wySL
9TiTkF3CMzoaLenVU+U1BhtZO0Z0BfVCqHBuLticg4XKDat/fpD8YPIpz0THzfqqxUjhgXKwkMdq
ET4XudbcTl+70GnazqeG/yVsW6I63NvJ6oOaSmEC8cXUFPIiIZd86kZhaJHVzO7bErfT2nQ1kEqi
8QD0lfu8dyYNvvS8psodvDKHvrcUqQZvS5UbW9LpuIyXyRyRdgnSkbw/Za5KC2Ve4If0LWGUfgl7
xXbtfmNjILGnhTpa+Dn5aN0bvkPULL2t4hUtU6YuER7MyACI0GrIEDZwtXLhSlB8SM8PEk9S28vh
4X930RandSCHhPUTR56aG/stEogFVueJBJ0j+Abmy4SG7urGxQf60ACGV1kOe0AjZmz4iTlpH3Xj
eCzGLCHlB9eVDy6ZLspWG6dlsTLQQgfl8A/MH6/Usp+UtBqxQwIzjYTcnZ+ec3jjsllee2XCYoaP
lbK3Z3JNBSdTX/3nhv7H8wKUNIEC7GZDoY3OPwQqdEGkGtib9fdjU2zKS8BLuVFGk2GpL+NeILVE
wB2PoJWfknGBFEf6eYKck/DYdjnxdT6boBHWz0WH/dfDaiuUBMvSVVP7dJrzXEkBBscpWE1V6qvX
KEGNGsqRVALh1IsHkzz4BV8+4uSon82envDeDJ/6/uF7OZaNIkcvw9/LDwVhyvnWtGPDpkFbbFs7
h9Ryo63w0ZlK4mRZ4u1vHxev3yHSKAms8EgKPrX1y7MTzlAv2DnARTE7EkNvGz8fDcjaRhRI888D
Fofuct9WoCRY6tAhawkIOzbYRPdUCauVx7dXXZ0/jmB181o+26gN6Sw8bCie6Qeh/3BzL3+XX5zV
ImaVgqu+Qs/7DGkEvJMcq49hC0bwNB0AnBg5H5gNqBMmLSAQTywjpgmkWfi689WfJVffpbkCDoMP
Rf7NQj+RaZUgWLde9tKsJcAzbf1TMM0Q0GP9MyvzTIoMup+Ay4+sSjNPt0toBLdXy3CtvqwyDnzS
viEV0RNexPjtHi67twXgvYp3u5lVtSdOJGwswhNhdBujFnuozmbTgPbCK3B4fcXpRBcyyEnNP2G8
Fp5hGBpmXBoc9WQ7RPIqo9E0mqYUOCC3cPlShBl23B2IzqwUkE4xu98PPAMHWBaHeAFgLCGpl9Om
7hbXXxgD5n0DmDQS3Q4jHhXO3xWEZlNeDm0mv160SxCSj8dpN7ugoyVih2MfM4mJ1Z3pM/nUuKjm
9WXfMKJGWugieoiO1YYEwbPNp64jP94qlH7GKJZdJQNJ/EBSwfEcSBwLNVUlPKJeBEtsXP+OtFy0
ZbnMNKLYd35vPKq48TMVO6J4QSPeDIeShiKlPeP7RXdSh+0iYuKn6xZGtPpeZGbIu87lyZcW8LPA
w/fFtm1SaNfgCbzlktG8SUaG0uPVI83+BAFmsPauNAnvAcAvYL+GUdLMM79vn/b4JEd2+B8BW5x9
HycOO6OCoBZapVCdam6fnMcwjTxqZ1pc19V3eOHiHaVDCrQ9Es8JgaMVzeWQ9yJSroA2wSOzaWMf
oPZCxba5UMxmqiiT173fiCuu87dKALzc2InGCl71yNUEa2BGBf18P2V6cyz5BT29tnIuB0VHVfLJ
7jJFukY189TnJxE5wQjpYFq1Op8PsGloafb59DK5OoS6S8gYVYZqHny3irty1N1SaNL5KOpifOR9
IbaqUqDaXNHFoPGF3KGOQtYmCHgm4eGiFpV1Yc9YSEutM0yGuDpvL0i/8rIR5Yx257dmTUTRLWCW
CKPnbvUwEvKkzHbwTnThDgqSsJ3CdiL7LraPPCTfR1QjUpq74MFjXK8vHf2ZWu01+N2pBD/QMJw/
QTfoLfkZZ3DUA8+qPUf2ZtEMHqoynw61FLRZ3kk24wjbkt9fIEMvKvSSFvSpIpEcX6MNvb97OZr4
2VdAzd8Zt5+gQtB2rVjOArWQggz7u5aeuMZrP9lntbAfptpnIYWwhzAEYNXnO1hal9kL8qSL2Dj+
p8CMaycCSMTLKHdz6VJ1/A62KlvEnzoFwcqydeJglSQt240QqoSBnowu3wsiH5RqtgtohEh9TeNj
S1i1CsNkxqE1sbCoMk/ejuGKZdty9lDO+iX6Xk33NOT8GOUWahXvDx97YO4sYCaDm7w1aICK01Ww
/3FhrRALML6Uajumx3UjII6uv7cLkvkjuXIsVvLJQnjUZj08PirE3BqwFx0Z4zioBMFFOn/ZV3hR
3gQp7QUQ6YThEg2wYj7RSkK6j+kfe0ayCjtNEdiTIm9FwphoW8SVmhxSllE7AyzHh0ZIDaOIvUDR
4rrm/DlAbjKD013hDPr1+XjVGaOWdrvn38uMHo/gN1PKlP15icM6vx5rbdox9y5p5UnjLGHm4LNj
s24DBSICGgqUb8q7t6HeSObdzcZ21dRr4sSs0RbS9g8qZUgdg0dK8kKIZ3aitytHyWy8gjnA2nAG
F40kEHIf5WKbCcj45u4oC0RGl3JW8xFMxb32sIuLRSMTwPp0CARFJqm4+OGB8lO3Zse0Czwh7+K6
7sdd+26nQWRgRS8OIrba27O5zlKRU/HCY+rZhx7YWPb+GTT6PjVhgcqaTZc7br7Wrn3+4dnkmuXx
pS2eXWDf4kSz44sc1IyUUU4VlL5ict0ChCVRE46ii1tyXfXQycXxr8Aai92fy0ek78rOupa8htkk
jsJi1lfudzBL8S82JLISjkik7kkPt1OzyiPNXhTiTg24dGJ6XnKySWq785/kOoVg9u+RDSOSN4wF
ngSQxQUx4wtJ/SxSnRTn0d0DJ/yhN1kccG1417GqMNOI6A37fBnYcJhgDZ6gz6cGvC4bgf7XgLvn
TF1+4K6iY2ev2GvYtsjB1xKcTaEaucqkMYnRvuIzPBN/yPonFJXtvIcl6wX3p6Ry4LBTFnJRwzXE
/KBfQUpy7DpNqq/s7SxZUVrxadLkedb/AE/co/Z/k36opbgq7C3AswdYKuMiBbs8q06TUSW8QTfm
OVKhcPv/01trPfFDxwJKkXWmc/vIi2Awoeshve0tNARaHYc191fPKUDG6jskG0bMOACcChBjgn9Q
+7rPOkvJCRPX0jZSCu7ZnFu+3rfO17AWIZQX/SFNRuilqVWZyQYDcJXkgSQulrmTJPfXc9LzOOBo
16+krUSW42X+53HdRobWMBgFLSzShEF5mQ0rzailIpWAstct/bCNPGT/btgI61PQFd4nHjxBeLTv
7UZuwVQN//Z+2d5SlTy8B2m1oyMEstlPWufYf8kMlmlZhoPGDTExacgWweyYutowSb8n+8j8X4c1
zxWfGs5fAj7BvBIss94fRHJSz9QL7OM4m/pPGTAgfzKUvP68kVxPNBbWzq8LWEA9TMa78uHGDoon
MMD3B5bn8meyScg/4iiAa77yvy0B6XtquzsBNS5Z5bu0Pd8onTvyWVPTEItLjVXHY0ypPt1ZGXWp
/tfYVg25yo8FJiSrxNvoEYb2N5ELop5BlZ0Ifd0o5XET3s7h6mAmjO6L/xa0o1eh9x8ie7w6W5D0
ZoiEbAz2yiCpCNF8Ajh7HdzTBcnGHauz0aKTVxsOumIdTjEXlwI/O3KUbvaWJ7Suia4Mv1J9Dw31
HybG94GTXB8iJow7SZptTxnlf7T7Y6lRgsG6R3RrC7V3I1FaZIzxIODWGPLjAmBnoIT9FMaBE3pS
rSKHh7t0QgJUMRMhJWKW3/uFAAJxcxTLoTZzxANcz4i6Df7sgVLq7oAEx7/L+vIvEVzp7wAodRVa
HEToEoLvPMxHYpayxmNo/de00HkTkvF755jsIf+4AwhvEFEnwqPaM/EMGzKo+KARSEvVDWnX0oLY
Q7cDKPSY+xk5nYFP+heJCcOYX+GaI2Cb6mpa7sYRCAjjrrrxj0t4cMfvpZ6xbN2IMraFldRbSE18
NmNi9zHuhZ/quyQ/RGALKWPUwgy8keIHUO+ceEHn4FFxIhdq+WHHjCfHCzOm4oJugEUjVGBbjZs9
lg+cHR76WenwYPWBHRm4p99NUPXmXhJFpIg6tcn0y+IhTBiBMHTiXjAnMSQNB5pD0e3isjd3N61F
2vACPfxtwvZi1I8dm+Jz872ljwuXeBmEM3Oh0ECHZSjF8R2ZimNU9N4GoEz/dT5n7xn4i++kzABD
3mOBjzz6S2/5n02JuGf6KazZZlvLf3f0dzxuJZgpF+jq/tLaqyazXFuMyFiqR95Yme2y36WDQJxC
XKPmfzV2Ohh9BF+oSbKGWwKbgYdaB5U8bRRqXSEFR5/3unIhHy55GQT06cn5NSFwgincnpWlpeLC
LgqxmEddLQUW/sSe/ggdzUT6ZqVG5rGSuTb3HixjKZfbFgEp2rco0sP5IJoz44FWEX8zl3RCdFeP
v8cpoWT0Z2bGS8Tg7fDkhkcazPb+Tu93ods/JWMB/gTwU+7rKMABAJT+yC85p4NgeML4Ks+10ueL
6/DKcSiGAiuinqai8n9gPheOjLBfjoaTIoqmBKUWCMasDhxANIKaCRop5YNQm35kGJ/XBvsKo5nz
751/foO5MfZH+jUOq33HYWMFmZBqvsUtllYpDLwflzdYgREZ0kEzdJ0K7SNVRzPtgmoN9yOFthbE
5FIn5cJY6skVcjp6AJaA7lSBo2GPNCCWUI8qJKk3uayA52WyTDCgY1sPJPiGUOiBpk4Ekl+fR97N
XO4riUmqnjf1gp2nYnwQRHQ+H3HMLHB6R6UIQjsLr8Ou9c9eD0+BAAZ61cDgnjGB1LNQQDO74I2V
ZCniv+BWt69aq6PRIve0a1g0VoKmIjtYA1WpEFGYqD7lBKKhNBKZYwhC0pIouorxtXy4+79RAdWz
KRsCiKNA3XchwZdPtmT7q9HYZsH68NZ7gMjG30PHi/Gid5DLPCCC4LXGdB4iRZrrGcyNg4nFH6N8
h9f+IYYn+ORvUsr8LVwK/0bQKgxnJt04WSNgin8GtwMvDLLduvTMSvfckdF9A4P9n2Ak4HkJ/DI4
4Yw2oFXL+lazFuO7jju0jPFQQlcpAwhSp96FjK16rXagE9ReQvAfCaDZC9KkvtTQeSIsn+OH2y0G
OZ+ntTcHS5SB2/wdFfme5LWqWr9DXfVuvaEwtE305kgAQ1lYNlE5i33g+EbRttlzyCVrTDeg3ffs
XmrryrdJrKP7zKvz9K9Wf/OzxPjDQxBktu4mVLnz2Zp3r+k/qj86Nzi2qMuDIm8qavsfSkby+l2S
/3+kcoeYnqIEA1C3et6G0e7XIQBF9WzDwRzsmKhDg6DT7IjxcOqkRaWmqjTRCCJsLpOukM1bGhYs
QmuPLanhjCOs4OqOOFkfvlunU6J7SFB+izwRQH6pxqb1uZs4BcrrHXIEf3gF2xqVhh4Hwp4U4lub
AESjFoNaE1z1f45sdFE3R23IUZ2t73roY9IUE8QhXe8ZB/FSrHN385eJ8b5MGpmd9+Tl/lpi5hNX
IlQqJkwIIXwrDjNHMsit2GzoZVbyK3cXOxKCYctP+QNqv/2+AeFgt1SHp9yt9tmhwG0rx8BF2PLn
Nm6k9R3r+e0rCtb+03zkwb8YeWcPBtQPPjkJXCiBLgBxR/26ldIy0PSU5KZNO0QrsKEbfc7RL/Hd
qdNL9Tm8ZpXXSSMguJQEZ6ijzPIIBf7k3jlN/h7F0yx5FjgeE1hWoAi7AtCnauub9qTfc0xNmw+W
1jy1hzHhkFgn6UYMMVrDjYmtiRp32NFl+7Iq+3ZdVj+cEwgfaEaA+xsm6P8VFli2OGoWLS6ujN8Q
wsfdb99sUq77zq+1L0fzOPqVdsEAXunNXcEDwFWu7xrkNpHayx3xp5xRm13Q7kpCNcLQ2p3V7gkk
3r9RlyIkjy0manA1qtfQeCuLMFQv2og/qdfu89bHc6TEDUJLDfUFHW6tdWm4OhJVqi4qC09zB4w6
5/lyRxWW2Waf2KLwxRqh5n+OJVPKprs0QRevdTY4tJh1AJSmdxbx7dvOiWkTpLEikHGoZKFbHh0I
/96BkTkgRcLPVVEUx8l94ykBaigJQzTxqq9AeNJaIV5cU6Yeg3Pmp+Rss0BgzUkXIr+I3hIRvHMn
cgIstDXl1y9hmtbLtoPwdaJ94ImUQCGG3O2cYijm4AAu4oC1JZQAzG6k7ohDrom1+PbCPoUAghiX
J6lCnn91J8lZOxhkzT/O1CDxDTngsbLhKnm9UbfOn95TD0omBKZbtiuJXJtZ4NO0J8fhiqJfpCF7
c4hcf31SIdZCa/HfsG/8CjKALKBpQnDXU/+YFIGQJT5yztJhA0HP/KfL2dMTXaDBwqG8K6QfMPzb
hgNFwfTleA9QNUPZfadSiQOXF9qUMWWOTFwF2EMx0twVvj4h6JnG82uI2zwQJSNA6STFmiFDrKc8
LyGhUEJLGepJU3SLJwrfjT2JlwxDsqbdRPuKbtzklsJukT32FUiOt/QRQwYIQDjVXS/CTF6aevEb
4IYUDioJERrSrmTFy449OZO0l/mm6bU1jGMtlJK9AHg/WIO6PrGPsy1G8rYCMDNwkCtp/DIT6zeG
fTncZijQhduWVXWRl9rw9nvJyYUtZeojekq1CULrKtc99q3NhzxGILKCcaseN5CY/SOGhMdm3/et
doZMW5hbRKKrC6ohwb6U9elmf/zOjR1ZyQwCM87uUcJ5Extg66pwdQL0XhGnT3U3dAgkjb9NXvcC
Y1pPZctKwQK2B6rHqCgLVQcywtir6fZYv69W0ITDhhCkQCeeqdYJGXDTMlRzbZyKIXXv+au9jTma
Twx5ypNHZnydcDlalkmGmxgf7kjefDw9ZkR7jVqwnBgrdBBpfeBV0/ELplEKLaYcuTj4sLTRoiEF
UudLXmd+r8nP3SbBGAF+e+hUFjUAeYxni7Wovnksd824QgQgqBmoic9IpZzAnj3mJmN/7pwtf+5/
lwiT6pRqhcpTVjkQrsKXWqrJxvix+hl1gF8DANvJmNmNrDFLUgf3JObnY0OgOoMEYNuine3ICydp
/rBX96whlFAfcezuxTgaTbSHOD6gzGS2zHakq//oBeEVnWQXpbNxityodMknh5/0TPxVNGs5AfSG
uOCiq3Q+AwK6fBA230EtNTv+sk/My33ghzxZbrfqTb84tNzntvqlj+jGOGOoXp8/RFVqPQz3vCtr
thtqtr44Rn3KrGng68A+ZT2dpExbQq3mTUBtP8X8t1QmDRmAhLLyNQGvs9TEFgt/63RC7UcyCecF
ORfApvFsE8tri7kvlm8oSKLTLZNTKwVbkjcqm/2/DxNahki2fQQN0BP+6/rqUXZLxE9IRMvXifQl
fu6KSwkKgaGKv/7AF7NO2ruJysvzxRbbKpStjx5PAsG5YxeL9sHIT1ITFrvOQLoUXhzAK23/ij0c
tIJDXBQXcx19ZLK4IXPoT+IxiPvL87+NAW7e31gamYJR4tQmpvTJx/HVvjXs5P40as7CmqdMyqWn
bxAb+WMm0dn9l0DQd7qnKX7Mf75Tx4uMCxbHYf2Q+iP0CQAAyM6e+PlwIdqqSP8TS9aZ00x3V+H8
DUAuSMU105A/jOmdkgltaFc3azAMIE3X28GckP9baGwrizwzQI+f6PSEzbRAhcYA5hu3UiXJFVRd
YB3mJbQofgXYdEJiI5PYWCE8xHRyE1/32M584tCSlql8EiqLmr/GMxIRFrhjbGCGfRyGY8EhLcJC
nj4PMCtdhH0WbRujC4apTfav1rnOqipy7ZVSpyv2ssiLuhfjVcplIk0+NhgNRbUIWQCXQHjZeCmL
bXfnu9OyLkAe07oq+gMo+VZsxextTTZsZIf28nKMkY9f4WAT66LYsZ2Nu9R2jL+n0gQxUEpLfqKa
jdsI68VDc2KiWIVgabVOtQypGY2G2bFi3OHhwtt6jYOTzyw0RuDzZe/ZF8D5GbME7V7esVaOTcvW
gPmx3FafwDNoy7Q66vhtFXSNFlwG6cVuIY0dKQulohJb4fK/mY5eCJr6sJVo3naUncos73fRltaN
Rfel+bFmEc6x33oRuUDqmyQWXvKpvh8kX/S2X6CWYbtFsEpmbsNlOyzVJYy4NGb0LnhVboG7wgHN
B3Q9QNw28didfSLNaGOnmVZ4dnYN7OJURNjz/B77my7BpNLF6tmfNChW/DQ6fDsZhQvp4oiaTluG
q4IGyy0+2TgkfX8aYMJGX0NW3ZbHsomfGS3u+NuSc8btBvn0ODxbsGYL40QucDlr8fZrC2npp+C6
Qz6aQn0JGcbPq374ufQp8tdiPFHG//HsKatR4RbntWK1Wd2iMgyk19LGykF0ilN1H8BFP+LNJHAO
LhEbVcjD9lGqWP4JPtVgNOdH3wplaPPZ3+5rBGt7DfCzNPV/w4TB8M2f7Zx9T10LikDW9mRCqZsz
mwdsp53pPTpSgdLg7gicYYG02hoZ+DY/+pgdyV6U3VgkDFGdQu6d2vAJcwtbKrXU2KRFV2+Aqxza
xukLydy3K8Kr5NDvXiUKBLYRKtSWGBFksRuFXOt0nqh2LfbI4w3S/rS5J6amk3SD9EXQ0rNDmTsp
eeXcWc9Evx15NYOImZQlTqwDLYgExxA0zNBsJqeq0ivelLFB6m6J5mdQsNXlYX5uKSjP7WxC7aFo
PifA36pD5EP6bSKzjE0avaZIA6vuh+O3v0UzcjpKXmxOKrq033JVE1uv9986uoFLoJBmQoTF9brs
QJhoIBJUWR4+Qfms2MblJMQ98AaDfrmv9fpEj6pRmW/L2M1OPhZs8QDQPLSs77TgXD1npMa9j+w4
E8KmUk05E77jPSg+zAM0CSBXec2erpLq1L/irHo46MR3Gy1YHp9BIl/Z1jm7n8H9EkUn8m2nfH9K
7YbrJN6Gl4ET2WRcz1sJ9dXOkLfvXZQJ/F+PzxZTymFnWBzlptaA9zz0/NPVajdlt0o0BYDTerG4
6dWobsfYtYopiDskfRXlFdSsLkDS6ymkhrZ7WneSxG7z+n4F+slPsHB0Tk/ZBL07+VykCL9Tt1Qk
Xpj/ueV1TGKVsLKumFuNlzwC+sQ6fGbhl+eFTMt6zKVkBqHbODVzPSTYtyublS0lKoUVby8Xb5gy
xzfiaoY7+tb5EOfZAnPqTMCkLwyZrjinb/paDkBxQUz6i1q3XClJfyMIR51rQMZUjs52xb9IBdTR
4G3tzIkQCn1t2HAbWaNylwwkVCqNfUVOzVECcNTYL4MpScgT37hMxS2eE7I0oMuw/s3flFdM2VNm
mcnIz3fuYmY51UYdEUIH7ZTOYdbfPXxBij48oU1gygxGxcvMflp7nUzDfWiwWchIdPxNR8LV2UKA
DzavEpRMAcPy61iEPI3dvWazOzKVit5bn99HYj3ahhRYHyf+06vEivZa2XQlNZ7y+mnDVXQRPVsN
vfEiO6mWnz5EnPnsorHcCa5ICwPnVK8Y4+gNMaTNIe+MqvsetDbKU7EXbGCyVGOtDH7XRQp3P6xt
Be0y6b/NODagRiVyjf1TSUibfMQcC95/YMJK1GvsLCblj3NxTWqiAxX6R/ZOnWwgkY0zaQebg7eJ
1xIYF3xn+Io+0QUs+E8Tf1hsLaOC2EZwVuFwZpRAN9wjRuMLEST3df5gzvUckMmn+/w9y0Di3WH2
KkxGwSgWoHaRGRrq94NppGDigYFtdRtXFd0JXCIKw4pJmIDviM5ew9CuRv56PrARQnt+CvffeEWg
e69YESdXrrh6Ld6lcB+xPEdqXVtnNLtZ+ol+zKfiNZyCCpOgwUamZAN2P2M6mP0HVc2e2hykAqQh
BwDN0dakZt4pRIca6g4CMoREFOsKsEXQZGjvqwA2gSnN2VxU/JcZAEj/kaXmM8BTzQILykXZvxpW
KkRlH5so6NJSIDU+ck+C3S5s5biqmcrkswmgMtobuyxd/9/gaQS69Klvn/XVtNA5j3jtynLUUhWE
TsakulMqcytsStoHc2mpzst+oUWES8rTeAb8YpBflYy/j+C36eAvAIvpMpDsymSrfydb7r0h5xGA
6Cd0ZNupWcrxpTF8alSFDgflZ99fBW+Tf/i/LDeChjvNK3fs+egrH632fUSvoyDUzFDSZn3VKRmg
aaJ6UdLEPAl2+3JLUuilr9UoFhcjZLwq5J6EI8gnNrjT/s4ujF4BDAFohH5OKV/z5QnlQ1V91UnR
Dk6/JqYy48PqxI7t5/6zw2Ag239NA9jPgAJ4ceXLZhg8pefoMA2HZKoK9arO0BYMEeUgRtiSaXOh
byWB+LnZ7Cls0RI6drMcNrgRtNNUdRwT1yGTvbON9GQ6+H24LVJCW70muHPjchH33gjo5CyFzwB+
xRphwjDDF6F1EYFwFPtwFhvMcq9wqKKSJVCtZaJiDjReFGh6Usb0c0E9R4G/ZEZv5fVnJhxDPCDv
uAZRmvyDx2jFUL99vI9UyZ32zD1lW4tTKnGXQ0P31Gar/SjvpF2ArU9qAv6eyr1TRXoEEyuTEbq2
BvTQYq3BAv7pbKNTh/24N768sLgncmGmS3mFtqLGzXMNJrdgHguQBiusOwJBP8clwCGePrUl+OLz
AY99tRdCuRNQaxpYQopnmQXy+0e+VXxRUtxf3NP8w4VPVyNqztWc+i5S1wgfyYmlsbNpwV1ycHwM
sQKqERB0gbxsdFNQqVTYqWVEuAcRGKAvls1N/KCb07vEEi2rfY8BEeoPCxjs2mOEHJZy+RU7lRR1
3j9Hd8HvmCNN91q6p0Cs2AXgeJoRlwgvA8XUxsa/rSFBBMcK26f4W7Ccnbyl+da4ou9B7m4sPTOF
TWzfy8PHVMDTtWhS+uEtPkRGDPTt0Ut0T3gV1tWpAy+hA12AGlhiL8M3fcR5GyfUhANEjz84Ok+x
X72YSEb/bP8sNNQSefE6jJ48yQItPX6EYoZtwdL+XJm/mBD5WP6Z+GAWYdiN9eqg0vwr3cGYTzPu
OOL/HO9gcCFVgBdTsYgb4bapcd7MTgTjdv31opYwOcUjHxwEyyBsRHXARHdls0YIEBOZKeqigl91
8NN5fl6jI7g9E1bYG3UuEB24sJiz2ARObU/mWQc3ZZtEp87ywbbTDw/fwCjl6fUqaUWyvWvlRQaK
BQ2r0/y6skmpokcMIO8oCKCyekOKM7DbQxXwRUFZ7YHOnZBPcgAaHMd3DOeYZQou4UZLLIKuDk+V
KLZFcFYBKABZqfutfv6Ydi4hF9m0JDPTiSbITbYOuqss60TKcKOfv5JB6l+oBJlwVSY7hSbe130H
+Be0bd6+A/HFlgt4FK0c1dLbv/XfNsH4KXkeuQ1BXkClFIthV9feFqdeMmVEnAePrhLw0TRMLry8
jcsB0scZ2M/CjQplUThJP2DNzZ666MnrKd/flG86MvB5AwxZ11N8SHo39Wa/L/Etk9WT6vzEhnrM
Z+S6w2rpciWo4ATrLvD+dkXOhPxy9ZP5HiB/tYLU/V/LH+6hrlsL+OlL/kckP8nFLl5aZWoLYYG2
+zVCXltbNlIGfTB11mtXEs3jkdC0b87aEVgVpNUapsn03Op7jTL42fSkJaInRCWSg/lf6bstR2P6
f1lssWBTibxmsrx6EyfzuvDRwFzyCfOvZxPz0scJQwFic2KiC5ViV2bq68MoGjWYRVrzU1n7j9Iw
XRS8J3MJt1Ol+V7macvNsGltgKdwC3E557a8T00D4n/RBhs8mnOahhvYAv0kk8ps0JCMgFr4KEvi
mXx2siURIOjD3Ocf2oo0YX1ZPTwvpD+J/dQ7fKOWNwiqyzlB0dmjrVdxST7APR+zGLA+i9+voekV
q5DdyvkAxi1oEYvrxdBb+ghAkU7YUA0m5Tvn492tO0rQfWG6CA37t1NJjUYYGKiQkb+77BUZMaxZ
S8JcMKyXB4XWs+bzkHeuLZCHzmrFHfbi6sAWDPWmMz2JCVIYSvj53jsQTxZeHRcsOkxkReUBgtYR
R/noMu01YrfFy/MP3hVJ4UxOXfJE3XWd/rZRWwMDdLlXB49ByG1Wf2IhYwc5zKqWC8xzi7q6R+EY
bjRMpIyXXE3mmzdAjSnjCG8RONXEG8SHqDFyZYPyaflCMWI8u7U6AWQVaZE+4MzkKucLHqNBN8Rf
Ggnf5+9EypzPhJzAB/2Dtx3ljopw0zBKDPnlxh2z9fellV/Z1sIl+IDwDlRFE3exkFU6XitMUVSm
aSgt67kuZM4kSHvx7ugonnwm4v4for37O6Ej5EP7iAuQzEdfDUI9XW6MdkuM1Oj6FsHbsZUMO5GL
wqdav88z8xo9Fi9eWhguPmJnbVEnGHKQ9hwwF6KdML5zjx7NayA15Vm7BY/JKFIBBkJ+1GU4/i7j
5blxC0C3VP3Vu+QIwmB32E78cgF2+JY/xecJqaFQQnFJp6u+EXJZhCdl111CKD4s1ulx5xYl3zpm
EmG2vmUqd8cBPXy+oy2nc3wXfdxgTxFbBpg85WXNCvxutwTbGq5XbyOuI5O9Pae5Rm4LSFa7aCwR
+MKSyfEpp6fWBZUk/6xs0D4zsNFet21GGnA9PYsYvQb+hdbQTq7D4+qBGh8oq+c2Wj+uKkF83jPh
9T9qKSVlCZVZOtPDK3SFBsAYqTQMXXQXiTvT1kyWclnyqvc0ToRPFygxdMdOSzGbM0lwSOnEGWje
8RGKleiaJRfvcx6GSEAlJrLxGK+uJxkbgXnBM5y5lZFHn5pL9KKUk/IFyFdbK4suKZShPsvNQf6e
CLrj9WPtHZGtyZjhXQkoRp41bdh5Avv0xO5z7S4k2lHQHtXvRPsATtSFTAJAZSiQYXyGrpcluN31
vwT0YiP5Ok8lGvJ1R+uFw5bZh7r5FAwLJlGiMB2N7NhjBUi+/6mH1Qp08OsUvAq8iRFCK1X8Lh2K
wRnBLIXE2oL4qkkRXp4wNDku3fYlnjSES2d7AqVVmhrHAh5V1ybWWh1ZiPw96OwJRrVeP3IsK2FZ
9j27EZ+wLWswZd/1UetaJ38bpiVA64VG7hz0Qq5i+pGtnpT4fHJJ7/ErORJGoWIJSQu8IyMD95ZR
jmknATi54Cu2tkpeY0qgSghG1wMkSYV3t6e781QNjPXBBaigjl7nEKRGjFmn7qhUzNgMhnU+p6Cz
0ToTgAoLS6NFnlTxkyXav6FMGvr+hHeSJl/UzhoY03YtLvljTHlkf8NTEcl34yrkDe7hh8v/nqIP
rQ7E4Y26q7wR4fBFTc+9/omyLI/doUd1SridoJqiKoar2aE8SLdPoPXdWGrxeNUG5e50MKZ2u3KS
bT/qrGTaTAFMGVCfWkwkt8GbXrU+PESd9rPbEd5lYF/NxtnZnFvVoxOcE7dqphLSfQZ8lyMSOJWe
UxMWi6G1kgQt4FKkP7hFxYJ9MeNI4xKa6ItCH3teAGuSjwnQS3KNiWbLf2oVa+BhIEgzEJFYRWqb
5x6cJkmK3nQ3slha3CgjPS9CedNPKOnX3u35vXnXA4tjI0t84CDEKONfcoDKzqEv/SehT68sGQEg
8JPCKxUfNCQgx976jy561vIlChKybjOkzGB0jaerpDPHohJ5NHHmm6JI3+YODbu0/Mdu+Kxm3j6T
1mEV08TiAOUgdMJ3En3F4bNXIkehmBrpzjiyO28BKVIr1i4aaHOwF0hZncpCQy38MIxEs3ihlY0I
gng4VlW3Gi5dsDDeFD93YZSZLeVzQM9jELFqqTFOCj+MgDOqtt8QOiMqyXqUnHrawh+skPUbP3YY
PC+WRkikxwWN6MqwiSk9TsnsfqQnPMUZB97NUN7mI6Xud61lkPZy1t3GEiavToYLA8ZOj7eOPVqC
k1l+ak4SGINqG2Vi0smPL2KTxd3N2wmYY3zep17qwp2VoHPVOQmoguUOb5JPb9WFmDEePSHu52J2
Uoui5RW5V8T8kc/GUCMCXmx3yqeOy3hvKm7ofzAjhgiXrVddMsT/9Vcmrba+Fa9sJfP8YknsO+Cv
fg90kqw3Eqt5nSRAVD/ttjSbhYw/aSFEifHmtoJ9g538pauyPgL8et45k7lRnZNEru4kXx3lhlqi
Zr1EmLt9gems3X1yubJBnN9msmtPWuXu9u7cUmDNCc7gLFZ+YASju1O0cP1UGxz9HYYCiCjoTHDp
Ajn4PjH0s/0EQxEVvEKsCYqknRL0mkwp6zDY5+hQY2umSeXpreTs3JCGQ/UzQz/leBcgUKRj7WJs
o6Pfr61EchhYJXyPnJa3hgLzjVln8hVuVmdFHBqhn6xcDUOzAHz5WWZ91obFX8UuWzARJFtHxHu7
zP3T64K1YIVcZPREzkuUqTq3B7Q3HE0H2BvgyAf6EhWYbC4dQxtb2LoCnVGGyUp3DdnkkGb/P+Yy
wru1Qr0zDo4GpBq35HEA6yOI+7IYNZU1PTandLgPLxUa/iaqgPQaPkfge/Uv66mMFRp9+OQlzauS
XmT9XQNws2GM6ukaXZVz0/S7uja97DmS7J0q+jxFcMMDYVjy82/AmPwxNAyHNyrYivbcu9Cs+F7P
fjKKKyUEWlp89hhHRL5zv/abQ3d1zhvvqmq8aosQKpmrWGR5OCwB3yYeOeDdyF8NimOWZmC28Zno
6R5/P7tiR+9awxX8u9TMx1OnkdXnpe45eKKjANqHuAttePyJfE3UUaUP2cK3W/UDu1pT5uu6PJai
3WgU6aBqXOTu9l7oOFdR+knVLmy4nKzMk6JS1bK3mGokdMSHDUGSYlXytZ9U20GPStjUZtYnMFfs
AA8VYG1qoD1MX5gLmTuBNiTvaHrpgORsiLcq4jTrpCB9RnaWoT4RwKunnvqGOZZVWdLxh1Slx6DS
VlEB2m/mjPFtUxsgMzOrr5iGAHbDquIipwlKhvdSIbZwp6mPcr672U6TQUpa/BKEB2/9TgpQkqxY
clJ05nOg9u7T6m/cF2uafi0ecn4ia/GMSy26J++VuFRyh0Qaz9eV0LNe/lLr/iFX9LcVYNsJznPQ
KjcJfUFxc4c5ZAsS+DCLyKr4+d/QCrybYkF2RTAUEHUEAPOwhvUqV/SdAk9616JZyhAAB7E5sXgZ
+2IqdHPPMzzIUwF/fo/wMCvLev70DrMzqXKhDXZtkR6QI03s8wuwfdURJn3VlPJeJbJ8sjVbapit
I02xtAUU31JtPNpi8nVWg4cTWl83qd+9URJkYpPFGa2BO8I46fCkwktzIQFTaptzojtMnbu02FNf
EqfyPVdNRMK4AT5gyG6YofstftIMTIiddCJJD+M3ow7/8Alq0PZOd8IlVNjUhPeHqF49Di3xfX+f
54h6iNa5MfN13wDQh+ATsxVaEjwQKKB7puxw7pQY3Np51p5utPa/8VO6xKdzhtgfNA5mPeJdv45f
gsfHqzAB0VXVaPgl0wNGfTSLEHJPnQOuBo5ecl7uIE+jVJZfJQZL52jRTHGl10NhmOoKUqU0cgr+
5LITQIbs0jRCgiT+UFzubBhVBv/3KQXt3NlCjjl6VbqsrX6bxvJyuKF5cRrWHAEeIYXUHsiSPE/Y
BCGYD/hbKl9eEmxBHi7gG+iRQkuUUtdmQFYUnqiEU8YJxKIxU1QE/WiSxf48V5TqWupzGBDgWTIf
mQC1PuW5mYGEbgfFy1wbS3uSvN7fbi94EhWY7H6bAY79MczfIcA8XKp/+pDNumY5lmqqvazKGGvJ
x3BN8NOBb+xHL4IkMExXr2HvPA0vWhERR/gQOFZi8AsGBY/+d1yOSp3fU/89eJwufJUPa6BJJIPL
doktpXx4iD6DbQjQ7pDmMOXtIqGHINJZtHsaSo2MY0BoD6lwNmVDZHKnXmHsAY3qrOkLuynVzOtx
ZQ/YK+rvRznwKTHIhM/MDo9Dqxmir8pBTU0gknRzvl4rr4MiCdLQHLv8THTCe+Gmy/45z9xkv1Gm
jkVUEvWlHA4lMRHZj8AAD4Y7r6rFBNkLmaJmMwal8BfD214Xkp2y688GjYiUw1zcW5k1Dv+I+2HO
Psigrx+UscI5qxwFej8ICQNzJVEm4fg2Iz2+7nbuM13YF15EIZGpaGVqT0dhRg/Q4Y0og3DVffDz
iYEunKXY+6zzGUqTLKcMQqzEobRuZbsyG+Miw9etR7ZkRvg3rtsqSFtJ9ITO6c6sdjoMoetsbiNj
0dMB98WU/ZdgUO8grt7xNW2BNekx2chjTCFiVfmzvaqnn+y8ukR0Htz5Nsk+OA1j1DrQ/pwtBSO6
+SQsvMtaX5okZu9rXggU4Rx+hgCAP8t0876zVUkLUmTD4nj2jif0+Il8TxqIw9h+ipwTpKazVG9Q
HyEG3jRFg8yxKMqsAW7Bg3pOB1vvrSdCuq1G8tgOqnJp5p2gb7Awh+0jYkvjEm4uovPeUDMWMwnB
KZMrOIiLsPX0BV0oBp79LPeoM7vp6Sx7pOgLM6rq1bUFHfWs0LV5RVFmvfg/636OWSpyIpac5z9S
e5YvE20wH+gccRTI5inaLqEhoS8XUSc+TSZ2RPM0A9RSivmm5J8xguTBJjd7SpGMhHS8utSVSXro
C684b6Dhv1xrKTFvErosVUAcFdoySZZFhF4RGr/wXN2zbRVjP8jJA2Us0cfc4XagnHMZON3f2cyX
0LMZtKcqrWUH9FX4hht+XpRpnxh0kPeRorGZ7/EipXWRESb3oRy5TB7mWs+uJ3CBG9mqHUnIRhKy
iEZU8/8hugxyUhsFlp2DrjH8foD4ye5Oa+B+cESCYuReA/GXCu0akmoN2Nk4BZpJXNa7M3s5D2S9
gKC1ETtXPcE4SDAv5oQJiJ1cBSDStlAh7aqFjcbkOil+HGTyQC4dzlAIyEqNQpCUr+JgF+ESjZ93
/GD0gaj71fj5KkY5de1uwuC3/AdcsqUzowAmHy9S1YL14EK8UiDyBBRLM4cyS+RVA8uBKHQv3Nfp
rl8RIbxEpFvkQumplhdib5DOQJ/f3GndLs4LYbkWEZOqLCa/AcFi/F5MnzBlBG0Lg8a0FhKiJ7Dd
E/k119VNiQkfq9DVUum9Kk8OfcqTslWIbx8cGOOBCHLLLi1zj+nHyIUvwcWZrS2ghQlo5iVa7VZ8
3txEyh7ZLBcP4fGvDLEaDnNZqGIiAiIgbeI4YcuF/+b+Zxmibx1D+WajFi6hbtX+yWEUM+1VYgCF
AiJIrvlHDilK7W6FYIc0geKOMZdMXnmkajHelcgHfcVAlZagpcFRSWWZV2z6msQ8ZWsl8RJSdcyE
aOAhPvCsD4aM1Y7jDfday8HWMawH7ahtpFjDaBwsvFTyDE38NxvWvWXLAV3Hzi4AjOavnOErZkIG
rTp99lsZhmDDR5YDZgUNTwy27X9tqzZT7x77lytbsGznD4PbpjZr1p/fGV0Kldm3iaCR8kd8fxuX
LxgoQp2sAbML9REOnsYdXGWH/D9UC4cw9Yx1YfKhoH7KzYfzEjby3jPXfWW/DkRROrBfkbXouIv7
Qb35B2TXKsBp7XelgsxlbqlDR0QANmdxJ0JEChpXA/BPRWb+0fZlB1ngb0Q2gYDVdESB8T5rSPnu
yq9N0BOcxMiPnlsiveU0WSan9hQBRxsMG5hwFCjgmDVYWENn6Kn3V5GoovgFIfDbAuT3s4ArF0PY
fogWDU3C2QM3IGxmzj8I6pWf8ZpFcDJnjQsq/X0mlXX3xDfVNqIP5l+I93cYY6KQtWSRJ+htuEj7
qOK0aUpAO2RHucXaX0NvUM3qA1OW+oTbaGggsKz0zf7m+6Zye2hLpsH7oIiWURNwy4tpmxIBfVqE
w4FxVkccjlNDTnwRD/et0UfqyRRakTonNT4Z4RPCv5BjKigZr5Mnt2Ux5QYW+mXQ76mq7d3q3vdT
+bJU0gCvgTHZaTW8P9WQ5ulD1eCTQa3ZFw9yrGLoDkfgBhFwVVX6Ou60Yd1uTOQbzFreTlBmgGgt
aYmhNGvYchxeoSrYqb9YdAfuExcY1Tql1X6nCnjHDtcoc1XWJIvVS6ku+VriCU4OBg0DZheHQ8Mw
KLNewXixo3qtOBTwuq9P720g7Wkw7SdRlvuATvSQYxiOkklxq4kAAO8pfit/55eyXBeEiz/I1INb
0QtUuMByxx1jtL5YY3+v3Hb/+qrpLwCS6PLkiJJ4tuYUZ5/UxjqBtfr1Dc4sPYRwEP179SUd1paB
z+Kp7WSaD0lze1fOFqR5uhJsd4kR2LlPaS1rf69rz8HSuyfg6J6ofYSr0YIfH3d66d2CuxMZQtD9
8x4mbXLE0jpHsRdSkRYKSnthHAbnb54Wdg90H9Hau+m/CTifpy9CYSkAtkhdGEwAslR6vV554Qjo
pL/zciQHbqTU9a3/qfav035z3nPcV8+dSr/uqIr9NeZg3dh8Cst21sDkOrvVTVK4reJ566KPgB5J
MLSNOzp8fR1Fi0pyQxILi0D6HMR5iRw2fYFpH3RuwEaCZ7h2KBe/JupD5UCZb9QFddrDpGWVyqUh
xqhEsGgsPjlY6eMujnURrk25JJ6MjD9DmbaOvyzNnMLePvXMqnJZ6Nyl9PFv/glzEU2VvJ50uxqK
+GCCcpkBxnh0eeHzcKXD+/hG0a3K4PL9puYbkq7DCmG0cEx3Q1Ctlx83BldDGL7hIB/EOo25ikJL
bnROJCL97vJ7ksn0sp51JkF/o/cRZ5Enqxelmj0tDFqjsW6k/1rV0hEmK22EL00ea5vekPlVaRjw
lPm2GzWxSIfUjNuCc/BMuniwFy8+bmR7jAsIHfP7FYWDTgsXIkZ5ae/oEUPIZtAT+ewkCZK5Khe8
Lk2DT3YTUbXaqT3FA5V0tKk3gDxUuWBY/PpU3WwEjsTMv17t2yPndptaV+Qa1ag9mP+RjIQgsM+h
lkCCazVMck7K0KguVYaZuxUA+DLaO432KlaJBqF83OU/vhG6JfpBXiFO/UIJWKOfiQtx/kuJJicu
QdfjGp4eOcU7Re9HZTpHmGIa0Tf4LDCwVSALE1vAv5sE3NI4HiYIdwKbeYOf8qJT9aFoPtJ/gX6C
PNmyLEXby7OUZnLAFKrIii92hI7h/zl+nzUobCz3V+eDBMD/f0fv2skSPj+A+TihnWbeNxGCB+iU
cb0MOdrSHMQiQb7A/4X23RkAYK6ReN+DNoLmN2n4PXtynr8102I1uUPkOFMuyskCJggD0VCHqKAd
hoJAKhLSaIzhKncT1yPU2qjLS7Xr1MjVXRsZ0MxPHff3WpqWDIOlosog4I86fNmbyAWZBgJ5FOsl
K30dcM9s5pLLwuXKHJuDbyIST68AQ1Hm4sz4ktHZbxJdnCVRpxoDU5R813MWKRuSzjEpfVyMRvRk
7zRJkP2bZ/WmnEt2o3n+p8q1ARDV4doDKe3tVDRxVVxUVHueQnGz6waAmBt7UTcGAj1g2IFvS/0z
QaQ36VL2VLkGVJwkDxwaSIWOeX3QdlSgUMRvpcDSMpQgTG/vhD7E6ir1vbGB3EhcnbqR2L2di03y
UFqWtaOPc2eNQTx/J9jylFK+hGrtti7AFn3Ut1P0Ok+7meI/VHI0LbBFSfiM2rSZ76Oeh+hj11pa
vlRWNzfqoYQ2AxOlDN0u2yWVjK2esNrDDqgBm1NP5KqqBaGGz88PSlKtJhDJJ8BCK1yrwZ+RmUxi
sFxJ94KTMGo6MUsG3gl7jJgPl3z0FfGsYINF/pPFPw5Et7BZlbzDFxEusgbcYHGDAVipC5x7DLnD
puXLuDYUki3aQ76epl8YYGMtJoYlySojFWmD58TtvxjfIj5PvQLBo6cbhS6xt+NU6Ctc1pCjvxZ3
mv1ajj7IpzvPhaVV4WetyXWx+Ej8qOqhmx70B4H7ruVJhBsCLA/R0t6unDxxqNSzkU01QJcWK07T
+Lu5qtMHdUStHdBZEOZvO9MJFyfsKxYyIVQ6c7/UXd6j7+h9JE5BLSuKQt9yr9O2RcViUPyR++C0
N7GhqRge85dNr9XX0WE1BR0zeAhrLDxo+Xlk0Tcb6+Lzoh+MhQ5CjRHJVTTvBvnP6uf860ul3O/k
jw8HGOfsTpH4mXWFj/8f4fXTDF4e1yuJTzm/FZq44peE4JynXkrclWtagvYCyaOWxjEduSau6GvR
5IP5GdaQ+2gTce69n3PbyzVvN2ciMUyhji1xBxrmBM0zCMQmP6sQ7hlk+b86MmjnLutOYHiqXj/e
oRu2oyVbqWmEtxjVt26bldrDYnYnzRWgzJ2NW04bPNIIeAA0CRIIBNI2p35qG9cnTTAeXT2AqClV
d5XBNVjaWSc4nETZPcKkL3XUMJn8ur+ddYrSXpPWYWdL5U8QqjEK/s/mPdZ+3WVZ9Qkx0lcYtD0m
dcpp09/6rUnZ2mAEAZYqQnTcuXOQNrYQDcVbaHyQL70LrsF8hSpU5AAcJP/rL8La687JVkxTmf7Z
zpPzjxAtGMi73d4Tz6ra3uViOdaVhhfRhrGq0OnqTW1ClUxF31OAEbLV0vn1jYWdLCA+H6+ijDUr
HQVEvDxhihDsbrj/yVi+mBvAzar1gXZAGwnVSm82yv1Q6nhJWbDsQFSNnVTA13Rk4lM9O0d8AaBc
J3n+wh6lYKXZCq6zpRj3bAKA9yjR4osWp/5EKW9UqIJbgSUpFN5SQjPrwpH5ZshZp87egtkGoEfY
73SMJ7dIXg45OipcSr9e/VnTzlZVKM7vsZDj6CgiHi+Ww0IgDKhnuPlvRsNodJneLhO1QBFjiH/h
9+f3a4w02X32s01mShcuEMmj2vuEyUIApD51hoYgqaP0VO8pnIyWdnRHW57Kp4E7/Ob329wDnubC
jui+5wSi6wZi70sPkY+7tRsRYcK2QJ2c0rO9T7mvCqr0lS6KcHw5VikceDFBAmJdwf+CiNeSZgYy
GC07AZ1PLal7T9ZgQUmEy6S5iY+p7761egdiUBSxHCYDh0DshuSKCaOYj2U6YG7D9hLjjJCaKtK3
TvjaafNSQPY9DJF8nLXs6V58KBZnRKM8166bu/5xpVLhyNPaLywptnPCPoq86E/xITPnYiI08U11
uOpjyme6VDg4XscB9OmJqQu9FHU3WO7Q5qzy+UFRj/kMVR5YeuakhlXv/9YznhJJdci3p9fIaFyJ
W+sbCnAhWWfxfR3bxmFwO/8vEVdFrq9GSA4VjYyCPkorMYh3KZPGoMsLcJdJGiGXLJJL29BHNX3Z
ePfi0AslhgtYuQqyLb1PEUuqC3Xct/WBASFLjtoNX+S/T2ttEosLa5+QJdYfc65+zf0pLyDetESl
z3vhlfg3B7aatrcccMKRfWr0aRzbSnWIrwtCQW3dN2qNP5d4zr5PVjgrx8A5CxI/GNu8pIXVF+DI
KKUXGZNB7kYvDsfd6AQPMdJJdMTPci8S+1nLAXMz/6qzHcQyBU3GSQ9kwmAAIAGx5JvTOogrVrWP
8ML4GXR8cH3DOdrraeg4t8BH06PyCY00wyd/pyO/ok2GBp9bJGCnQNM0ykdtGToC0kbyYoHAccOR
2ElsT2H3fflMxWgoVrPkNIaJ2MOF5t5SSveZXSIBd55ZtBCGuYxGw77xC5OS5pCA02TjQnTP/FqY
YjgleX0nhV+IQHPKT9RAsw0iVlpEpAliW5y2V8+ND2jlOwKUbo1vj3pt+p2pumHx2t+UT8KB879H
WxKV2kj3y2qd24cuw50OjamvVTDcx6F+F59IjEIHuX5wrb9tyjCHqMAnbrCWug4M88CL22zvSzLP
HwbE+7RKaUps8r5LwMS/LlYI8CIec2Tb7me/9JX/T9R2iGiZCwBUP8ygmTRASk/pEBoiKsZP3xlM
I13lTKLdtc/U/aIhYUphPz+8hggP0GFnmWjKBAI+2VPJkRrXsvT+xDa2dUxjLFiMc3hA7hq3uJ17
SQqxCWECWuE8uep3gk6usuHC/Gcxut5AMf+Dko8MzrkdNQ0JfgifzBlyhAR4/kplwjnC5beriaqx
YdX8CjS6QZ4chzfivC5QOUoagW8O2VO3XwZ6fkqiexJf1gTKiWvX9pk+bg07XxKpJ8IpUTWCYFOq
noj+nka94o23CDrXbiRuSXPgy/xiZuTkSdGcZj2kBkZHeC+SZ4rjTCZWDerNBVT2XA+2ZJbTEi06
GIGfAeum+rxOKzkRpia7eDWrRjUfMEIZX/nmHrb3OLTm7npOWdfKIioJMhgGHQXfu29p8CmuUXDL
quauvVT2pscoxcm9xRHJqyGKPpsdaRavoo+FWnVx1iWiBPhybRmVuMqsQzBhVFYJbuHzycy8Xvnb
UO1IqxhXR6atjvzP3Qq+SdBjbGtxuRQCRGhUzGv1MsVJsxWkzgmP3eKbGI1AfETYWvRmLHOFj7/C
Nw9wk/uqPD9WRPE7dFO+MEMAESaPXr61U9zPYyTxx4TKwbvBt+zj18fx3LJdXSlw8rHdOWn9Nabb
3D5TrqPJ087TtjcBaIT/l2vl7J8jT0gksZgL8hQH52GCsj+1TozAspKl7AV5X93UovvlZo2MvNcX
01Gh5OQqqFRRdhZujnGwkpZM01b8vUYJZ3xUwuB28D41PS1mY6qETnaoc70ujUUzgE4nGCA8OBK9
XQKKjmVwnW86xMWUglv46o1Zv4pjNfD7lbp1kbPxLW4X8ObcEWY2V1AoW9/eolFXoTj6LKAskcLY
rNVS4KYiymy0tUg9+LyA5bzb690cThRUKLTUeOWkeJVAsWdfVZ6tVGIRhEP2xgJ0xeu9d7t4D71k
dT2cEjdKJVQc7q8JCtFG4jtoSKBvhJlusybW/6s8UvE77xih5+YINb2Gk7elq7yu3rxREb5yiKyr
ZLGP//okaH9DQMRhDXh2GRG0oJ4X4X3lqjJEbMR7MDwoDKVHEnC1J4bpFZjtc9t9OfB825MPuVZw
Rp9OlYZOrlDj884Vu+kVkjWVTHYTgNe7vEzuWqy4Vvf0nczxY0OFDrdhmF6IMcEyEW8i9gQ7WTwc
k4FjV7K/xcXhxr79kmj63ZVErMJ560TvLZTsh/rCjjWUlwWzhtRR8Mu4ZevXCj3LpG+mvYvpl9fC
9yWKGaZR1lH+E43eNOQ8ZoCkg7J3uZbl88+zidrt9Hew+f9dzr4Gn52H2aOaxuiyYkAGn6Ui0Zud
OQjMy2YDWU3+CB0Xq3sSzFWurTLbb2BYfryZuKBi9UXmx0T2ISRuui6IHIbwEFjzRN1gjLqHDgok
aOlPpmSkWQF8U4Vmoel8U6cuckg749N5BethKcAmWEysW+XDKiRM4TsrvAd3vt/PySUaLgoe2RZ7
eo8ofP9CiM+yu3UE8Q4mdrtnbS1ES50OZRUFONDYUOQSEvYgFnO3HfGdwxFnAgSgcE3x/SwIUuKI
9yxGwfXepemiQcsXeU/V3MEv3OuD3TgTojHMnRhZInKyiGk4OET5p7w+Qt2Mu3/6kFJMR6idTFkV
YWlnV/Oski3P3xCIfm/fN/34VZBa2UaX5djVPM/oTDGvCMzFc9iQzICcYKOSjbeMpYl34x//DOTm
PiXGjr7MNWF4xJkSao7Qtbwnn64oiBHfIRMbehmRDshUmzorMZ7AkVw2DsfrY5VXHeZqeBLB3FHx
wvd9nRMTiGD2EXTJEOVQGTbvHOBXtR45YtjRwMX0TGbRa4yn1PVYSKPSEAY8qj7OJbSfz4zvG7LJ
7fE/0WiXZAzgFm9S3SWMYFp9K9kARfvh2haWfneFY/xk4/jWQEPl05SR0xqp4UZErmdv5ZdZ+YEJ
H7e5zauSm+fUqm0jnziEfpEU0DElhC3PqeHn80vxJiHugTjfncQ8jLTuOUCjcfL/Zfa/JcqTYbE2
1OJRvlVOhR3BvlE4GhEgg3dCIUm6RsaSHnFWUnDQArgQrNEH56IECYmxxHECn5+Xo9yoibmliKGo
+XTLq+hj1KchUPgJirYQFW1SXs43wb6Z8G5YmmuuHzOh5EU+XVMpt8zZQzfdwdmS7DuYOT9FJhD8
NrezNGrkY2oY5LVpTzpddt5g9TOaC4sN3urWVdYvvveBGlWkvsucp60yf28p8VCufk3qi4ThVQiF
U3W2Ucqq/hoExYJuXFNC9ezHEnb4Di30+5C9yFcZXvtkMJ94BcyAbHoHN+kDH5XajPkzlN8uiwu/
Eg53YD2Pb36g5wjB5EJK+If/azhJxjap3jKFeGqQVlbX/1+a0vsRCyTlYknzl9PFOdGnywY8XrEb
NPPfEudJLjWjjjVwMvv7WPrRCJQaXAMA5gZfuLuYqx30VFhZzcgpaNhiMnh1M15ApOZ/Y7iN/ZPU
v0wDHwRWlXpOmIYa4jlIdPjvSpxxzs9FE8xx0dOa/9nS2E9rcMYQPdkT3aoeQAIBQ+UsDYOhWfu2
1kAtaBXGJ1pVqSKe1fk1sfWaPZcWWE+sQNooAGgIELRQkQaINsnXrYdJES6OeBK93c5OLhr39+Fd
nlsegaffD+bN5OhgV5kpRlJvGjg+y4DPgQGSI0ygWFDle4wDioPrnbetS955eQDVY7Ud7EVxoTaB
ZGl2x9Jp/c5a+odjSr7T1b0hsZ0T6aFfR9ZucdylaPmWhBeiN5+1MkZkIbJ3QHqk6JskGWedGEvW
EdN7Kc9Aj3vQ17uZ9N2dNWHDTK6cKCw946Q14ZaIn2+0wdomD0257T0c3ofKHP9e+eRzhevFiwjE
GRfir0ytC1fS9qAV6V9s9ksr+hYh2pAzfn7oNg+qqJIeQmgTHoiprmzJpLysa09lQ5uRFHbqbest
atE0zFPbdq2iP/7G7i1LbMJZk6lxBm8+cGA+QdSM/h31Nd+lZ/F45BeAVz8FyywNjdyrIWmuZPAG
dSRhgUsbaYDN6G0zfV4o12GtMbdD5fGugjiBMqg6Yp/ZJP+yJ6O0Q3TCDQ6WbTMJzfPrxeDYmNPu
3T5BvnZd7+z41k1xVmVq4e2upfmRANk5+xb7lrJblwxgKZGE3SvyKrtW2m7ief+/gIWv98gfblhm
ARpkWGh36ri4YKn9Lce5joUo2nhJf4tRwtaA42iEIDbIf3nm8f2utXzc/oV7OsoPODGk/JoiOyFr
/o6P/sTY/lJEV3euYBkDj4TdFKpV4dvL4RLTsdVruH16xqL4olKYPOvCC9C0CrDsaDYy4Nk45hix
VzTayzFOv19OCzSAVGR690ze+5WdtokaYQJV4hKAOENIMxPvktOJW1LzG/H6CnPo40+aOAtE5L9V
n36uCrspzRFzjcYV0trNpZO8AFWwsxDugempOj0c48zIUQlIeEWVrsjOqRVMRqAiK1k8+YmhxtFe
i10pcBiWI6UaKLYMvY984QAo/N0HH4Qvz+PNMDOcLeyuBPgtrUeTC9fbYWKF8eVcxQSIAF8r3LYE
YiGce4PhWdvM4BpNP6qxYvn+Np6ny4x0tFViZLEutldqR4MssSEvihlaU+9slKXr5OK/oEIm7jYo
92GhQMUeibK3vsdhkhR+dy89lqDgd/tDL0uSwJTjbo6FICoP3/G9pGt34wvg1GWp0QGohiEP6YtR
7leb6xB3Z8FWfE2mYh+MOhnxHMAJuYH5M04WZt7ofwXaVvmA9xy8w2svc2hCTk4gLQf99A29vD18
1i9pnfEHraE/WdsBlr4teuSN2q2IkWleEyN6JgMGj21mFXhEZRFI8ZbkGvmnI1M9u5PC6CcuEaFB
bH7gH9CJM05PJAu89eEQ3JC1Orpzp04/1DqhdzZuXLUpYVvXZY7+nadN7NgGQQP+Ws4pl+GlnKxK
Q0QSPbFPpRc6SUO7IXWld4Hc/yCd2b7P3z6D51vboWP3R6XvCSBHKP7IPLfPuhlT3NzVOCrJjDHH
pL1SdsvSC1LY7LAXuBzoZzIWdjYRqBYhDnyP0GF2KSYjId3u4/bjlzVIOJR1imLoKUpLFLgJltC9
0tgy1lbZsJ3u7Wz92HCoIrC3EDFbs1oJjdmzPINawEJSPy2RppJi6D+29Ty/v/kYINCGuWDSuLI8
yy+cG87dSEJ/NUxUa5J7lfsRCjLPwFML6/XuONjEf2jWHtnH1rXvOQRwuIM7AFIlD3scdvsNwuRt
j5V3JXoXOhnHA77Infj/cjXRtPWAwHiGkvhwxgyU/klTCBD4LAziyEmc+4IHe4Op4aaIVI4ob9t4
E2NHq65/hyJEi9zSw9YtTf5sTp1azTZSIc0qbSRM0bWfLrTIRFztKHHs+QCA8yHRWh6N5N33wLYw
sLMziXb0zS8fZnDKy4GmcbNfnb1KnhXAOAxQsYG1bcFAfZrF09DdaL7peu9Xw8RboeUqis37D/8I
exm0DuX54kq8efkdQoKEwVyT4+yCjqDtstiNY66MSGhYvu20DpbwvXjTmNjbzki/5t+VWHn4bmUJ
jnHrc7yH0JetXnnOXDIwAzkpEG4OkVYuZplD4u5g7I9kNC8l+KauBtsFP1jO8TUfPfZXMj5IS1Hk
fpCwryfq3XVz928Voy5lDzVZ3v6o2l1bQT2U+GtaZK+4MgzZDZzP0C8KWTALUGycnGt/Qvouk9yT
nUBD90SL1VBVDKrmdmC3e6VpHotnZYweo9GbwWGeScLWH8y8PkuP07d7uVz1ZHTCgfq5notPMBkR
g0vwtGbSW82wn2DptR2JcNPZldnRu3fLbmwKLw1hydqJUU3dg53alh0D5PWASWuB5fxzeBbkA51U
gIZMbTf27tDW6XZSM93DwkgRuw5v2BcdtGNG36URG78YHSAK+E73Fb1k1/iP7VwX6J08pEtCVDnw
ZgDdGnJ5C7sX883sv+dxj/dt8n1FbxE+8qQrAqincmTG+n4lcO5VTiN5iN4Oq2oQCjqD/OQfXR4O
QxGljj6yubnubmSlI2K/aFWsvyWp+sRQM6uZbDaYjC+AbUJ3tfBUGtI6Oza3u40icd9XcbdEoAh8
9YEvmXw7V+NU3RxO1uiH8vJL7Piwm1MLLLltFbhs9VDE81TJWw9zeZZ06BrpqBLSrLU0BzSPetDe
w48Deg5BFUIv0lKv/Z6AmKbBd2vLHze9vfMAZ6M+dJ7RTNrw/XLVSvnZQPwguKuxZX/uGoh4prpd
67Ypn7VgmUWZ6Lzpd+VbE3hPCptmzRU/y9Qm3pg29fK/BOAFc2dF8DxizHBeiazMVcGLMsr368ko
9b+5qXxQRIVm00x6bnf8bRG5PumX47lVFA1mdPf0wZWVDtEQEcaTOLyobukxgjv+BhOUQ/FNU7mp
rWZ6RekUKnttTzD7ZG5EBYT1jtxUCIZrL93i22xwtTUX10f/DMJkIpECHl38CP5pxHA8zASSBgpW
8WJ0SxxINNfKHTsyfB75bg8Yt7an8Cub2mFBI2Y+65aXV6oS7PjnekGqwcsHQoMzCftkZzGpYAtS
8XeGPASKeiOiIyqt6U+ZXsvYPFNhGsiYEceOHrJIYsBBxX1rHoLyw98WE166V9Ll4CwL649P1co1
TTnSqDlzJKGb0klAjqKg8MpjLd44/utPy+vspsxjALA8WhlI3sBwc53xA+Cy/VapxKPVB31O1T8o
QDs/tIw+/yKfFe16aCOOiM724RXKTPhk/biQlzbyf+LU/MZwHVDc+cq7jvIrGh1VKWi2yUr/OYOT
iP1BI33KOrXBtue3X7+flwOy9uG5BZUT8I6v61G2Zy5gxptHX5KDtyiQ3bY+mwSMXyKnzF2aoYLH
nuacHl7PHVNKlTfzgmE6/+/MCAdtEEcF/IZoBEqlgeNqItbhgf96xDYnwiGERR+L9770wKRShabX
7aCLNkHG4KbxfOMoZAVd6S+JpnuqW6Jm1jdD/UsjtBNAALGThMmx/j946PZ75sXRkr5zr5Rxs5LP
PRvhyziUQWUCaa8qcICoe7VIqHCjasEcUjwodlIbpZZWEf0/IE88mENz05KAOC8JR5pysEjfe0xN
CujRKd+2Nr7DzKCVMEXMODiMBSqWbiemN3vM5XchjKcRIzyp7Ifuqpu+Nm3ce5y+PojN07XDIM1D
/HkvnPmJFKTtSpXOPv0PybPmOuvTC3eFuXlclPNrvYWQ5ngI0tRq8pnzRmR6NsyjxBGC5wxeNwSm
THIue3vqAUtUb8GiIqJ5MlK9JIGgaAUpwWtxVFnROx3fgYxA4UIX6GuuoR+DWV/XOrlILqTK4B4x
AoZ2osUrqBGl4tZXx0lqBHDMvVV6pSer4wVXyv/U3yOp6D1AdYkiOywfCmDvxT9wYMThr48eQYlS
2nBaDF+E4qy5IGX6ODPm/e/W7KxeoTW/7sAFOYmPUaYoNF207hiUmf+yBws7LCH6e7TVRyFp8QGP
kxGAo1600zdaR0NNMfrxH7IryQOqvbNTTW2ZnsZSjUeVC84WDAQZ2GHwjXhvXrNwi9wmXlZrxZyk
tyAAyFc9lYGthSxug/ltHCYLXrTbHbv+cIS1TXQj1ySp8Fd7DkChx/a40hdg47H9UnDP9rtqxEM1
/WjvpIcjD3JYoerf7WpEVFgJeXYRxZZ0cqqiREk+3nPL4Km+Fw5VK2VM5j19vqwQcqlM7/D3Dqzk
ljBEL7pvVgJlxtFVvImhw9NQqncjfjfjqMbUwr4Myp1U0i0eCI4E4mWgPD7zkXk3XxwUXr5pVwDh
T18g10IqCGPdwTzz2jIjnk+9v5v7EL2jozVqjJQwV20ykCcsmzDSZl2B5SLwZ8W5qhubyEYDZmYB
FiawXu2Y/mGoGuSHe4L4+YXTtSPCLtqS4x6FeRCFNOSy0GW5auKbD+j+DMYrLXd7ujJlxjpMRmfN
77dWr5j43pNq54Qbsrcs8v5MqnExE+HNvGfZrjmptPmpp10hfW/KsK0Ks81+ROxbeZXJ1BMHc/QA
0oLE4K/tmJxlVwpl1qMzlbLH2Mr4OnflVzqyrxceWnLeDXg+Pv9rcz1/aVlZbMQlc9KFEpaRaJmY
FtWMSxBy1T13DCpvJ3RPtAzZtJ1r+oCmqm7GyZjpK11jek+cuM3V+K4/P/h6u3q3xXi2zWykoPW1
C874xQEuUZ3NkcvwFpG3yvw+f07g/pVsE3h7KidWk/2IpH/iMn5syjJtHRWOmdEoN6yPNxzcEnAo
87DLCGbfp+W95q6KbGVHUr4QTAc31Acyeym/uE6cCqXcXE1zFYUfHUZSbEmUUS9h7pvE42Sht2gN
p4xknuSM1ESKb1XWOz5GNsM/oRQldotR+VhlZySyRG/93U3CrKhdJ/crtVXrX/ZTEXiPP6gk3Lu/
Skc/gks5t8XN+myp98JmAIJh3I8AqSM82x/c+ip8rvVBph9pG1Pugnyv3pSRS7+8xI5jiPXR5RA+
7NgJNUrdZMIQPZTc3T4+PiGR92oYJsJaXGJpFGE5rqv7W6wiKS3mxnw0zWFojZscImcX6nl0wL8g
P8yJKCXW+M+WMYNDoFP9rBVCQ2b2VGgZ6KI3f2XUjS4pzdf+9u1p/J1vKJEw1Z+S8Q2d4CxdnH5V
7LcT+djgZcJSj104MvvTAJICijUaX1HY4TA+UYROGNoe3TZ5o2lMotRQOklQLFldBtxdm98k7bRu
p48z1VRKMtvUuzET1MP1BTUeh8moHgRxmePNGadSv0Qxs8UtAjy1rxCsNNA1hhwFeKZeb/UJdR8h
3raycVby6tAY7PBVNaX+iFXV7D0ZsmSJSQiTaaNzKZp9Zi5/gjDl0QL0SP+IDKpJu9Uq9/IPfq30
fLNHiUhRrLU/qu9FP4h0yto+PG+bbfdlBpMBtcAWP+GcnZPEiUYeQNkxC6Pt+dIYdPNpbw9g5+Rq
nSYp0w5oxKhNlJLmVFkxVNMjXPoAypE1AppEt2BwXq4FVU7G1HHpoznwFdMTeR9r9wD3FHCV7ENZ
dPd8+AGo7Qgzy3pg+a42P0DkZsX38WdwY2NCunpZ1VE4H7BePgTlyZKYD9EGTxL4AAl2qJhj1sN7
LiFnoR6yvgekUXGTH0y4TnB5VSSUOm4LGnNSiZIHxDoLDphimeOizPa4Nir4NjwVijOejKnraCXQ
ntPB5a+n6FsUYEoM75K/GpymVvaNuDPlZsjKxt9/JCYpE6Jc2zRannsy+PcxftO9Depw6Rjon3q5
/ULGzsN3CoTv3xkddZzFG6o7Sb6jvKogAZanDbbqCTwB+urNS1QU6+KDmiIEbZZNj6O58GPQ/szn
KR9+Y7A2JqxnhAMr5q7jN0Bd4v//GM+CWCi5X/SGOob3yvMDDfTVEumeGLZlVGRmfW/8QEUJO1M8
9DYv7Rw9z/nyZ2qtvTpoF3nVgzzOn311+J3oRd0VEX5JIYv6Ir+ksxqRXYDN/urSt5+TnihQnVab
luOJaIq3jpLbkLn1ZMvXcCGGxqP88PpJdM2IGNmQYma49gR+j0rzVJLCEGfHVajpheGp1FSsHPO+
pJmHjebvKszFHmkGZ3qGH2V+l7vsvPz4hmqrBbKtL9ta733o3b5XD4/1rcOVU9H54GxkCFg4O191
j5scKPy2zwxv0VLUW2MBDfGFQgG1sJ1voaR0LLIngTCfpTy4coiKgmxy2uJxGlPQE4HF3kWBagBz
+Ttqtk7h9Yf29Zp6kJR7hKjvA3rWgb2QuSkUhFnqRcTA/OPFHmXKi3BbvZ/300JdJNzCLbeuh7G4
qxXvliWCvS34jnqyir7ZpOyLdIXAXzdDiUErmfxz5K2CSwzVRSAvFvDCsO1fXnAOviScHJMvBI9a
9NoUbpN9kSBObUeNtuqvl+zOyM/j07mwp/QOg4UZM14J694w06jWksAw1vTRKk/FehTIlWSongQ0
NFjqdIgT7FkB2hoai528/14WRNHzNW5cpNx/vujJP1A6YgV5MJboPSDXj6l3Awq1n5RVhYpbnOFL
jqkp0um2eEtgha88LNjXG7mugB8mVELS7+6jeUlF7SBhRvfsWdP8hAfebFSvT7jxdZz0pR0xZow+
DeRdOst1TfTCf0i05kA2xk2qq/c5BnojXE4T2tRUwCOavfYCAdPg1ixA8MhBaFvYJ45nZXlgy/a6
lNf8UwvrmS8lR5qAhB85XpHSb8B7z+jFx8QakLKb7hCOLXObrP8zeDuIblndyOrHXL8eKyUeAmrx
4I/05qWPsaHtRyZvqZVjQMnHqrcYEAu66i5gTSbx5dT9ZyYK342V2G++WuDsssP9b3e6iNzzq8WA
dgqgfABhSV/kTTk85wX2CvFvOXQeyFXZQ08EAT3ejPRpX2c3Grfnj6jN3kmXrt+ITNnMlwlHKG4X
adeJnNXdmi6jHSnM8v8PlK5LBIPRb/RqYGiKc/CRPBcAER655L7CxYlCj/VVXAA20vi2Rq640ypP
PEr/Ffl57O0prL2PCVm/3G5LGdPI5YnP1fANKxsbLZxd6tRlOTs4z/a11A67BuXQssId4aDHbwWy
MjNXuJvxP1BxI1ZEH5JMBwDm5GDj+0UP0ybRF6BGkPQynKGJNFFO69Ktam+MjEsljFIwUe334Ya7
qlYBx2DpN+eFFReLeUUfFSKDhie0M1G+QT/R+T/l+TakSCPT7k5oKF/2SYXGJv633Ji57IBxJ9TQ
Kc1wtc4jRMcS5jpBm4CDd7LwB7j0r8mVm9FI2gOw//T003I88rjnbgpNLTDliR+86+gJglk7MW/f
HhHDC5lo3jdCBPmrqmthU+aHvxFQ4A0V+F5bqIsg/DIPvpGMqpqlBBfQunHCSb+BQE/d/3HptbUf
z8SWyThIxFnZkoMan5mV5NOKOhWOYAmEyMbG3K7+qm3H7gtWRj9kG1U7cdi6pUKU8ghTHUKTRdCi
eZhPOQdcJQxySlvFQNwsKf9SLmLbg11ub5TtNlxxDAhZdZiINYtVxick5z8mi9FF2HmbC3NHtekK
o3NGjBFy/VEpjcbdvcpvHuYCr032oyTTg/Bx5jHW+fO1wC50hTWDBSXSXjLTdmwOTFHC4Vtztv1d
Fg/gKQPqKP3iFRdHzm04VODMqpC+ABm+Aj1EQ26OAsdRTOuSdeidScmgZDJzs6CvuGLRCFdGzpU6
oUkSvzLRLUA3KGqtIqP329V41F6OOkNrIVgyyYmPDL0sp+lzBDYEesXxTeYR7QajUQoiuxyLZaIL
7lF9DJj9iw4+q0j2JzWwRovfBmzIdienkZmf7+Q91q3tAk3JWnXwRrlz9LFjthu4I/eMN5w2k7gH
L38RwBC5oUgYqn4F+5PaQYPgx2WtMnhqERMiSOrxR/q6uO4la3cQqaCniMMP2zCdOo64RwWe91wL
mm5gM25S5wLYEosBIGFErNrrLB4iJN/paXn3dqSDWPN2DtT4vsAukKycG1L+0Sn2pxuXEtvCsapL
l5SAXyMyJZgY0ZPUnvEZE72hbRU4mwKSwXXYgeNKLqdChQ1hxaJGFfd1PblfolVJ0PKHRDE+V0T/
Y1mcoLIpYzS3+J7g/elZ+nBuK4T5HsX8JeK1syBhHA99AtL9MqgQbAX3V4sUlkQNQ6GTmvnHhLpa
DiAiu+f6I5Fhdp6LAskYYL0/dAlkME5XmDEd2v7+lzu+yVVn+qo8rhKh2MvdfwAIKElCf2L1P6US
yqDTJSy45HUGu7eFeayBFBdzAkvv5YsFtidG+4gzja/bty1vy8RfLHV/rCEWTv1ABcpFQn+voo7W
SDh/gI9gPpcr7Dtr4IREPx/Kucr4IaVnQltcPPk3mGVqhi5+a7b8JJ53gQwfhgv55g7aG5HUZEZh
+0NU084Auwk0i415VP1omPR9wlsNkIqT0Opw+XwNeeBZ/Fgx3wStcLD+kictZpvTyz61WTdQl9sK
5NwwBlPzPko964yOMZH/sPkYJGD6U1yTP74v3OfcicivDZrp0HUG/5UeSgDOceEjgxkWVK9goUmQ
ipe4jlAF9cZ9lms9NxLYuwd5HibwP+2o6+MReN/beHAaqHlxIV96pYPmHII5GQbbbzl2u4bDyxDf
O7uEE45F7P/AzZRKvF+dexwcER5mShlTDBHJMQZw1ZMt6VsKcz4Sg+N6RnwFrkxozbkpR6BxESxq
QMoXDKszCIzOYZ0x0OPjfyPby1h5hYl7fpyPBiGScEwhbUTLPxwAku9wJ3FAoNW4vAAuBaPD2smS
DDGb9G4LaHTXgLj0aTtp+rPTTmM8b1H3PofW3WTZDRR7GFR3mKoY97GvmaaWZPSVTqn0tr0h/5FW
EJiqLhzRqyb7uwxKd5Mt/Bezjxcyli2qdBc+RhC2IWGdqPF17aWIfJoU6+LLLq7niFxUjmHRixKu
zHdeRsWKh9T77yhK/jNwfHXBprb0YUlke0F8FO7/nsuo/8SJVuuV2cvO6heR2xmdWeCLAKBoN+Sl
yB4edmxpwGIJFOhxTDGXCm0cbEFnS2tpZswRN7NeYcfVG9cr5ClS+3hAT+98f8ngXcmqZBuoslYH
JUh1zdY98swFp1bS9TjuyKi6L4gRbohGAdoUIzs4GZUPoEuisHI7tSCExn2v+eDL0h+YLFag62/D
VrAPq9GcXxBYQmnXZBcQFizm8ajlEl5nKDwKnCmZMxXIv260G+QVqkziVYY2f6x7gvmNlUFa6hyh
TxXF6UBStsOOd8bOi1zEyMufMuwBx3JCRfMYi3w9w08M+7EwDB/83ex6J896nF840QvzIpBg6Z45
AuV9p1HZv2SC27ZlQ1TVuuqHQW9PBEClYe9mbg80H1UP6ko8QG0LIu9OYKCcvqHFy2zSGTf2+RBU
oGAI8TXID5j0B7Ilkya7yOio4p4uCUoRiZPcUBJgrKTbSSeTEvq37FXFWQbKOxM799JruWlZquH+
kfDJWWiBnbXZuSs8MFTVyhNpIE5eQ+bS3OfAvL08CbApF8k/q1m8ozyZGDW95Ci3o6e6RERP/CdH
oeV04cm47S33/AzqjDiUebnZ6KmuVX9QMrpQfWzqEKmiqsX+F/rjqvPWMBzIkZkEwCm1pROkI/lf
EgDIQuWzaVs7RXRltIlLycDoUrve2VqZbE/0C+mKR7a0iYlQcSZwjCCFiZpJaoiIhXj+oF3eH3zc
qW9NrzegU71kt2BoVNGTST5IR+migVsgN/aXbD2+jFzNC0uiyYIteEz9mbJO7Cb3cefUEAO8K/JM
F20GSwi0vmFV1A46Xi9pCMOKtm2wKaTU1sPZ5CKoIE9BLAsfn6Yr8MdhiNCRKoNmQaTP6bSveJKn
jTx2vLercAicPPXR8/VVzLr2yqOl7qgLirqunbCigB4drJ88jj7uAUOecKmUI0rUqpv25m+LCp1P
7iXr68EWxmtqFQA6bkX4EUw2ijnZyzUpR7mfNUaMInX7OGmhth0OorWnWgzcz0PZ+2KYs4IXXNfF
IGhWWgRyCb8x+RCRexmP78mf5ov0OPJ52ofBg87cY3VoyYYcvMGsuYvEz3yHm0w2Xi2P3n2pLBJq
K7m8AqPby4ioKMEDw1uUdUum/0ed3XzMpSUc5+U5rnGON/Hjna067Rr5SQZMYy+MvUPisnvjiEWe
cGSm1X1gUO7r50NaA0urhEyYDIMM4J0DCP00GL13ghrCyzPQxp5KBWCu3OJBMDD9Z3N62P+NBxaU
9WMkMR9nQR2IMHx/sZhwX/dX7VC00PKOzFBabnYlZ+gbALtS81Fj9Df+Ju4Pn8OEx4l+K6u2nopG
nZcrq1EPuCsM46Ib6ruN55AUS03E4X4fKMBuWTQKZZqQ9XWTNQcQbA2Z82R1gBeG0/JHzujt3zEw
hLGsPJ+IQyLCITVIt+7N3XbO8qchoUSCxHSPO4fPHXyaMKpQtAaAhMhROz17uTkI4XS11B6vFwDM
iNBP6aRLerfgdtFvk8vRk6PRnisWfhBDMax/7giR/DIEPhDIitaC5aX7S4dQsYXmw8gv3yicrhZ5
aQknrbfpmxhx91ekodTxQAuzoajqTgbPAXS8jUI7sqOm+4DMzb0rW3nAUWUjF7ca5/YfaKXnoU2V
cUvOo/IGerhZeuZnlNCa+I3+6KjTgkjE0T7OO6r1i7zH2JnuJaa+Kd7458ZyB9tL9jcSc+wOzsfu
vnfZwE8x4PLjmAGe4KpbJNB+9dNb1sGA76iyG359XQvK6sYSHsEwGKLE27Pl8FqzVwHGd1IvjzZn
vikJowepJdPR5I0XXNUW+lX3Jh2H+vbVWnkNJx9qQirjxjTONMmVw4Jh6KyuR3WVLusEttZ0ukRW
/4EX3I6WQOJvuquIGnSuyqPzIHahKAP7AZd0WdXyEKeL+tUSnXoIdw1uya34S2HhJGCxNtEVmKmo
AScCLv7YdJReC5s5d9Ndh17h2ZojJO9mBPt1iUl8N1k1xbwlwaVZEM73LHsUbLTxn2GOo8XEJQen
IUrKWgayAQsFn2kLWxtA9d4OYA4Y/QFcyWKGv59bQTu7MXE6l8nCN9d7az5X6ZAl56MqxWygJ+XA
TW9APFpRD2o5OKZh/Gp0ATT3lX83yptAdR1xVhuGarx7GYH7M6x1d91FPfchc83vpmsubA5NZ9Ap
LcBaRn5hbiGjbWvRBAr87/UBSkGrZ00zHlzvbjXOAU7XNOwqLlL/a0HKmgulMqf71gcvEbVMKzwc
ihTE1ovYNWjRtLCB9rG/oMx48cn7ImPjqrVFReDkl6OCIh9Pkas4+RAwITlkeKzULu4yEPNGFDb0
MnkDjB9ZiEN5XY8WbxG1KGZtY7vz+/NlEcrTYTgqieF9UYF3e0QrD9XaDuFs/Z5ECX7b8pB9F2NA
y+uJRCPy35X/BdmZlcGNDD2QORA1s+UDTzl918VQbyQ+1j55pzYFmtTXltVEoWOwPhfDRfUV8nIM
+0oWvTVAHHnLS5uawVh+q7YkUe/3RF1uE/teeYRiOSPxF/xJMpD11mMmJmTOlrWAK8YjfReg8T39
uYoNvQMzx3I4JEPl+msyyAIhsIep6PZD65CmYZusK7Exn6BWQf0BKbPgeFLSoEbnHhWGUFIv03yc
HLQh/kj7Zf6Qh3RSlUja8RW13YIcxCtLpKy6p5UiKcQomEQ0WYIsCwP8CqZAVimiHMUWtnsP9ylA
9cw6iPh0B7C6LUIbOkPm7IYG7rboTQbFWAczTzmb0WDfNlzNKE34KUl9jrvnjS3gIv8KXJCqAqAv
MwVFypA4iYveaLYclUvhAQph0pNIviqiBZ4MavQvfYvQ3Kn6MwmxsbJ09bNVGCNKsWETVMXrUqio
cukOg3G7yMrnzxZI4PLqLZ3OGqZ5hmTkOC2zMx+hXacnkojiZocMUQq1idJG2h+rhhhKqnRRDScQ
OJu8MaPv4T4kS7pAqEipoqlJ1+8axcgG2qGPIbOamq8Gs+bFuVo6ZPxrfdlNOeECM5DDwtIyKgT0
1QCjC7FNau3my/YqLZRqJKqlwOP7udtZn2R07g2GD2aXGYpmupkXXWjKis6bowZ1RtI3oXZiiZcx
7x49aAITWOQrkjvT4z58gmgYDkoVDtJgLOJtFjOkrr03tv22M6TMmxisUU/GO9R9Vc7pOfyTO6nw
viP02/DtoL1piJUHhTpnjfo8wlo+0Hh4h10nCsRLIHYXFVJHvlQz7tAsMjH2JRMLjXxxf5vim2Vy
h9etPcJqZbxlQuPzzX9JoNFc5z0G84U/OukIZ/T1ch5WypYSIAiCj/dpztIhxPwIq3QTDdVw6unI
UUuZXXUsMId2O6zDErrFliIsNRPFR2NNXk1YSosrfnYvaRNXsEYBCE2Vywfos63Im568dBuBUYBm
FSLSDe5c1b1WMa4yXYNliUZtlER2DZYT2Zq2fUSj30mqp76+YeMrJW1ZqN9EkeznSpXrmjqxteBd
DDasRBTR38gC+do5kndG10anSP3kJy+KNbqwjGQxVb4TNSrAse+OLrtDlh9iD1Eno5FEP32tPNz5
Iybtx0Ql/iNg2CFM8+x+PT9YJtff9MqdTw8zHcclx07BHEqh9wYHUVYCgwMP2rhKeJbjw2aEVZ6z
ioX6NZ62LzVRpahz9r2WCpu+87TOWuvzkI6JLl8yXplumrUw1BvFSrdBzVGArDgh7hvfRg3hxVJp
ltNAKBi4KhB9JtRhIKw2e2G+jQ8YVKSGD+YLFlOFnztFrEkJRLLAWIP8uc8bnxOoRdTFiU394eAa
Xnrb1xwxml5ap6K6GKgNIffipjTN21dhnFLOV/m9L7aWw7dVsjT2CUALXDawu1GLBHvpFxanlUiF
6M8NyuXP+sRPlFn15ljgJbkxjEl2nRKf/f3b/iUEntyASfDw+/bWaqv9mvG5pXeZtCYAH6jhN6ts
FQpETrX3MhJVAI7fMexLtcSbvnOICiybG+hbUI20GGPFS8t2nb+GoVQFnxU7LIks6aZnYcDjRgdQ
9YnNvNIXzU/pGzxpDe7r7WwHdRYo1aZU5iyi5sfpWEt4GE2gLgcotTXL7D6ZRqhKBwuoR+DsnXug
IUTcYU59zRmY+vMsI2OJ7pn9QonIWFnwDAcNRyh2dK7ZCiPr5RMavfAYGfoDv61/ls81W2Lvzgvb
NYMnl3gYs3l/Rlls88xdXTcQV7M7s2rWS2JDqX/uLOueXRPg9N22lPrt4RCwGUPUIG7lafupf38u
edLahEO8IY7CxEhFfPNI99J16HSwJwpBxwqn454EHrmvg6lQH+4dJakWM2khtz60k3RcvYPS0Aok
kjzMo6Ruh/qkX+/3sNUU6ptl7ZcPEfbhcn25PawRrI5vGT5wTYrI525WJmHzLx/0ZtBEdK3R0W0p
AmnJ8dUKPTA64afUuzSw1HuvZWY7Ub3DqJ+qb0EXsZihKnT3wuENuiHVNv5ODg8T/+ibf0T+Gfni
LJgRxOumvPnixSqGUUXnCIuvzH72JL+WByFOokQihylRxUDZBpNuouMt5A56VqkBaLcqOmed9zIb
fhGe/K70jd4xPrVjBS9uluNvVkCV+zOnH8X5todiFYUj0mxNBH9r5k2COzFxa1TqNpPRQQ//yrf6
atXIexIJwFIy7b0VUu6TXLYaltpUzzXT7FEk44j+N3n6NW1ff2MtKHIV2kgg6xeaDSJqxwflMI3S
lIKM5poAG7Y4+wPWJt3k0iGUz26ZV4+1knktjKhbMi9j9Bfzvjm4Lh+8NrOgjrSvjLZwACwVTpCT
6p0tgF0eTetiSPn7C993UFZVMUZK44Fnr28i6Bb65J2vEsEA0nRdvvR7IMMNfFG4+iJa08INYCQF
SYBOdeqDvZP9dt+71wym6GPHh/0/XYtXFSQkH4tkxLM3pFAZKcq0TG3DDLPJH1PkxFRLkZPkYInz
oDb3FDqeFcgtEdsyMNlKJHIeLzjbB533UxIFu3HpXYtM7Iw8i2XjWexsN1FVU45HZgHN75KqDZ3f
/0CaN53PpxKs9t+m1iSGciW/Cb7LCfZ81SreJDCMILSVhKgrLUA4MyAWcw0JnbCWFiNoRXPtkcGJ
CsTa/QIzgO9tmYCZONPSvQpG3FfFCjji9Qad1TLwCdperDYWTtkRo/YU5uPCSlpfDCekHuKKE6yX
Lu6VsM/hwwHo4S1NoUHtoGpqtcv8eB/3Z3OTe3p6zkuVQCQALt46yp28mcQuFIEi2zAJGGbXj1VM
yaZfQ8M6oitCP7s+TRIRy+zuAKCnjtTGhaCn2PaBoPw5gVL0BlBLDh6Iy7HGRT5r6LgTbbSYhwOo
OSwVoxtc5HOtmaPZ9sN+GlE/qL8RFQJvycExFEYoImxyA+Wku4qh11lvWnErieVMMUBXLQAScV7R
o85z1icA0QnrcstQh9slxXHlzlrEFKPPpdrI5P578UHH71mZFaMPUJkJkSp9HVLFHeQv561pRkxN
CEgg/reBtNC8+tzvD939yoaOFRZzj9PzYv6z8UG2AH/DF/sWAqDWWmWfF07j2tHmvCP898DHadBN
9TWDI3jg3uZXBHzp/dS5Q0POCeoFH0LN6rZaMz16/XDXqMGkZDnFk+uDn/AxtkO+AqpUqM/vE6Ou
dohr5337TfQU1WXK34sQ/6rUtO6L6HXch/oOhjbRC9MGKp2aSP64+8UiAl3c2z1Ss/eEyO8+bQCf
hN2YijyIQpBqYbhkJNNqAxGceywJ6KkN5Z7XErJ5lXlAN4d0MPgnHIIngxkuwzU2RUx88CP6/kE2
BLLaqQb2Qca473/EUtA8GlTjT3+yRjWisaBopvSYogV1PIZFN/pWoTtJk3CJpIIRQaJEtRrIySZ9
x9FrW+qoAaV2o0nSGJmmaevOsMcqn5r/uwNkpJFfgTCZbVN8j9OMWkB1zNdWfAmmWhaiaUjYDN5L
q9fe8Oy2c6igMGTOLhJkKyDVBIsyQPwWcukRtJl6BdjuNNo4WSTDtAN3BJc7T9fP7Z6b2Nbg9dqC
8lvQmZp9SBJQV8yexnXixxO12cFXJFMUkNod4Y48cn3Mqk0TIXK7FHzDgN//DQrPFrng/dAnT019
XfGSSgQhYEVjCP7RJt3buw9Gj1geUUoHnizkELWX3wuEWV+zvciKszNN3zkpYBEfOIkKOtmlcWfX
F918+N/6sc94iH4ty73X/LpsTVAcB738X8Oq9XnWEVCEUanosF5hjCOyoR8a4V9tlFyaMN9kMNpm
0t6G3EqHA39G7whSMsLcL2yqyEcke+S2+lcTLMsxzGjMaUNGqVcgtPW0D0Szz4GcP67dLJlYk5K3
oZPHwY4lGpli7evG9xaYlebmflex8PLUT4MvzgqfXaj1rzwUnjnxCg8+PKRMURH87hF/fyM+zb61
qN1d6L5aGMCaVivmBOJH5L6h2rXMI9FTVPIpi5CavsFDq+yd1SJ3GCTzOiWgSwEQ3rkqHFVnBqnF
whFP6+4/u7CvA6KwUTY1zJllgXcStaOgaNZj6bqO57nqDr2XHU5wEMTwgeJ80D49eKI8dHW0N+xJ
zRMHErCEYLJ74v0HRhgFudVsQ6sB/RElfCOefc2co4HSu6D4s/I/WYz2dcg05lQz99sj08jA6qdI
LCGPzHWsYza1ON9b00PLk124yXxAZKHjYfqAu3fMWj3awXocjZ+LYySzTfo8YYKUQKENA/65SlBt
Tyb+BXOqXan7IImx+IQXL8K+JrjwmUdxUsuqyVHUKuTa4c6ZztLhs5e2EWFwf28cakr3mbm0gnLc
pysVHBMQf7wjXRCyGfCC3x+G4kXmiQgcTPsq9W9LhVamrDG3rfEGtlCc3f4HPw/YoRC+ylOITIe8
n633cXyNXolIJydYybrjGbNx5zqPTrk7w62ps6J8R2RrbBUpeOACSRBYupw0QvEW3TDg2P0ZfFth
4jkUaPw8SUk1PlQaodHvuRyde9FzJS+U+Y6Pem72kb1MsFCXrYy6kBP1efV0LcjImo0+/3RUKn3E
VEYTndRfuiCYN+4P04mf5i3cMfjomYHUCueDzZkGc4l/FaHVXA57Jz7fgzvkIPXRYA8bz5jzM3ak
2dPZpGs9PC/LIEN19RaECzTf4ZUZOJhOZqvS5zGvuhpBsd7YXf5N6evSbj+87DIm4+/w6j773jqC
wyyQc7XMZTNzNqb76qeqfBdIM3swYwznA7j1aHrSclODqhYe+hhfOC0Q+/vuhSfSEmKZYVpnEyJt
tMbTmXPnt03kI7G7OlNVqyRGVe1bM2xQO25CTxsQ3dgm4UYDcmLl2E6HzXLu6+7J3+CtFLEMY0yE
M3logDtuTN1jfUN8y3Kalsc7RIPOOtRYxFk22fqKLWeQB+2DMtZaPOiQWg3FpphxE96etL9Yqb/d
BSSkFN2VwlJO8G8T8XS4vJZqzbOyzAkvANla6EesyFS8vv39ZcmfXxBEtA3W1AX3cpGe9YkuPUHc
0M4K4Fsn6mMntCLADwxwvkXOB1KeFFlVDD+PrYrcC0ee99B0xaf3S89tt5shzPSCSY/OWAohT1LE
t0dt2V1NY9lNXJRyIMVlPKBs6eGz4pVQE7DYc6orZGKok5D3/cde0YJnRHHVypfoR7Nnwfn1yikp
VBnBjJb/E8Sa2TYGqsOG1Q7rlMF4J0ubpiyGIaBn+CF+aUEXC4SCqj9Zb4rBao0USDunSxAuJOxx
1B/LuD58sqTSvUTvxBVa0nqR40dq8HLcYL8gQqs0OQY+Jnm5npm0Ho5PF7JGMP1EsxdofzVqVywx
+hv2VmnFxPOMHgx9sC60wzOPD6rTnp+g+TBZoZTm/VBvLGMVYjlM1XUmJ0EwCCktNcFG01lxErZi
dZau1VBGmacZu8ZES2EfqVU/WTQ1sl5sCwOFOXQQnk+8eXS5gnc+bt6AUiAVQ7WU2Gc8EnhVlNws
7+2LI3F8wXuRuhKrWAvEC6uIm4JgsHXFy/RpnXRc7xSCWIVb8viMVOHfLO+7XyWgExNRSqL7PO8f
Ywjfi5a++8uSNrivIoSD03ab2W/BYbycxJi2XzEgaIypnITPIOsC6cP4cEA4Kero7L4u4bcfr2ZN
nSA2hzLDiwlKU1v2YS4lFVS1+FBcdkijTjB7gZOiE7zK+K6p5gNcxwnE1DzdhYz9nbvZPL1YDI9E
sT2f3E0y1sNgOGG8s7tZVAJ1FR+a6Iv6GKhyuGv54Vq1/+2ecLUwN+hejxga2//QRCBL4pKTgB1v
igGu0K1yUOFULjAOIUt5Bu1pzb2OHCtfUKE23SA8vLsQZIsdxoa1ZVStmMDFt/6niJiZJuhJneV1
y9KxJBtYlLbVxt6/0YwsGXnyYiPVfBBEtaJqmNqcgn7puPKPYEl637liwpZrgrqYkU/iqQSSrZx5
tneRzycxnObgA0B1vDmqH42H9EDVwcz50L+FxppA528dFhfB+YL1Zr+4AyQcCOAsfgeK602Jw+iy
hZAiwwWvYucUwQ5zeJMMBjdkBU1WJrxf6/aQPqCwObRzHqYQbUfM2GCiNYdq3JUpvMdDcvpKJVVt
OxL9fPmsUygyrTJQQBQ8CL5PvzkFoZoyDy/l68Ir3B3is+N/5HblWKgjJ19/dNs81Cv/O7CbNW0D
Y8vjzIjhB638P4qxcAD8nWUoa4PcZzQz/xgq9DYRDWngPOHpm8rjOjtPfET5/duuSKQfU396n0kJ
m0C2YfMT3LGP5ObTSu22v9QcjgDu75lFmKUuNJpGXhnpixGiYdbibcoswuDwXsW0MvcT4A39TfwD
TblJ9EhLhfBWUC2o62BpPQYjcFnhHOhNFh/ofyZWbUJoY1bKDUNHkt4EWxMsMGcJgBzOz9VWPFhG
MppbkGr1aXRoLYbv+96Ri/OAOF/0aAISQK8O0POBV+xVFDy9Gr6vP5mf7AqbwGsJaPs3ByGlvFKx
UDHSJ/CPIT4uThHORKdxy0Fj6HynGSS2kfQUx2lPjLantUXiqYu52rhE6ae0oy3a1OQ6JmNMpj8G
RWTedhPs642cVd9WJ0+u6kUGM00DvtwtZSP56C/GXIwU+SnHxYl+yIrgpGroAH/9qiJN8E74gmMn
h6CDRwYNCV4m8tN9ADveodLYUeYXWMRgffojWNQAJZ77lTRuPy4pwKKn49vZJLsLiEXpm+u58pVn
rRtDXl2tjdBDVtz+0VUomTXhk9r3VJi3wRkWr6iL7plVA98qoYt6kRI+7XQ3WeHG73sckwnHoqOS
HZTc5xD8bng6AeE8oWAntOKHWdDCdGvmyWwgiEVWJ6KXbR9roPlDp1o9+1BkIZEEjPhfgBe3G/Yl
YCMbYRGpvtvVB/ycrIJCXkSqI3pAU53a6iw/d5SiIhQEY0MyX1Y3QuKww4MbuIpLqQEn8uDZ34nB
532ydz3OawagG+8Okvkidtt2/03zyCJ1IlqF0vI9S4XohN6kFHtArqYv/iTpENm64kaRLhxtWbrw
nJWW/gDs7yg1nWoSCzWSZBDRHNY01a2VwpyE7amA9OftpZ7g7E0S296uNkM/tNKOe1BtxQ2hg9C3
l5w3OfduKdW630kf94Mjq0e0ki4rtRtYjpC6MOlEA0Vr0m2sICdTU+4ifTGQ+HhP9H+AGcZPYJKq
wVlRUfP5keG5Ayp/ilfsycsOW1CFs6r4TcPfrkAGFsrtYV8mEOJ+awCgYG79IMPOc+6RXtfeyvyb
Fz7k+OnlDexMdb78qRHfipWBr2GSuiMOTnxsEjoBqE2+RYv9jYTQowAHd/yKOj0uHtH7w30m/DtF
1ge1UwK2T7qyNcxREfscIeDQGMdbLk5KKFbqvCd/6ReDGXkJ9nSC4dRK9pVBQru/Pwvz6ewWh7Dl
L4mws3pkSOvqVKCH4r2/dItFIJt8Vxsb7syecWuInbmYgEyQ1Stg9jFK5bb8LxdmP0huD4BxwYGn
djmfus0QlOErEDgdzEXiK+Rcyyufz+qptXvCzKz4E1bKQtfi+XkfabRBs839paxgQX5YKRbisSAD
M25AunFO+CPnTUSupCv0OEeT8Djnt5KDNrzsuaTGFlnlYrgBaSssv64qn9nVVCYUTtLb2TDgHNRA
bDql1xct8uUTDF9VkMwZTCT5H72J5fH9+0OgBM3FmvoZXR3iPbiY0G7i7L1Vaa7Y5npzTi5vSiC4
lJiBYe1/qF6/7+kWeLcxGHtJWTxURT/IVJmDqFEicF59+/Y6bxcQNR3mDrfVF+Y1QZ8ZN9FhaGCv
TyXjzYoip00143ZdbokfEYHMt3Elp6v2wz8IkWp/wZbQ5Cky5oePWcu78OCT5rFok7VfE1s7XmL5
k0xcoNhAseArbs6hMvzK/DMyKbUADHv87mMdENDfRkz/3DZQeHiRUMXJ8J3PMHs67q8FevbgLtb3
G5GYvqjVtbDITcGwPmcbBrtRkS8nCJs3k3sXUQnJnvGPmYdkHxGydo/JO/PGM6pscym11O5duDWS
lydXgBgNW3EYChxqp7LEs8RIEMQUbKjb/G+izrWMJn0W1GFFylvZU6xU0BGiDKFR+fklkySYgJuP
MDgf8VZoJjn0EEHPjH4hPnEJPARE0227ONbhPbDQNkfKea1Uzv5jy7F4LWk6KK4G8ZipM4Oio9OL
NiieixkWcnlL0FnWr/5wgXG5nC0+3xWPByyV23yrriXHCdR5F4Uupf5I+ItxPBoFdvih1L4UQ6GB
p0vckvJ0iUxbazAdDON2ucBaYtveOutiHl8Jil6CjAoZBARyeBIcVZ9M0/sma11jRQ6qi4S304hq
avfni4E1tzY3mAiI2o5uEI2Y+xJPe7zRAPdrvqgjtR4YR+RXWwl2DzGNEj+HQxDAwvScxTIXnWdb
8UrQtv2S1IalQ1NbIZgmtWZanpYYJ+NMWyrfodUzIoRxZSKf/55zGlz/SkG2Sez8mTy+InOwpme3
LU0eubm9LQ4ZwbKbs7+GdXUXaxLrGRcItf6jLEa0dYK9lnwW9Y2wJaSaB3t+ng5MvvAN1elX3CLX
amTRQkxs3fmwzJH+YhMiH+C+ZcZjzNpiPWLA/9OUk+bw75EyS48YsUQC3GbSvqOyG6bv1oh0eyLl
1av2i4nMiM6NgiUGiz/uFjil5zgZu/yC2QFBgSl4HHF2Y6KCIzvZaBfXMohmXsqn2ccBtcQCcsvv
5BrpVp6k73R61PCS3R0gCFPD7nPczWaZ1IG7qB51UWJyYPKxnGqTaZ1CIyV64HFgRLX7P1cx33/t
MdvAGvNsMqxR4oyr6k4y+r8lb2knbIAoAPw2tUgGjFPtRjO234xP/mnkqXsJzU89PCOTVX/moXLB
JuiZWQTODbm4wkOZ9chFkJDelmSW6wBbDdWTzoANtstqCcNtpUUoUhnHEsyIzNrQKnzuKW8iusCq
AY9yvYzo9YgG3+BgyQbMB95XqQS5fVqM24zYnQZujunoPssUcdDrirSrpFfdBVlwmngWk2y+Tov3
ZRc4OB+eo0sVHfrFn3PmfygwOn9WG0pBWe9mBMQnnxayE8vTbmSLUSG2Y9cKMlobW0P60BuEk6/5
3xOgq/TR0vDOT11idnvWYhpgQvmWSTR6OQiB2uCd/JJyDAxNE9ZZ6oZe0+sq3x0GWHTY1iZWabUH
wYBDe2lexoNnzyrritE6AvMsqsrQS/DNaDYyWtkInmAPyWRFo7Da3snvmImSDt0HSWoVy95IYu7I
NldNGx4AUb0hVmYltNmrntvRlsbrysPaqRRbS9aiLhAXJcwfsTfK8nNmV8pARindrpLrSgC/gVly
SynH8uDkricytVKvrntOej8qiQB6WPNKj/t3veM0xIREC8sKBDOrzlXVg8PlTVMdeWnI+qizcN6Y
F+s2eCzkSAlePQJaH3mRFkS4QavBou6ruikMNC+AsQdZMVw+usodvfy1Q5EvuvNDsMerOkVJzPV+
MEQtYR4h1P3WX55Y0J5SpV4F6sgOM14EqMtt1o91/8FW82i83rMUfms4l562mFyoUAwmJgfUQKxX
mchnIQlkNHOk3bHj+W9FKpPLeoNuvQI3IxmRslXBAh2EhSArT/JURdSaDgkJhZ3ssJtd6p8IXJ46
5hkycoSLge2iyovggQ8w9+dyyVwxTIGsFB8WT+OOF2FobZy3B5bWfX8xt05YaWXPwALkrtVE8yeK
GolBfmoYzRq2pNlakrAFQx7Dm0/JgpHYiJrimt0/IK9zDto8Z+XBmidK+Rt+MnU/LK7vjReMzEO7
YLMXYqKtkExzF9wkcGLoWX3T/yq5y7QevTZx4BpzQuVOgbrUmnc6aFUxHzHPXVSakAMD/09YYjFm
KCLMP/eQ9NCjOEZ4/i/BFZyyY4UeZXHbjRgqvvk4AAhooVoMwPTvQQ5q8zqd7rTiXpYdMyouWj+1
zim4ptG3zZ1a4JkTCeX6d2F0oZiWUHOwtIj/HGQJmimZ+UEXR7176ef+7QbaNsfnQPPjQzszHq0S
2ztb2HC390R+omDn6DC7oJ1lKtnaifk/ztWDTjI38IqCgkCVKgkAmHSMzyBxNFS1g/L76/ZeJPNc
hS2b+Eg7xZYSJiVw5qBDg3nSn9V34AZs1wZWeiHaE1fmKQijNBtJet8ahi9nkdv8x8+xS6E688+T
30TeRqTwKYlcnmI0nkcgOaFGwE/9+xqS0H29/7ukcPX+xkitU8V3RjflHYa64ov0CeT3aILSiUOb
KQti37TLaxzNTonVzYeJERqFcXX/HnUHCUfrJN0eZDdLgbS8+xl3X/Vfhbgzm6Q/W6LP2UxNKuod
+8sR8mzwwzwNhMLrtNScqh0vORLhFQ5GlEv+hHfd9vnoD0bmNW1XTpcehh2uDoG0WDGdyUqMffdm
LtRiQl9NYjVwPkpYIV3kRfiHBO9uhrZKnzK/tFIDAXOGMkh15cUBKOsIV/fwGOExaEYR1zs5pa5m
8ThMlsnqTlH0eGHVcpBRMlCEU8V0Hn68g3uDbGoPd2xD1/oJ+9b//b0NWvr+E61jPSdbykoVJcOJ
9jQlTygtwhNh1R+VPEOE57fZm2J+nITdjUGlXpXlkPAmrIfjEPwYjnPcfWHAq3gJAAsRVqRb1tlW
raII8f4EI/dgl5bOMeIYpqpBprrTjWHiKqqFui3VMRHkofFkVD9j3HqPP0IC3sYsOsIh/QIrQumS
rw0kh9kbDqS26IhLayA1HlvV5NJl0zBCD1VZq4jfMHAgT5SqTyzAuu8XLN+/leaRIXRAdAHrLwGN
Y4sMGiu4O8a/5FwrsZHuHeCF7PSSndZ5JzGMrNuSZE1mAMWlrB646R7hOtCiyZivfHWEQ8hOqhpK
MxQ4Nm70FLZwxYpH4JDghM9hsjnZnKCBFmytRyt5j30dIZB/k8N23tvxvasPu5JEwuimxd78Szop
UbP/tsZmRcevxtGHFoqSADMUo2/emFJED+afzJ9N4FyaF32V8aM9RZHrpe3A5i0/1k3nbxrB2kgW
wlfLBNTimpuf4NYbP5kpxu96j4h18BL86rvvt2WvPsUv1TCkCa7+By+rfO0JGNbJbGZW3iXT/lTw
p3bBViQkkzYe+fsat6BV/xPGQLl+e2X0XiT3350rbK0rxytPp1qSqlaJpWPd73WPb0kUq9NqYZ1k
TVdRLS6GPH4g/7tYTxQ4sVrzsCZo2oFPctwtfpGeDZo9jkAviCtfp5Uqa3pOv5QHYelMWrP8I+nY
M4ODfadJbgGx8rOp35nUliAz0ftJg/JPuDW/zcwr8ZNGjwjx2RWPnAXPcwpzald+fmL7j6HJUD/M
ngqpDpTCcjR3YGTIdx/xIrYBjkM9Lbk8iIZ6Nbtw8oV3LCEQ3TFFaOmRBCfXlOkUQTzYwLQ9aRGm
efcJVc8bVaEjunDkVJu+GQqu3uz4vm7NnN31S7c9I/wJ7mwp5ZajeQGBCNkSagXmRMaB3cc7iktP
DFUGWu7oSEgRW5yPoHCzBXQoYkmo/tI3dk53U9AaYmrc+fGMmiAjeImp0aRcROc6l77XIrjRB3vW
c3aZ+n2VGgG9mnyMfIoAEpHRq+sK/HCSh5wmHxv8WCBqGS7uRNBXOEArvr8Q1EtOBwpO1X586W80
Mp5y97/XJsnz6K7+pt2CBwaMVkAb6YZleJuIwTwj9tAKVSBwVoHI3ntJPEXBCPyweBEzS9G4Nxux
L3Io/i4gYatF5SdQaujYItyx2CMBQg6/jUbTqHzLXkKK9Q3ggZzjFcJysrzv0m2rcBY7qgOBXxC5
mAvncroE3xAfId7eV3p85KvFlOMLGzB7nBTp2vLMnTH3UXrzZkBAgnJeGER1DqTrMmT0kuFhjQdR
8l6/JBxI8E9NcWd1+6f+w2olnck7eCZRw84c1bJV6Mlm/l8/HgHXD2aeTmQP1p1A7BKFq566+/7y
O1ZZS6F4B64+9DcfeXMTXy65Zf2/iz+7AJApHL3gzxISQVPeL3cHxy33x7Eey/o7DAN7I6gBn+Mq
vviTvMYKknF+4ZO/rlxRWLq3x5PcEpyJ8JVVgYKKDADkxk8Tq0k3xZ2XLTs32Ntg4e/LrekwPLbH
0X2zDzvnzlfqOzuzCYaqDJwNCMVN28xJUH/iaYX7z1hFaQsSZIbxyPIoHjxNVz9ezP43aQzR3FQF
R97X74TBrPSceM4IQyY2OEARgqcaZsE61Wsnq4jDOFTWcKZGM1Uw9V8Lqi5m6GI4v4lprpMekAY6
9gs6lYbPnaqHdtAjDXL0r6Zm15yrkbLR9Px65zi8cL22I6eztrqgtc3x6HqHM8ekwCUmN1p4i/MG
QLeKBxdl6u8S7vtrPBH67FjO+rxO5kdHP1eu+53lVmp8xRKvneXHJMw80pB3R8PBsVmsJXiymmYL
l9M4qSRxRtnp5cOcwCGHwVtRxwDQ2CYISSZGYkPo2BAq3QqAboyd1h5g84t/15esh2wzWX6eh7PV
0HOveW7I4Q7TOAlkF95kPDAP+LmvUx+g9AGzGYmCUjQttCt1HJkAwsDzKaaWW83momGpALNtsOQ1
n4jjxl71gZyU1qX0gMgnYfKAZmm8TPziAnC5UwltdEbXtLgeYcIMvVI9PO10SN2o2EGkC6S4fLMO
HFaryDUgk7/R6VN9EtX4r/w6XdsHXNTSNpLgBqSc/c3DpFEklkGHumHwiYGDTMiUKAlQd/qW5cF7
xd4vXeZVSUh0tadSIuf90bRxNU0iQ4YNpV/dSnv3EMQRRCJ2ufNpc9jnyF7V268x9V6JIak8OfRs
KjkmlfqS2YiOZ9t9a5/T4gsEBiVQB6AjfpepDmIi/We4vqVfsDuT4jIDaa9q0ak0w8A4iT6HGLSi
x6MXzYYphcEgWjpa4oEIt1JG20c0XZU+5RIMr/qr9bb6z/diHHPCXlOYftdJTZfy08GrhbgzvjKB
pbMcETknFiwYeXHnQzmM8ce33zee9vNIPQWH4s7K6n1sWnD+RG4tmA5UHi0AyQxmENmA+aAjrvA9
9ZFB3glVTlg93jIcF40LYvn0lHyBiSKYxH3wV2tu/oBwSmFW8PQDaWvrPgvfao/Ej508koB9p5gY
8Am4uifH25ivmu0bP37KQdOxy4+YyqbDaKkGJAiTnp4LY7TZBsmSbBjLY5UkeV8lhP59qL3jyeYm
msn6ZbYydWa7fv+KLS4Mfvdqr89J/irUAjj8bTUxCHKRDPI4NWoOVvXvbGjaGxkmucvWm7Xw+ady
xJE0+kW3oMIEYbt84a2TPJE/3XnF+6jpx77xRxs1aXD4XyJiEEZmQUO/n7jM3aqrgST/+nN12MiA
srJln6o6V1XZS1FNcwJ+WTF4tJou4wNqjrHhbvB80XSWD/do8/ogfMTo9sJWqxKEq0zE9q1dU7Q7
BzmSCdQt7Uj6zdQFIKQORCTfddD/AiSX0iMzKEV5LFNPEY1g5Qd74Lg1jrG1ZJy/Y0wJvmrZOOnQ
3J5pswJcNeExuUCN4TeU2oJQbuttxSpa1KHZP9xr6umnk0rqw6CYDeq3aeNxGevDZkDMrR7QzVvn
Srz+haRNoMD2t+3hsWph1seHQ0HpxOzZngXo17/kH1bNZ+6XxSpkLKB7jF8aD6pxOOWMxlWbqrED
xBgoTZVmPfEWo1ZgQV+91zMprwRSuhzzkoIVRbPOMwHCHbV5ugYlyypsn6+DDfeZ/ur3YyNqIUBa
4UMI0U8xNrdbNLJ2dUTazO0WmiAiQtAwCgUhPMmUdoancUX9gJx3+CSBn8qcqwGbs9Q30TBYXoLD
YvjuDExYnnwk5c4//U59RNsCVbDgpfSnYYPg0OyLdgAtrIgYQtXwaMkUcH6X755heuPaLVdgbFNp
oJDbSFAQn6n/ocRQ69mc23bQUSMNvDt6XkaXLFI6P+yJX3VvdlfZZ/DTIk76QOtVZ68jEa1rRiJB
jXlUrSgHWxF9/ZYMbUORaA2YgQI9Pz+A3/tQx+m/rjyKu1Bh+8e8uNVoUhzyAAETdlbfK7LD+uvE
ugv/sBCCP+og5jLId5thxbsB4XfRyncGL0xoSQKDxUmI0cyeegxSEqsGnHc0C+9dDgVFX4Mbi3XG
OfXZCqK1o9uhRySxROBZXh2G8HlIevUmN19pnaHqVUGl71g3B7jqUuYT/s+wlEW9MkrwyEA8LUE2
/3FjgTWP90BHCP44mcEoME1ZKEKwy2MmBVZnx9DzP0yL+csRvt9b2e18kE9DoMQ61WAFcfvkW96p
B32OV1E3SAWswFD7PZQQIiAdBAiSWY5xGD7pPF5mfmcGqjxBZa9wiFteAKuQTV//yjGUkNu0+RQw
6JJvbJ5lCcbef9vrITePp5auXuXBDi5fIdcGZLZtDQTEZyX/ygNdqMEOCvdHG+YdI4dwfSUZ2Qbr
vnWCf8RuoZLZJu8hvsg5UYALnBufHpZsifdFCwc6Vse5pNW0nxybsY+dcWS5FupzpF3yqB8bt442
zZlP5STqksJItfWqncmxaU6HSqBISVzEHug+WDJj7ygOkmen5CZ8z8xjmn5e7ILXgbTHvXDUoaWr
ur/G9WQTdMKIUT0fjRqdYxIQt3caE6P1f5X2KZL3Rcu3MTgzv5gVWuADXtGtNSoyHtnlonV8Mko1
mik7R1bpkH3muX0UiYJ2vUQZs2SRmmP8LU+9TRZr3HjsCdyM+izJQMg6VMddtJZdNECHee3DrHrj
B4JYg77xHl26qxsBP1gNDJiEmgzObctP6gaLMhDOmt+HzZoyxG0ttAZj9HBx0L0BrR2LV9uc/8fq
TCNvpzkHf350URfBwjLjd9MOv1rB0cNPQOOw/97Ze6e5TfxQ/Gx+ZZ+k8aris0QN1Xb3gjaQ1BNQ
Dnov+rlu77KuJ9xn7RZp6Y5hbl0AbIm44TAZHW0ryD+EmJPwaUFYYJl1r4pV7F/B8k+9++zJ0D+k
lWe4W21+Cv9QGo3CFhGl3DSnV2d7pYhqVuXeL1ivR4MYCmPHfv+qy7uWLExdMFHTQXOPGRuGFGil
sZCHk1ebhXb8FBAIlY3GGsowalfFXlwrm+TeM4HDWVcGEY/iUipLmEvKkEEo93C7lQYKxuYmxFWj
RNfATD3EJyC6YryDjPC3Hr+MUk3jGV2yJV0+CvTVyPnBdbMrCKTQ9guNiQE3n3L3eO1XIBpl0A82
Z2Txke+Eh9li4+KGbVLp+dnljzyhGp5eKjthrMZkzjNfrcEjjmgw5fb1/DeSEXr171z17glcRtEp
agIBH7F8LfaThIAmNj+BV4ymP028trsjrxg9jlk8mEnnSVCIihb+yk/iDl3BeoHWXXMLfihtmSL+
tKeK0u+3RtKp0TTji7Ls9leYVCwwj/9riUHAqrgHeD9Jon1gnVmnfmJu4T+UzGeSomdTeDdwtjjj
paaytr/Af7dGbLaU4yT9R3PFPqBGd1VtCHsGb7ryuEd0z6e5bsOBzwtsOHkqI97VcCs+3NQ8/Y44
MHpilFEg2OlCKkhhknYS6fKqlkviOpt9zGPu+z+39Wcih20GDAO7Z/ZKEpvEcii0ahHgHj9/AELS
0itsfhmkN2okPzRvvJf7a8Hyf6XmFv0vlW76qHgeHdc0Qha1u4pZ6sSxC0wRO2DNARYKxIi68Yi/
/8AjO30XMKaVFf3QMNDyzZA/5bKEto/D2TmTggm+5lHzPhjbUQBZcatplppnbmIcbwPyT4ao9fg1
3DufKl/7fUSVQjDA81SpDYhmcqwztI+aynv4YA9AjrG0D6g4q38MGyDkdDMmRUSm5Weal3+JeFxB
NQf5Zli2v8wyIrcRntXEamKE+xFeOLye4w2Z+52rmDdGaqBa8r6/7ZKnJBp5T+im/sBkWbffnF0z
7Gg43Al83D4Vpq0DyKkeqDoUR0zEF8xRzUECjkE0puzLVweR9fF8vTMn+EhL1Uz0TzJBKxMNQeZp
bXMn60exhwmc6eHoXXpVteiuCqKYnsnnMtgKD7sNTeSm8IFN3qhx+gtsDVZUVJQwBDUR7ELn5abz
SB08CGYPf63RoydmEPgRE1dtzYWgQ8vrPJLGKZ9IUHRnyp3/w5zfnp+fvlLvO8fWiiLMRV4PcvWm
KjZ1Qj3SKeQlxOkWcDUqzFPZBwQfaAchXb/wY7tM+g1tL2//rEZrRqNijVYtWxK/FYukv3jd1aRO
AqMwC5GBL6RuRwqU4ykzK6QJz5Q12kiHX/nAW/A+NWKzwRcc2nnJdACAk5JEG/eHAvzM/PJfexzD
SjxASNcRvM5lSL1goZjinU43dPBKjSoo82HGG1kxRwsujmFnBNnYPETTWJuBZeffH8wGyU9GafFx
JUXmzvL3NOlN6XkvCOTIMUvsexBmTTOLxuz3o76FoS53FaJzOYky230Jp07ZtftRDdKSl0rPlKYQ
KDk9ftu0mmCCM4PITRK/wt7R8Cyd7WLOFMAUEKsYBtMwYelVd8b8YiL5hkEEfMfihmzoyBwOy0hE
mh5S+EI4XZ+Cp2s2Ojjkd8ExRsiIZccTzANQJPMvOAuvl9V2d05gOgSGVE7yDGoVBp0necJdL58y
1YGZw6YqBgIW8Gcyk6yTMo5uJ8ICKoZeFHi7GEULB5muk9JLnVJdh3znR7EnANsdJrAgomb9YmiP
3u6cB1CRRyUTh2+9dudHe5PBUOaj5oDEPLwFCVmAQo59gePV9/kSTqBOU9R2iwZZw7GMZnffm/fJ
nDFlypZGSxQatDwbWpGsEX3s7PvBdThs/eFfADrzzu1apIGl5FLw80R1DN2+FBFfMlDU7LDRvyGZ
RIoJkSOcUMvIAHjlxv2t08TnVI8D7FHek6UZ8sgUHDZrBVXCuTGbfBLilKrjYKIfW4rmCsKTYV5u
BWr1I5khTOKFhtAvDaP5AiUY1CpecXbT3YH5O7OQorRDAa2UBeP/Xdoh+fKTol4q6fM0G/1JpPVA
mQJCN9YxHCqgnyM2r8LQK40Q/49lmpverASpKv7YImW/B8b77Ilj9zz9CNzhntvus0n/fCyoxCEL
Y/rMyBvhqj/VrD7JyNR38sA+W+ll8BAn4hNwLbMeNEN0YlzJgOytPn5TpPxrLUBvkxnthE0USNFE
vzaiMZz936ydMTzPjLIFK2jcDbby+HuuoVO8kLxBmluv5uIbUSL9ty/p2lMZ4TKgeFOUK+4vNV3m
WgzzM1vz9gf9/Ixi5mliwqCXgZyEZjIs2MHzyakojpwF7lDvkCpXMiDaZlfWuwX/DeRKZd2z7x8g
vWq3wiTN1UWQB+K0WSVVl0U0bLK7zehyq7mCNztNyX9CfNkHu92fvv7hWL+V/SpCIJqEAoXxWiX/
vMv011MbReCmE6iBGqrUvc0L4f2pjERnkyKoUf7qAqHjnXwQbG2F8VsWNjhTU4NjQbDZY7PIZZgi
H3c0JbTT0ykvl36c32tnQc3grVQHyPllh8R6PLpV0Ezr7QfuGY5Z+2oloUWzxkSck3icBhG5E4fJ
DXUMOqz0Ek3l8FOcbX8QTbDbbmz6lEPRbfY6TC7p96EIpiqNnkAjkrhjzWzKbco77PDkipZBGxdx
b7NGaxWNrOAkvJhycQMk/AjXPlnmsn3vtVoSqfF9Rf9cOSIPF5qa6bCymeZZSoyC7rC48XUIuWMa
F4NgxITlsqVEH03dcx27FX4dJnzBJMMdXvmAz8NNj94uhWa5jvzctjA7oKDMwOtas4ESMttjJaCh
Xfl2wAqpFJixfXumf0Lj3uCcHLYjipTyuDkcmnMr9dfnulY4P/APE73iQwHcuNiq1oA+tkedObvI
WXzk+Nz8VwUslXfjqQtaRY56lQ3ZTGArQ+r1m9cKo+eq3cLw5q7xzWQM0axiByaEPiwfcoFp8SDL
WGHsrnDr2ewQQswo5Z/KSpNmUk5onYzVta+XL2p0kHq4unySndPnSgbHzudBkH9AcprjYSvrI30j
KCC2kk75AXwWviJbhwIf5aGKlAVkwXv3JjUZNoknynnMBgcIeweVbgUi53o0Ry59HJLMj+ikiXzE
V6TEcQ8j0BdfiXnVgd/62vxA5kx1IEDgWuHF4cZXl9UlHkGTYfn57+rPTxbN7w1S0g4JzjEcwbjA
hs+quZRFeAr93Bkw3zN2kCvQj4iiC4408jJ8HUNNNULyxejCmvw4wUm8zjaGWjE9AXFcx25UUzJH
kMREeRUU7G3dzSxiUuBcMG3exnQpajjd8+uTnXQpv3hgyBOF9CIDXtUTDNs2QfvxrjtAunxS2/dO
azaNmNJoRZE0kXKYTQ7sRvmzmGg6TYSg9ISBxfmg31pnS6Vegz3n9+i7Df/GE47eKHM/zEv2VveX
hW/3ryat7XQhBmqTyqIE5Ybv/lgtjfycOK/g1YVfz6MBfrRAJcgw7Le8AmUMK0dG3LvO3bQmQB/O
dltmFVPqMGXn1ZFhncslNkVyaCZPKyOOq4ZlQSDj09x1gtsZQWCYpxSV1XD0KurjegzPlHuwIMLi
+ZD6e8TkSmHMwap1WXsPgrDE+sAskohu78ayqjgkbMKm2Tff/E59Ove35C5pnXjI8wlID2P+/2Qk
iXDVUiug1NxShoO0Pmy325WRjne3SJpLQzvjCUj3YtaB7hRhs89mvY4YgeAnALFrKRjLDqiZ+AWM
VtH23/ud2dQUycffE+z1bB9riiK392j/PSc1GcE9nM2bYnoJNMIUK56Rc9AGUIoWdivZj2Ho1Qp5
W+3Z0tVrhsaU+HhYY5sdasscD9E72s8CqrtyPUjRyAJdwiwnL71GEE6nvpEAT8bNjfkZ0ocZpKRi
2Fy2t2225AWkueKGAqPULepx6mBtPSfYXD6AkV6+cWAWHYngzEM1mhVQ6qwpN/n9KaorGzlxt+Co
VZdUmqNB0JwZHQwtYgKbNpMmF/WcNhVN5ylQ9utX2nbMAMGZGKdURRfuhwCQLC001HAloJmdWiZN
Nr3XuJAVwe5MxDdPUB0VOu8cxSL6rd6TmU6vZ3uDQTqJq73IX41se0i5rVtR+qvFK1lSAadNIRFf
lSitTWHiKwhsJMMbhqMFiIzTSZaeXRppM3kGTmw5fiUNPg53Uza6+j/Gy/mLMxipQe8IdF/nxnF7
ZBih63QHoFjvYa7nLpJKkqfMecNifK7/jBYXulLVFnsNjOz2lHsg1AtfYfz87iLZww4iDwlXqCn3
4vi7oL7GxlxBQMvsB1+RIzLoP9NIL+giziPC4wiUFArfht3YZai+kuS0mBUFp9t3SwaNVgOMJxsY
LKuQU0almKxFYgxB86Pd0X8QNpMdhxWd5c+A5VhoZZNB6xMhApcE6JgYvRvJJ6Ob9YtJY2u8xhEY
58AHnEBeF9bb6NKhX52/xVk6PMvIRZH6+MOlapRorNYDorGbcRQGbfQQxkaf/fuG9pVLyzvnAaf2
5M65ODldkWfB4G05S9GvaDpgjQCWztHsDpE0D/jDO6sVi/IEtMWTwlMxbyW9mwJIKotkmFpXYYaX
OKG13wlL/WcvuaxlAv8RwOfmlx/PKLO5pHcHseTMMs8rKz3ibBHz1JSPCibEpN3qr05LiHvTLr1n
aHE5rCVIoh0zVc0luI98faoJNOjkUmMOYu6Bvdqs3i3D6iYYXECTBb3jsF8ph07D8ZH02WYUburC
44glrvGHcSeZe0jMxHrfM7BoddhZayIY/3ox7HBUbXGNiOXO7G3Qa+kdP8xklNcQIpCnweOTUYPk
sO7NyJBt9pgQkW4pUy9TQM39HZNCWiKX2oA5K8mPbbxe1yTJEd0vJAlHlzhITsz6RH+jeq6qZCT7
3t9H++balsbaJb289U8iwAE2zpqtGfYe1m3rc48M83QigtYP96hOaKqzpIA/hs91vwAsMZxxmuSL
KQuM9GBgVWNJqfRvbX+7hA9roFSPGE6IXuZYPI7K3O+nAXmTW4kkTd0PisPQhRTc87sEL7JVbP2W
nqUP9dZy8+ZGzH4hVhKdSPEduoul6Uhu+BcVhkMKXW16BpLEBNL0kn/PnchVxj+RTNkhDlu6mmUf
VU3tUWLf1u6fi2dR/p15bMqtaSemS+cN5v5zipVa8Qzaj/ls6f5C5WAw/6WHd4CQ/QOOfFyOxCEA
MmDM4LY4iIyGoCp7Nk08cQVsGeTpwpnUEqRgNPp99Qj46QDrFCk1My6WIAaOZTZ46ve4cCHwAzrm
S0Ter1Q/yjbe8SAVuBGcZRPx9iQSI77FMtMHIQbqTrvZ0JTwi/NwIZk3nUzAMQAAOMtdnIhwCNgg
0R3SdZq+nB6Rb/Ej2Ghdqs9m9LYeJURZp0uszz/E6jpSvITvAynWATizbP3pQxEr0ofAWJtrHeWt
+OkQUNO7ugh15crR6yPkD/FYEUYOxHvTMiMxcX5esc5uAqWC0VH1u8yUs+r/SMSRuBKneQLgzgEz
bUexA9HHchiTZ2ZnN3Yd6SKQiM6ort7TO1OfNgDN90L1x1cy4AQpzMeRewDBy2InuCVeQ2+hcrKB
amQ8M4YPd9CYboauk8y+rQlOrqCrHD++22XLxbtUJFJnJGkKafubeQeExyMa8F6Ta4m+jLfrM/MK
vNSVnKPfpSUSEgmd/bv4/0Tb0NouvtdThD45cIisXRSxb/sRVZDXH2Q1Isl9af8bZHk9JSwKOuTa
VUd8yKyInzpIHa33N09kmHHZiToeJEEdPCbam6BtZmymr+OdGFCONPmV0pFU1AfkDtfGyK/dab6I
bCFPAR4hc4WwwEdR2BWWne1wtRop0l/9KEUvG0LFvdqvMhosesKWh+bZ4KKG8TY153fBVXbZx7k3
kRwlxdxw14S3btbF46Op9C85ZymkU1vLd/dOgwe05U82uQ7Hhmeij5M+HqqEFXC4e4o5GO8oZl9Z
nNDPrV7ghdDSHYrMLV3j/VZcyH0cFUjEdVH4N8bCiHAw4nINIZqLvSAo4OtUE3lfv/OavfSj79Yc
dVVQzsRTwa8IRAtj4jB+kab4zh7OHTRiJmH6Kr1X9JrWWR1epyMRwDS26YVAK/6mjIiLLS6OzSIF
27cDdalj0j4Yn1nsJY0A+fd2L0oiMZAnmD6nw7Om3qLlLeptfSkrSmDv/rjvYFncOlVZsvQ1yVR1
aFmXjYyhZ/EcX4+opg2VfFxr12ky4bZjdon2g9bPt7FFVjSW6PN0y1TWZ+/YT71HWhhEioRQtR4z
+Ug1PkmZob11g4JuANscqbtcMGka+N9aZJENCD9VHoC53o7NR3djxMA7YlWnQacadTHbnHqPrcds
+I92WPgaUcIlPlQugzWaPMNzY57MukF6PctZd0Vom2ubvqcLtVqJxmhXHEFYxVYxeTx8DT4lD8fv
llCfL1Rk7YhvQcwzGVXVv2J5YJx9n6DUtTTfpYbBCmLyHqsoIeRfAl6p6XJyhlFIXXMR/ltxaT17
e7GqKhXUQ+L84fxzhkcWttUUIrRwIk/ouoyOULSi6ndbIg3mi6G0CuwTwJaBwX0LYTNDPX7G+5pI
m4SGU+gHYgLqEJiHkLZeT1NV18yPZagN4c/+/fJHfQtOU8EQkmpvuPkOAk4rVpJE0cB3N1vgR/s4
a/MxmvFdrozatwimNCc17o/A2TTfIZH34WsglOS1hBjVSPO6EPayB2PNu1neuN5q3zHJRUDNIa8o
6SFXJTxSFVMmOCi7aTpmdosRV/elAuGTUSYEHzaYYJNpoWKCHaTCbiG8oklqHqY+7XwQZ6+02CMe
c2DZtg4ydKUyZDcG7WWcPTsnuZgKw2p0KcL/4YJ7AH4/TMOQlTJsOWQe1Q4t6Qa+E/ci+JlTCjd4
83VRLdMUy3GyuSScmk0ynb15yGP/YDkerBDbrTJDbetGSyCgal8pRKH+YGBRg5Wp1Ec/xZPHf+ug
YUg/bFOvfh1eiJFvuFeLMyqE4iWOPEdJUZ1kt1RD17TZG7dv8XRWb4u9TLRBThBBSGzVPVF53i45
LRqyAEsXCzu14VhSsxYgnV0iEsqKiPzxxMGKYnixm6MaLGAHoZ4oA8RtglfSxzcMGTTKFiBfLZBq
LctK5eZGWC6+Hf517jWPpQT5c21b4UjnV0bE0M1uHq43I0rHrMaiDCMukdGustyJl9VKD07fx/9o
RZpEG351grJcH9iDs90JHYrsEPvnc8kBCLAXhbyRweR2Ty58ExW/9jbW8aQUKS7IT/pg2eBThBEm
Cx5KcALg+R7TWYsz9ElBucirirQwMZgMkNI7rzjiUXKjr37jABeAMzE+uUxDRmEvBluj7xo9nsLL
bYhAP91aSucqTyGNA/Rz75uVaZRMMZDsb398s90VD9NGgkwLNNHWAmOCqF9Zk6Oh9JyQgEDNbVR7
yFKM9cRMg7Bc3pHbTXqXhgj/oHF/WCcNn9z7r7wVDEg5SKcHGLhkldAsyH0JPmUgiOBQdqFKCw4o
MfHcVDm7LKXjEBE0sdZFPqnWbyEm7uFPTxDBJjDUpxgD0b5ou0H1Y51Yd6WnUQL60LjgiV+8sCnO
3bpXOiS7imcKgCqWSwgmYOARJczY8K5X53fEC0AVX9ifm13F9kAv1nQdtp5MRnu6hVVrrq03hqdY
kLwi8VJVlXv+EqFhoiZFpQYCCl34TF12J2CNJnMqoh4bjK0C9+YuUMFRTdDE0rltx9d74SEztNTZ
JpYTh1BAr3Rdv1HpWh00Q7Dl6wfuNwBKMDO2vnD06YlMSHsxa2r+VlBW2TR65hlICCVEnrW7hVfr
CRV8Q0Gk/Fy8hDxRo0qqMjcN35HPz7WTPl/FXcILtjLAkf6/M/li6oiSKbD0ZAB/KDz3nJkHIyCk
G922YI7Yz0ZjHBuMs3vSgOmfdVTDgfhLlb9ppfj0ZFgiaVLjy92LlFbjSdgOawuHtUYYcJ6UFGZs
4dm592koSaEKGjf2fgeuIOlRBiXC8Mm+wI3arwmCxbAD9+fYGdkm2jHSPTdyrIqMx79Ia9uqVmhw
QsO/vBJ9JtypQoG6uNvIp8mhSHKrZqYNx6P58ddDrbiKyjP4R7CQmNAZbD81fX7IUzxF2MZ+o0i/
Y05agQy7ID/U54/86MM9dXtqUXyMlNIB4BoNbT2fNZKXHUwyVv0P1Y6F0E4XtpNNOb8156KbP4wu
v4WAXOBJHPkY8JeO8/jCltaMNYllkZGhf1FLQtePZ+TahK3S1Ty94hwcyV+v1XmTgFkrsVIklJ4N
T2SfPngJa/oqpDye8bJIr8nFiRB36Pba9SAlOWD39e4RTrL6jI4A9L+9T4/4UvunBoma5o2PxoC3
klIsz9rMo9ScvqcIRSq0/Re2/LivBgqQFm77GiCaKfTpo0X/5sePLE/u1M3UnUI4VERQM+LvZQvz
vH8KXrCdeAzOazGtyz4XZu8yyImDB5xNlobDIwcNDjhU7u1GUzN9mMLfPLodb1hShpqsxiHmAMuJ
1TNdab4t1YyaPYzdBppCD1/eS1r9xGqns2Qvfm4UT+lVGRxsG2faqWvsCBrUyo0Ipn1Ma+b8khUH
tvccodaFe6gUn/vh4upxZK+ahRagTYtkwaaggQsg6ECUdRJ0ff7aBU2CioyVeA3w6IMHcj/lglE2
9H3dLw2mSvjq1jhahqWC9pFiQiN41RyL9uK4c2QPOsC6/r+OsXvhNu2ocPAjJqVntNA/btEtp/zz
KOhtjpV8p7bIXeMD/Emiu8Vy94/t3dIda1QOLSn8esUzVCEEcQz/8fuyivPPCff/GTT4WtQPm+Cu
E3o7SldKytPEupdtZ33X22EyGq+vszBbo8QKRtrkhR1n/pXwkCvhVV7plkpqbPP16IOTG6TV9WSL
8o/SABkZ1qG51rfaU1taeqeuYPNNIYmcUjSRSXvBaYUY+8kQjOvrOEpXXw/PUEoAd5e4rjgzzeiU
jILUBhHeVvgaGidDmbEvoHwkhAHxUjTOJhJYCIt44Tfn9ZzHIsulDaJca7QilL2fmHC/QhChYB9N
jU3wbCx+cZ35wsBnSx4J1rgEXV5u8vl10OZCjXm1ll+5J2Qh7nDwGTGLLXFBaBrp0Po02YoaQAK9
0N/fHf5Dx2n7AhXvvDi98M1F1FWT0wyJVXr8JGt0F1D7XzeAihcwezEf8/CXKpGXtc2R6HYoN+oo
PwkMPQe/pOURP0V5hHW28TyfPpkvd+8vXJn6KHlO0BF5JRGpZRH8MeSVT196FwXBmhIl5Kg8Tz7H
7Gqyh/BDJUUZ1oKwc8eEbTR86xCaEaHFgNqL5Lj0bnRc0O0f4486M+bLp3BfCGmcKJ1oOwkrAfIx
brKyf7p7G5mL2x6veZYAqglssU6xxsnxqwjiWrtIwEl5/yWmO8n1Ma4haFeVmX0WPrIi5actGPqj
bxIg/yuch6gBImPqobP9T5LQQNwyFD8E8zo6ajI5aUEZq2JK9SVAlJ6v6alHagalfn9oMGB9tDlP
V1EJgNWDPl6xquz0SnwCuzP/zoARAU3v0YLAmruAHmOq8qt7KP2jElgemYIpi4Nsa3W2Y1cX0Si4
ieyAB7egDs2ekdpizQyh9mVTYYxw5k5fZxKz/8RrnbyUZeYcEmqjgKTWIgu+YMu/iscfJz7guJJ7
sOnYk09ddXLXolOyPeI6JM0byN0ORj7fjBvt2Ys5z2vl9vG+C9WZCBgnN3pZaEzQuBu5mEpP4ijV
ntjTc93I1kEznNWmRepWo2sB74HLRWqld3irvc3Q7aXzVzE4KAdpWhqNyL8qTmtKdf3Rh6XBnTTZ
7duRRjoVjO2o2fPtcAtUoF4ChrMvPiqFe7a6fKQkyau9GS60zayN6rDJZWfxNiKZcDdIe6/PXKrs
UkUFzruhBTdRXtztAvQtLN3kf7xawTCmXzXNY04F6mkJjAbtHc2+n7Oit+NUW3bfOtPmWSkALE9A
gK63BHEBCYqeAHcJMzRy/frKfCI0MYDIO34vMOm2aHj5VYSrerESb/EzuPV8WmoKOBEMrc1yXy7h
GeKSmgBX/uSNxPQQpEuB3X/BuuAeh+WNkrWB//A6DgiMFSGqD2dCQCFzcOLw5XGkBpoNXci+mLwT
VIyVjdk/k0wpGwvTlI2i/33C3Tbrq6hrmAeXZzX081Chw82rHB5OnJGlA7B0EOKVRba6aP2pKFhv
TuykVpujsd7i3RBixMTFLYyYe49ma7faX5gSSeebB1rs2vAk+gTLmbY4jdAXjxNTrFVex7pelnYg
5KqcUe+e/2JTvv3mhzRSIq30GC+40nDuS9AgcP1zjmzmCAygaKnv9yhGw6WMR0deax3eWhuRmGZs
32e6lbRWlylMU4O5GwL1/Q07YewyFO9VDiLWX4dE0O76G0GiMVNCyl9YgJ6qyNCl7cHaEzyMKLI4
8ZqlzwVb8+8K10DcT+a56eAFVqjJ69Olp+jxT63L8hojADGYpzYoqVYdTLWPi9Ihnt95vdjbp3jh
6AdleG6p3Siwwle9oL7Z1rq3fBJE1TCoWE6VOwG2R26qRpp8n8sRh318FZ5fg57B5N0m0BKoIDJ+
wXJE54LaRKlwOm3WKzL/5mJrNQK/cfMewoIX73WXaqo/vU6lmbnzZFXcAZaagbbdZoMiJCzT7SWW
dWpw5YFNF+aiVcohwGnf+uWT2FTkAHxt35MQDBl58sTA+HYSlBAHxZk2V1duRmUtIlAlfWH9v86c
/7zERPHxjAtQg/Rm6xJ/KW44/HWDI8VMz39b//o4qHe4fVjKyTZ0sDyGcV1lGgqRUt4s2zPIduBB
8IfWAoFtbj8xFU0p9hZteiVIkOl6bXI4lEz3ZOmmTG/mAVAALdTlq7K/2qIEVDz5EUCskhxrOjla
50XgwsJynCaGVL64u2xmRJWQo2CwPXp4VtdoQR5wKEXrRrnSopfe1wv95rvrDdQzpUpwRxqZXiTB
kC6bYvY/z6SRZReiFTVQDryH+DIGBG4ORrm2T4vsjZmP2zo0lSB0obUwth3X6+deF4KRTXrgtO9P
3mjSNcL4YVnarEuF4NLTY+reR6pRkqfx5AnMpyx4YGhGL+/dhyouCAW8azDXiJAU6qKMxnxTmYHg
VZSmPu0tNzG1eTz+wHGMCLD6ZZpvze0qdMk1kIA7pagjMhIrRxkg7l5mZT8cBqgC8iVG+z8mZqBc
5zZRiukgmt3YTnloI13F1an0tmRyCoqb0GG2IO/RjDSIIJqpLQk784DoCXySvyPRjxx5Y981Ldq5
hLYCeRGrkk4dxIwDmcvqz8vAqAgTGr2SW3ASbux5rYsXFDYLEVkO+VxrjeS6mid7xxq4Q6XkbAYJ
WsLaDHe1GDG9Ypvacw86F9eedK2GJO92lJ6HdjkrTmAFQuVPYgp9fVap+yuqUHKYBJuO0jOP/Ima
PB5wzuhLwj3YbH9M3ojgmLFLzrWNPDVr8OdBEcLae2cxpqrACHIUf4YBk9ISo8gVjIrsvO1aTNm5
1gGeMC8Jzqx8gPoUh/jb7mHgXypdq+1JU9YY+nrtiLk8SNxj5XXXYxce1YtkExmOktAF/uKzEeUu
jihzl6THc/HTMHSxEh8QJVYvVOgI+LoQEiZoFQetXRKMRQSStHduLVyqEojXu4nLGG7CDez67jbb
ZYgKOuNRS/808/hy4RsySSPaDJEI2GfOR3ww90NARlc3RCHebq15xOwo9yslESC+8LoGsuxFj++I
SndaL/TIxCx2KAUGCOl176HRIMLut06vmawu97PIKXlEYGzd6+Lc6FGh4/J21iIXGTcOD1m+qzJw
icDRomuYFs+/JJ0HKF2zc6lrntv/TZp8h1waXan5fxa31dr5r7mZZypRI48QdLDspm4Bd+stsLVh
nzHR21CnY/y2dcZcCzjdlmvKCZj5eX5SA1FrqsjumgVHFO9fB1kunyaz3qSUPFnyKYqI7NMxPbSp
U9+UpW+gBCRwUhD3ecKbSVoYqV7zAfEh8tkmG3OrA6msb7W9WewValX9vq3aR/GpbSYaW1WNVpRG
pdTkyA7vL15Pii/8gy+foSsmtyjG4pmZFvovhisYFskXWfBNdKUv5enYmkUoaPx2S/33CmoHAWpE
DiDxJScfeWOtm8byxaiEJethqcpalhiDFATOEG7qAj7lTLz0+pw94LARiIzbCgq4jJqDj9K0yoJx
59YnejN2dlIlvQDUpS9n2PsNcZCpMiuXmdr6AxdRbwqGMK2/4S5XXcDwS52NPTHS0HSOFqJsasdm
zkVmpeaQbEgGjtFIACrsgcsB0U4AxMaq6QpGAq+HS918pAF72kd19e+Q+/wUuN0fk/t0BLXGgOlq
nSUu5r4+B9Gsw95uuCV7MqA2OHMc/XyyphZB29q8AVcCb2URwpltb3zCumuLL0IQuSqCM8M2N64K
Tg9GiVpeAxgfUx81T1uM6H5Xh3kmuwXvL0+U3QNWsdHgBy3q8crVJOywJ+lKbNSJ+RqRKew7csPT
yECEdlxTivsiD+Uy5hbEqII0aSWnODWr76BigXyhYcTn3KqTMuhF2iXyRV6MVwoAjCHtEv+QlPJi
nYSlpg9j7M7Oau38jVsPEqheM64A5FWphJAFtUiaCtCso5ZqFugPRl2cbVeXgXlarVpezUecm1oS
hfS4FDvZefDoQ54uZO0NeVodehgwhbo5T42j7jUDzt+Z6f3Kp0kcQ31XW7oDSoUPkX3D/jNugYeb
9WbHCuCl+L3v8M2Au1LG7aWruDSovqR1SK+bzNzlZbCmcHRs2PD1Tc0GdoG8UiR/e3jOxy6ISuro
Q9UOmxFisM7S3asdtZF5E297BMIKaX+pNLT4CnZS/+LJ3gwTp6WxLhJtB0moL/OeeQFlFCyK3Oyt
uQIoPrHnJ1qFwAVgifnpUsZiEpr/kkGCX6s70gRDiKkJ0gWQ3OzddDx964eDe6d248gIjGMEHJeP
xVG/fmZgtF0QYJbuRCQahIz/E5iJy2oCqO4pgOw7eaC/wmaT2qLP+cyXoalxfSJuxT2xkCkVwC+i
FX8usDd9CY6l7AK8zbT587mAvT51dGlV1TiQ6Vs1htf3QI4gTbxn2VzORhE7FgAOR1oolX1HZI74
IU01mLWutTeHOcgb0H+wcBxScnekq3sKF8lY0gtSgk23ESP/1FQWkCzccY56paZdo8UQ+EaGsrxm
ipz123tpMEmbUp6+d4YOk3o10fVR8YipHypr20LgLTDFGkiFwASKOIRMmrvSBAm47ZeSZEfovzpN
QGmAySQ+08P1njPpirM/MBYcGTqdTV6kTVDXR+ITiC3Hv5GokKq30IoaRpns+R3TkMuPeQm4BpEM
Sfir4Pl3dF8dDiqvWPkJMEt6MSqL6t4tbM1oxhs0lHBvX3Yt0mXXrUgaztRhxXkrJ1OYzJVsd/Oy
mefUm0zZNc8ERVbXVjtTtzAwMZLZUPd884Fey7HdnF9nRf/H5dI44EHx+3W6f8oZhz89Da0Huqnx
PvjE5dNymN9+f3TLEOAWggYlgcXirS7fhEdqe7Z1A8s/4ElWKItvKcGe4q2r08pgADBEbRcPrOd9
dgT55CxZgvI1lVK2LGO2BZFjLQ1raR4Jc08eONNMPh6ZzJGGlZZ7P5/0YMgofxe5hSihwoFVTBZc
Z2Ce7Z3vqUDQ7+xX+C1FuM69scvbFuA4OnrlpagpBHsVG8GSOiRVknZ3reRS2vi4gvdcTvjm00Bg
2RcK18jds27NDEPcpAClMkhrIyoEFQFy/HuvxmP9eeCrbraG1bc3Yc1hHZ5pZ+ULU9ux7I1KE3Qg
6upX2I0jj0Rl82sjpYVzcSat8UoEV1Rg2IlBzGMmr2GGoo4rI44+ieD9rw34f3jrcyoQckgHDj6A
rMlBHELPIfHyt6A8I/cQyAHAVUpVgRignI2XCDyJgDKbkDQGZI8RQZS2XYHaG1yG4fI+PmGSviFv
ggnFGDRkCwZ/yi1oPN6Yod3TFpofAdJFgbpsfbwJNKNHRWHRnGnsmJLi9grcjOSzOTGGV4aZBZIT
2G8zKGzshjy2HvZzzUn41uaz/XlkFy2a1OQ4mfIs7raj2PGWzSRg29ppALv8g4KFzsoK2jFIwH2J
0ANha4dGttCcd3yIROcoATo3O9SQUPXEok/u/M9+kX1f7EQJwfJVifdBN8B4s8ImIl9OXcsTH2cs
gLB0tBrPRJvjTkZsf/pcnP0jpwygeyoumnNDIVFHi+/5/s3gJIsX6xhG8dNTJgoeUP0GbbaxWiL5
5EeGvTAu5H8qJspiUBTFTpqQ0OXXopyEAmWSwCNtoAtp+4YiGkzkn+PN0mNRRYE7xCliunNc2WBc
JWmRCcTg13uAaM5P9FfEq+3kyN4kUYbPo4tbw5xblbV1RGzZsoQguvejGQwrL0/ConoZ71I+Vqa4
hPvZd83J6jmKlUXz0S4IzcmEk9LDZO+uvaCh8kdTWC99YYvlgGGQUeiu0zRhzaloX84xKwyc19mk
wr5YJJfd/DjkfmZwMiSuMpObTNFu3NiLzQ0d6uVP1VQAmRWBwl9TMFu8pXjWFuDSAYbYeE/EtExS
8eh43yIJFgUWP25cEeQBU9aGt6bMtyltsLhmGSDvjF6J3GP+vFcbvFMGFevGBXLpPs3SHNwesTnb
tqAdPe/S7AhNqxO0WOwJ//gdjYiqo0MWssxeUDw5aN4uo1yswsZTTejtM2ALSMW/CKwRoAsek/gi
3CfL0gVbdx8y5LgRqQp9TkUPh+3OB2kxwfQ8HtMLNybuc/Hfbg1LKkULWjdatNS8W1A+BIxaIVhL
LQOL06s7f98GrKtrB1c6U5KiMJ+Sln5/yL37K8WwXzv9lhGduX9bqIUdmMMvFHsG/SSj2y3yFLdR
0BJjM6BelZW9vS3zh1Kk6m1zZhBuo0yVV3FRj1CJk1CQogTMwi3GQ75eeU03JRSesN+S/7A5mZlw
/ZWNXANdsp1clVj+dNpvUlDMpiWaHY7h3b8YmswJftaEIrJeYoI12qaiDSjZ9MW76bj24cAtnpVI
pC+fgtWPV/zPQJYsh5MAz1I4iN3LOV01nYH4Du5DG0Mymj+u0ZZ0LEPrwvYxn3xRZBRsCmbON6+w
sJEid5BGogK6DgdgCtB08oi9F2Rl+1SWD2J5KdNYXh4tY+7+PmxKrxw72vdOAFhKCM8BLH9AW/i2
hN0RBtHiUKTkknHybPJlZufsdiIQQ3+rL9ugK6bncsF9U5duzJdAlWP8xsM0ji3XMa8QuRBY5Fnc
mZkV+L+lIwRHl5fdf14rtSROz1kKi20/tBJkTIzx7swtsWcrikCDAxvoPLytzLVHTlcWNLJ2skXb
+2R4Sl6q09gsdWDKTX7Q1ygcZ0nMf2pfPZ31JLOj0TJAgaXkflqA8yEzT6P2cZ7nXdMDpNClzvgu
8Q08o77vsuIWA2JTFV9jh5rkOsKfGI0/zVhu8aZFFBA067iEeWNGJZvzjqHJXeSmTIVLOBfZnwiG
003joi7H6jHSpcXg5quaNwsJf2Q9/LXnwidiNR45eMOv/1DLSzDHCRYh3AxRJl6YaivSollNeNb3
4kvHMeXhQBnL2lGxlB6djxsBqdetuowcC87WhUdL4yHKfpBL5zPog9XcFFayZ5T6Yu/36Kzyi2og
cXgP1ZVEFzc/9jixtRH7FpDLWjrUSc/ZJfSFcTM90XP59UhpxB+tuZYJO3BMTCDI6CB2wC6RogV1
zQpBdl+6MUu4fX/KIe1w0LEmzcR0jPa2l7OKWW2G3+yopuT+szGlnAOqPLU6psFVaT7z9PCYRzCn
vTKhMPPvcp+JsR+ZQ5ZUOmRNxtapk5DRYO2EekGoH/qxP/+iKUQdpKk2XRDw92TnRnHT0jbTuhRl
tqhjMRXjbzzWiOEV3jtshQCMYkAbqK/PLDaa/IXlNRvhh8u6dEW7gRqp9F9viL91780cv7cuTz9I
DjAT5Rqk20/zyVmK85OhCWX6khoRxsRGQ3IwpE1AmiqTt0iFZkP33ZE37SMtO2CH/HK1D1NPcvWU
IPC6DrIM5Pt+OIlNzhCwez24VS3vO1vQ8A+FGG/yEPSq/8fzpWujD32oczwXw8RoG1p1a2PUH8RR
ShoRyQph8BkDb1IPESOqQMYhviEjlPmW4IdDhG7rpe3o2hn4jMB+U0hH8AubTcMpO/E2LmsKvVrR
CWWietQaBiZt4gcRwq7bY1Lp/aKoZlsF2iAcKzmV6UKwmUd6/fx/4lYmgH9zGPU3SY/84ns97DLy
OdUR+jSEFbxdq45a5bqK+k/XXHRRLnEdrtRTCxAtYz3A9wUNyvtD4XsEhCQ1Z9H9jQLOSPH6uHVR
RcCmA1ILe6ERxb6ioMl0RpVdHx8N9SU3MKIKSFl7C/2tDxiOeJi7YVif4ANXMQwpTl3cwKWH/fHl
B78ISPtPOgV30g5qua1Br+2EquMwQJZryWdnmQBjt9/DgS40j1OCILhcjPHwUwD8oQLUeyRwO6yc
xzVcM4qSQ9MJQRDacHyjJz2CWdszingmzU8PQi6lFBBPOV4lTsY226rcXtopYGm/GTDMttqeoBjH
uP2eZGZ/yx6OpgQ8vf+iuB9ghe5RAJRIWvaJ1L8yhYvkB7UCeiEbncLtjwZJO2l+z64MvatZnJjM
c/Eqy0RZ+rTVSRkIPAg5OBbvmxu9GDaEGcRZhI9dbr0hrpjT9vDyL2VhAyzic5P9eqS31yqdn2Gn
iZOtaypHZmfWc3Ze8qX/IISG1cJXP7kmNay/JwvXEwZ+HQdETdLkpIAhVrnlMnWnDs8x854vuDsG
pun2NjLigsN9xKGopZgxTNZx0YE5oXjRiAqwzDLeZ+vsgc2Bo0juMGijCTW3N8lIC6TuCbo6CrAy
HQs6lk5CQGBB8HnVXvKyXxT7v3UP9fvvVJ5iBGNVvmskJXDWjxjzP4AVqwRRJjtF3I0JA0G3BaBX
u0+DEgTLpt1OwWknDbeOTqmadO0yNd5T3iX2Cz5jPmm1LsPLSXiI4Rxp+XTrBpG89505a+0/39l2
QEXJqBkrBdFN0Je+xiVl1YLZugZXay944sXkuSY/0+wXwTC8eB6IXU9H1hu6m0fM6oURLKD64vDC
EJQMjT+tzfh9CEB9SQTCiqrcAROPlfifjN56kM/ZyRXNNV5el0k/IqpzvbxE/udh2Vb+IQHKI0Lp
ZSBvhbTGbMkyqvlstsTtjOtdMapyIU8NeOhits6fGj1bPXeyRGG2e8frokLCKY0bIWblt1H4N/Fc
Iw6aD5zzhTGY53At9judhfKh3ERmor7fVo3aUIjz4T3twOXupVVQnOdPvqTckWkSBH16A3VagTsR
TQ4qbE5ne0DwEwUhKyHJJfH/lSQtpK4OdM/g6tL97U2DKXf6CnmsfSTaS17pcSezUtvu3VvW/PXe
o6UYGnWF1Qi1WMd4Wd1ZvVU4NLnypoMap+npRQr17LHRU+tGfOgWilX+7DWZ449zZEoCsH0WDtCF
MdoRKHg/l/5wONZLrhctQYCsljcO2vCPY2N+weISAyD8+N8BD73LJduQPO+BauyzZJoZdu/Y/jLk
UmVg4u91C7LrwcTZ4hZ9gY3ziVYuf1073xUAaNDIDudENvYy6y7uurz9msBkQko9DHRpeUI8Zk0I
GdYDjgJ/HbFJn+atlzIaAmb10r4Q0DQWYcIEbKZ/WaFEX6ZLQKRGmVytIfhmF/r0/00zzxvGsRY+
1GrI09Kc3Eq/FpQxav0XUCoLpy5FkRJ6k1PmwEyb0b9xThV0qY6CRg9KRlRibB0FhsuE7uOJvW10
+2uBwvXP9FwOkK4pMr48zFrtIH6OcTdMaRAxzurZ6RSmYOxZ9d976qOM7KKbjuk+0CfWFbSJ87Jo
J52pxNchDwm/rTXr9npXDak3ocSeDOfTBQAhYQiQyUxMC/12dD4p0mBqxJteK6F+dd4otfz1tQQn
z6VMNzIVtwA9yD0T8j9shlsUrdVaBucJvdTrF9qwndn75+U6q6iqM90vk8w1v+DgFeHi7Q7F43Co
U3us6dlzec5YLVEwD0+5BYAnPTTbFoqp1GgzpWUVBs79VzAx22ShqCzouvqzc0o1x0+1icxm3udT
3Jcb9jnfmdgj3vYTKeCbpKH9WBUuo+VdID2MKCwzLMqcVG3Tq+2ZRtKUo5Y3kq9Ys/soKblEW8qw
GGWwuyIaIAqi0xbXA9IL1bnNalkCMel5BB/lLMwV4/WGdVpAnK26ZYHamG5y0WQvkSQpwIaq3BUb
Sc7Xy1f4m/9mx1czBKMe20tOU1f4BW/5oMQ3LkPlLjICrRdtZEocpvuqrJechKVRiloMIqp6rdGa
xN9pUfKGvx4mpeSktw7XTQyE03T/O21wRfpNLfWAeh6R5TbwR9ggp6p2yEAlqUb9xGKlqWbs/MUD
T2AIb0+M82WDqZLn1BfxSWz3c3b71A5ETyYCFRMvKuATUYqhBX4lgk54yqjPfjolwHIKug9BpEXf
k7xxHQc8Zp3iyuutAj4MIzzk3brq3Hi3E8X87tFCbNPQ8X+UFoBbLR2Kk2MVT8CwC7p9FpbtzeyB
Rn+8ZMN0V2Kv2K9p6T41Sf+wl6jHjCECtPZ6uuogIuW+MBBKxVF3v6L0xS1Hda3zPPE4BU83Rm/y
dJ8/C3TVWd5nP47LeNcxe3VG5/pYEzFe2jzTJ58YMObI894tGohUcFdKGB4gYji6z9bDu7pl83GC
gpuWbmHTGw6GOoXYPKoNLSy4ElFwoWQNir/Z2C6H+4ewKIzT8K4bLtyVyPuKaW5bFWmb2T3UMaU/
q+h6npSail/uwyc1NI/Y/Xji+qov+Gqr+h5YzyZwqDoQhXghd6SlXQ5fNJTogepkCINpxAv4HtoN
iTXbeQte8Uzdhb7jTwKht6llaUbUJTlGJ8OxnRLHFFexiLMkYWv/OpWH2cHb/+pZnH0apfIdY2lQ
JKot8b5thup8cYZ1VEf8Ot50MHApAOrEGxuutswEeZN7lIA1omxxocB2O2iPw9l6VNviK2f2U3uN
X93jVCjjuYLG/IHi8mhSVp5KGySScx85VRkOez6mnKmP1+mLbik7QynqNgFy7Tccy/X7dAnLTZkA
ljnAMdAPiwPsA9aoaI/XgmWz9dYcb2uBOeU20GTz0m1z1jSpFcOA8cp0vBfiHO47s6ITpEZ3bA3l
ijU5zicBmNLwGDpoU43scV7NTVKH5Me1UAbUmzIq4VDScc+uIQfj5oisGxN5HBkf00X9A2dH16PB
bXbawSkq/X7wFWDvbPMX0A6yv2hIM1c7rxHSjW1WCFIFWg+Z8tGRNbqn9SczFFtWSwA2YAupcVok
vxW5AK+3HM0UY5szyHqJLPJCCKcUndQ9jABXD5CJD4L7NGQ1C1ZXF36CWZfMug78mAi2qqsZFKVo
4Y1+PPdWxLClUs1zf4lYMDGk7FSa346HFk+fbvI0PyolJLtB5A6ku1d88bqvpsK5SQBHmEI3zSZN
5Tdob3Wna5kuELSqESiIg2EasouAWNDqxRqiAExOtOxF82ybUgCa+aAEotketC8o0yfDKAzt3upb
JFdjv1BSKUIlRM566vn7FUu5QAXBMMTS8PoWuXK/2hKTc57AtAEDeJXiQ6fjwl+Ud+ZSoZTCSlUo
1MWeglZaR9/KkYJ6coz6LxybatX0se43LyTFPnWY+xCupYNpNoLFFiZvzo+gYdftdsHIzi8Wr5RG
A3iOp4Qy2xIL6sXUjXRT6UYqHpRz+SqNYrFN9yZ9l1yXvgLisCzhaayOtmQdTE1LiW7Ib71bcUyJ
hM11nupuDPKUfw8trsSrXOGh3EuqHcACdm92hmO8cRHn18JuTMjAg1AdPVnWfkeYwcJhVlRzDen9
YdJb2l0csxwSOeSzaapT2qHRHqLmtN/QuZ9tyghhVu8IwPfPuacgztOsLRW1zVdzKzNkP2r0gUtG
XJznJ1jhrrAEP3oHNa52U/cFM4A6xfSriE+ExIucFD5qlTCM5fXMgvbC/dJQaDQpZ/8sUUYgTGWU
uBPDC+d+RYwojLLhOhyVb3tGT5nCywtiTN7/ijPpMEftUAkYH5l28Ghr0Vi1V4mAGj3D59gHkA8H
9LeKaBKnYlaWpmH9TAFzgPtsyRw24vE/bLN0h+HDxXhGwDCHEXZJ5XwfxMgNf9Qpn7NCLcHVDyQ1
DYFPwAsaq81RhqUdqqIQypE1WRYdiiNSsasrHkgnJVuDPQop4H47eH1Za4ZBpIFZ8AjVaR6DpUa6
6Mrcx/+v3GVzEtK/a3HDFd+b5dlo21TCOnwihHmSVHa8lQK3UD4TQSYgjtoB/yEwQP3EGuvXBZ7M
d5orzXoaeBfB8B3z+tRsxN0RYtSFxwVsQBUEZ1rvBuKq+zHLyRELJVmzPaHrLQrF/Nho88vY5khU
pXyYyKOO1cYtN4XlKRs7Bd3kbNxjUSKrVPMPCmjFQ3EAgEft2GMveI7DkZKAqjB52Gf1O99uSr2G
xJF67OVMYCSNiNcDKeuhVchobdnEwxhGMhlpzLb+9lyAwFnm+Gtt+ejVIhiyy4ALX9q8y/FZLc00
8EGup23LManbBu0hRK8oA3Yma2j4mjHzIzDKRv+Q1inj5nuBfqBYBWC+9nYEh8ucPcJE50/P2Hnz
tXZpPou3wVR0KJmX4rkn3kdbeC/KUtCrMz+jc5CCSUgRsrdlMjxoecSd5DVQZwiy2AoIMVavk1nL
U5ICGX2xW2/grAx89C2H/O9c76JZb9WlKgP5L06zuHBTRdwlU5Fz4rIhl/wWhE2xIf4PgN1U2rF1
GYdWU6WXvoTir2VjopXCC3S/U1py/PxxdE2Xo3NfFzzrbXMF4C3EANIQ7bQdvaxrawY/yvWSiaZS
0rE37cOTWnwX9HtORlkOLiynyOT8Q5CUZW4xtJnkEEAVloj8hJ4UiiSU4zmPOIp3/wRCCvazX2ry
fyoUJHTcu4LsGtxT5Qb34aSaqABjzF5vFniBziAw2FnF2+4gDEu+xLSHn1dPW/Y/EtJzm338tSMr
iSsTJW7HGxpEYTOhse/uxCXSiaenVnspLNrMCJBgQy7tU75G8EQStTjWhTLQd7zTTLeq/q73rbox
nUGNxCzxBHmgyQkJXNKvdnCYlVANSu1vAKz1Gol3N92fORu8N1P2AVMQUYywcHiVHss0jf9csHAi
BbXkLfCRK/XhQryelEHfrZx0N8NMBvL8ncsUjIQZ5jTfM2jTkgWMtowGsomTpaHHUMHpRPW1Whpu
2Z49Y70tWLVBV0zByp7mddizzlsSwbnxEkOQlePPzybxDVNUk9ihUwBlsUnpI5OPOddZH2Cc2+ma
lVhCA3P1bn3l+9Es1Lq93mMJB8QlpzCCQXDe4B/9/6KNCA5UZd/VGE/9/fb6M1eGwKPS0DxQ8WXR
fIlO1QcqEnmrcagpV4cIpzv5F5ceoTsTgb+68AE/OHQiJqE2A/VF7vUYcoikOz/bbjsHI5cW4h4a
QQvjXmcWcorkmsht5ds0ds1SSP4ikqOLZHc4e4PocjxHPq9fkqnDcfIiYoBS6oZAtfY0+4KN8IWh
qG9WYcRkNYTvBHfFkFu5yyHDGyvuUcURaG+PzDikL+QDqfFwSoXsxYwkK4nZGSlJKqZqgVMVNY6H
I74GjG0gW1uuIhqrqTUWmYoYg1dODFeaZbtFw4Xk56QDITPe7QnQkDL16JRP+33tOyM7UXWXzWND
PHXpmgw5RtMfTTGAaneaIl4haFJaApP6bAXYDK+WrOG79fJVN52oA4lqOSWzX8yaDP+AkyEKF1QR
yifCumHUc/LCVADumTQFyzPCkPUQIbggPcuQhdzbpKna7igkiK6bfxmovrTA1o1CNm/iFz2je8SC
GLfHbHYKjcN3PAtFhfFGze8mfldsdBzG/lCHzzK08bp5neEmgPOszDYLy6FWOnzkiQI8ZzgPIgnD
JkIboFllWvuuqnu/IU8d08VaSCfkL8Ml4ppTpeCoDMVm0IjuikVV6lgjUvUI6Yk9J/MLC+lNeCr1
j3yUY5vPd7hexix285v4KetmCZ69fbs8yS6GMVxdbZWgHnn2Mqi9hu7kY4dupwJ5d45d6zqhgc0m
NE8HfmQQ1lkVpeyOr5SPWhkK2QxbQvbTtOsMl4l7GMVCYIFEIYNQUp6a2FIkAYfGOIycxB73lJ3S
wuESsoR31PUsA/kP5SEER/yTPtjCjo1QDaujOg1HR7QxdIIURIrv4REggy178hNNTahNztqcCZ87
VUV2xlDIAIBgWjsEppLRVix1Qvs8xu9Elm8z9YdJ6zEaCAOD6UvYske1hHeJbgExDMJOtZlqPRNl
zFXkdafbOR6PuXMz3gDlHk9T6g4ROVCrISMD1Hl0QKdjTARx0tItqRrSyAOrJ7JpPBvWrsBWAFWP
oIC22AQeUAwzDycwbS+x5ipwE0Lm/a5HWQ6CMD9ZMbwU3F7VPZrVe7bfTvOlHFEFBGcWY2akrRIH
XnafWXx9Ce4zmQZaFWhzUvkGhnZlJhtfNfWpyCAP9CTiBCmwW9hMXbJQCD8lMiMaQdBw2f+iaeJC
33ECBaxwhCUHW5wV1jCS/nlqPUrmq6vGvjI091v4HELn6vWtrR7JZ2IeD6wBJBhpj/1dVKhAPl9l
QV4nYRRUiJAgdPQlLrSV1LVfv75VjiVlPRXjBc+y7hO+KUhkRprUq5GglQILngTZ+5r4zQnRk6P7
kHP3q5Lp7a/6grzQ5pzVoiX4jaA32BazT8DCuAeMePkF8qoObuPWk99qhp8ihjjXGD8iLt8HlFnU
tyfQgyXBrBHW4tDazIwzIZ9TNOk4BmgfDRHugW/Tn/dN37QYpYv+MC5moPwpPej+6IQsJZN1Ie70
qb1ywVyB0OupnDQw7bT0TL0r5NmBy1myIHWExTjgVvhptQC2gxdrDWe9heYCjubWo3Dk97GjE1qT
6vx/BWVd6TeIsPUsDneMU/R6W04Rlx4ZJ75VNnOP+NkO4g6h8ZJbPJMBE/VAKg80rqrI7wAWwMpn
+BZE6ODX8ykbdZ8CyryNOdtZGCmsAVoaUHtQG7RkJ7+T4HWuIpXJuYW7AZNRaD++OhnpIK1mRmoB
E84bVFLLsuwtRMPq85dTw/qmOVJ9o/cPN4BDBLjJjhpzovaiagi6vTj/SkXV/z1vEEdZ8fRZ8FJG
vJr6auwClW7jGiTFuJPeMjlAGzCyJwLZiD+N9zp+nDUQdVhhduADr9+jX6BydxXn2rl8RDhblj0u
cLpoG9t5P9tG0QrQF8NR4s8rZ2bOBmSPhG05dhZwoVYb3T5M6wlieb3Gq9M0MwZBLDFaaE5INoUd
BgKs4XeAeUEWg9BVzBlDH31Zh3AsZXq4bSsMCKyihR0Qq/yg45BeoqWeAEgNO93ZT+K6Llcv8vzH
TpuFbpMWq56gEtfKV3DQ1nQ7jHZT1YXqni3t9zKqK1T7NgApMbhVuKNpyZ2O1P1S8zPmuFmirE9p
wY9XIe4miMIF5jivkgIj1mkuKbYKDtk/ye3ypsHYpX+tJC6bCwNQ8wFwPU5Plg125ElHrNK5aPT2
yg6ZcpmHjyBRF1DHlec0J2Ooj4Lwh0tNqjfqpvCihVDIJhwBuIXSTxDnqIifk/nrox3m0neye0vj
IyqeYjNQfF/fyOtoKOh2I7p6WBpWRoRzILL1Ln7x79hQdxnK4H9As3W9XjnssYR84kISi7ZVIU2p
Rfk+UUrKlEThEZlrYrE5MZ7dyeb3LPomY9abp1EH/egtJnx29RLabAeQP0zgtiHNpTwFBfhV9/rs
TGG7NHAVOVIs7PN5Hka9RwYSby+PyrnkqZdEGHf5ydVXPt63ctjdJ/iA2kj7gUnamQioRFdd3Jm/
SjxJkloX4dd9zCnCTzIxD/xYr7i1XBXCafmcYzKMGGCjtk1SlDsvL6O8Pz/gazsp8piLp80RR6m2
Jc2td8HN+qUsJJ0E2GvQ3BgYzc8JN5/18I7hF/pWjFUK3tQTA7sfy5xYB5CvQW60sZXavqehbbNJ
iPagSeC5dtHcZeLhZug5YMrqAPZSBlFXpVkYV+EW3drPyfLpS1jhJkBGDQJKHyDpWsSexhYuhkS4
W4VWKpLtgqF3ukxyJWm2fWGq/xhxiNpqu6/RVkLWsX+BP+/s+6T4umy6G15h48Rw5x2oCTwOny1Y
JouPMpU1QZs32hhenGTfxEYfPprTsg/EE0f0kbOogWbhsvc62VxanLD1VduKC77COS9c/wrxE7Nc
vxNlg2mFlGEoDClBfdm2E41z7ZxDFm414I1kyuIR0qJVILmgo+LDFZDsemUe3Li5C7JnQGrV72oR
SSgakW8yXiCw6x1KnaYskKYtNNgQ7F6NaiicuKhJSHy9jWMzkOkNvScA6fUjfGcAqtRapx/Za/Tx
t0Y6Esb5kvC8meXkMIERbFpyBa0AsAiJ2fndLB4WwpNhcS6ZSrXEK7pmDaaVPawUcKQvDt5XOrw/
YemECLAaev1eUJUUXCbQqDfX8qqrb9ZHhgd3cZz7Nz39DUd1kFjF0giP8iIdSQU/kO1LJ4P59ngq
3h6Gy5Z/PbILjEDelMvcjg/hYB3jba+N19wojITOFicLHaQLEu/KkrMNgLXMEYdmaRKe+7pd8puS
fVE8fulwCYnJxeqMjI4/8rhb86sMOQi61RDhIErXG+TiELJC5dLSIUUWqc31tv3JLayuWaDilwq3
ljyhm3hPNFYdfZoKqyiDQ7QcWGGKQLdVxpNJH0RM8xA+M0y/hYHnByTlHRWMkcxCuiW4Qd6DbAvY
XpAvbQy0Aa35IbVNnYCsr+a/hDeP6KXbBPA88Jd8HVPLe8spCCQWH5ysCFksvFjm0CX+BDwK1rNX
bRxnkw3A6GwDuNJdam0QFBlMY7mBKNe0bf6Skt+CamUlH7FqE2zRl4qlAMHv2J0BGIZ783DNkWNW
xPhc3tuGMtEXgu+vxk6Of+/YE9qxMTNEisYmYpfloVfSga2ZzP+MtvADy/2/O/CDvUOO7PVLve7i
LEDxsc4Y/aVXw7ezxVlHbE9osNf+3HSJa9YDJykFBQJHmYz11kkx4I//6sbppFEJMLGnD4Dh2TZq
hM3x1xqzoy8uJyy+U2vxTcJQte0ApeiH/I4wnIB6gIvM19LEuO3GKJ5DQetUD9ae6FTzQVowPMBX
e+tNrXGL334cK4Hqj/X0kkWv9oaGxS4mY4ZEj+2y5ADRxdVzBNrB2TyL/YWgGwSc/f78nkitpi+1
pxHqNplOBk9FhHMrMe4/KKYropX56YY4eIxcq10VDqgpcrB1oRB0jUzPoBTk4VjziYVbjHOS1t5j
5UoZWMjH2JnoZsxsFuYbCPerzIBbvDJQw9btoH6vsNdQVnriqWSwPbp1wYkJmhVEDHnFHoSnSYEq
Y2QTO0qZQkJeRKihcLmHCM0Us/TOGXadAGtTmP4axhrhPMqhNhj/m1mPNgEdNtq1iz4rHsTZbuAh
se4MPOxmlCFGuhI2LIRIkoxVcf/ZF2QFSiP8FBt76NqEv3DvOwEFCpztOE7Aa7jSprQKu/bpzKa7
zT23xc2yf8mV5oyBFWAF75l/S8a4Ae6xv3IKJQJLDQCe377aVL2xux6k56+DkVQWNQ5jb8u3JRzP
WM1dpheNbi0cMJ69hYbTJe61nwAayTwvJJQG6KtiQH7rVQWUhdeTXXFn54tPziIJkHvN6bPHhUdc
iKu5QfF+TaQPtkO3rUrJ1K8wn8B1vUQ2wAJoM06RwnTPQWeJlfJjp8kN/kqq1K2ooqqh2345HX0G
Qa/xHMzzCHwMs92a4trz9jsz9jROBfzUw7zks7gzQ5wHHVnT7OtbKf+/1GCQJIuf3bGC5pXRMYvI
rZj1LG/ks01VzJHLzZJCpPYg1NkzQ0SClDexcUbCMP1lqmsuu2sGnt0KgXfLv/u3TEULcFDgS5p9
4GJ9AqnjC7L7Peh+ju4Y0FJxDxitGOw1PGkqTPCjDIR4JKyjDau/YNbJFvLy0w+SgOJpzuzH89rk
lXXxdv9kSKRNlVUX7vOgj9PqM6DzBuje3xrwZ94JJN5Q9ePn0fGxS3aDz5CutggtvrHCsUoh1GMH
CsvKSj/vplJiVaGT3vMWg6LpAlIQob4J++onK68fAzVBZbg/bwVIm73gkqHFaSfE2A9wpI/ZxOaD
Gi9fWhh3phOla/imM/JP21n3oCAyWOU7pE9FDZiM1ix8YleH0/xinE0Agy+OLprqOE4+WS/mIZUC
wrPHea26pirGz8nizH4CVOQNlCsNMmS8y/1W2BHQINz4NTKefd6Ei131ADYH0n8RV6CJhZ447uT/
2UWz9IUQy9mu4jdftp+hUAnJPwur+sNlTaZZZPrpxFOcs0JAf+dzst8532n14e9ybye1LAqx1lPb
6XqrBpvYQrr6qa4ZwNvLQcJ3oXCW7s1PmjF1Etr5q/ZFjBQeE78BPB0e7zVtOfvLOc6/xIE4g/25
aiEdoDA4di9a35CrOsXaqCL5yn2KtfIPwrkTBOfKS7NjHWAQkEhKdooBGq1Jadrr9JAzS5vfNM9S
z6Daiou/d7NvQfIpyq7CzF5n0puNae+SAlcAOxqqiXrCxnw7qblbUZHeB0Z2L0EC6g6N0vDo8Zix
y1aN5YTvvZJDtwuOrZvDOmldUhO5shKsVi55EP6+/afAQ7Q3xW8ABZlJpe9yozeqNMz36b43aOrv
0i4GusbhyKbC0n4Ymx+RPd0jbIArfhsslWO1X1fBSqaxgDXyjEfFXnd42hG7j7/b/gOE3yfRBzoS
+ix6UBllavDKTI6HhR8rg/zym7gSnjl+bCZu/SoN1HmME8k8CPp8eyqeqLGQPTBcYWaQ2stJSfOy
w1q+LyMV9ZucwTSp9G/wAhZFQSQYcaxcTVhQMkjAn/7DIesL3OcLCulW398E5YV7shCSTDUxRSsS
jZP6Uh2U+cA5meVqBdTDazhmxx68kE11vl9VUeMbpKfVUmnbyEtLSt1PdUmSnKnBzBYD9xAbeHvY
HmP96rypHBQTVal4g5L2nBJL9TsCLeOl+lJAMvrAe0Sh5mKVzvmCQlxs7OpHcTBk0sSv2voywfNF
BiHnVRFY4ofTGM94yJ/TQspNlWwoDSKnNWS+DxGPaBAUkzbJlh8GekK7sDlXgrK4ghcmkVXMu3wL
i/Lpo2rit1HaEzr4wTH7QqckEcmTW7peRu0D+VrbhEwBqMoqh40lcV/13FbWyUGrB0wjfaoNikgh
nGZykUmdkVDK7llRygXQwiEm+ROkFrmeWdpiTQK7c8jhUVi2ihuuCGtSdotsArHyaMH3pfcmzEhg
g85SuPRkuxE9oR0n6BINZ3KV4dCb/A43zEdg+PV4sb9SG7yNMwsCRnjkaHo8C2QUW6oIkI9pUn1a
rxAEk5mTTnw4XVYiYVRYok5XmFJiTSv8l5JVVk1fEqHCv5UTA1eeGnSrjT7BS1TAEOAFdljOwkIO
SWduSBcK+7DUm987rV/0AIYyi4csyhw1oB4LKUwcMa/AXBSTn9FwVEfG9ZQgY91w1yaWrxYE7+F9
N/JgDrDP9M7p08Ub2XGmLAhez9tnNqgATHFY6C24ruqgd7YBnu0rce9IFThNS/89ypQGab9dCGl5
4VUDR9vBOqd86zcSYkj5e2LbkW3J5G7A2XRj0MluEbj7BT/jheUupF6XA8ttu4aDdw/iHt1ix2SU
vSch6M9f70W/++InThjMwmqGNfJMsug2J9OPcVABW8YrpC0dqNG0BPzNqDXisMWF4EBu3IZcG9Xi
Gwd6s3h0vfxlW7Z3ODpW/VsqS8DZS4fIzHoXM8FnElg4Y5qFZ1OYSRhCBvc+vEUFAkpkcFRNtc4v
jmJO2DMDpK09ElxrOy9BlpdFwCVzYIp/t2VEcFt4/V7MAl8989p3s0YLmqy8GVXVDyt0mrEmm1jc
ZA96EmiAT0AmKgdyExB019p6vMtaeBZVaGLGmmJb8nhZREZpSOFcVOvt1zBypyxW2k++VBfTevN5
sz88mwAbOVJyYARklF3Nnch3LotRizYnNvbCdbCtZYFXczkpixCveDbqGMgwyHpKDT7MRP4qvDLs
LuhYfrbH9GPLLjZ/FiL+ti7cz1eSF027oKQtnLSXqipJwOgAm0Tu5RXXa7Wj1OZ0kAUNMvHyO1T9
VLtls0rpR87Rb8FiVF3+HF6ZbYMAiKaVpFtKXxroNyIeSW+dxvwxpm4LJJldQwKGZHPc1BX37BBK
Lp99u2nbC8qqn9RFkF87+tnnQ/AWJGKKogPNtHQDoH33IbOUvkG+axGLJx4ght8/O3DiwvRuIxXL
67MvfjRbzamqCQ94sy3ePJZEBfINM0JgeQj6L+OANdvhv2XsIzhZFTQ7PDsoTxeRwy6pQeVGaHtY
uMQyF3Jy5nI3UK2z6wwgSd69GEOuY51CWaB4cukJSNGXMaSZC1HWjLxMugFedfiBN6K3IscTCQj3
mKkd4CUFaZGryVE8xawwvOkyZUadyhFbJr0WgGerdRpEMHDe4PV1sC9OtxTEJHrKpwLBI7TYkJVu
ZILjB4acepnfdtu+DZ4L/Wrp898pjCWFvwNHR07+388P+Yno8PGlWhIuZNsPwEnS0avzB5QuU9L2
8oZW9uALPJ9FiOolrNGEL35IcAATwhCxRJ1nOVw8eiigi8LF+47h3WFbPrSjW1NwCEcr2l7DYyc8
mTtPTCl8lt9caUecwVpMmS+pt+kGUF0OhuR9o96MhSMVJPTRjPIqh0QO4044ZEVsj+Qc7rgCcW3J
f6cRl9QKkZL4BfKDYs5p9NEHXN78xDsQ5147Yf5cN33VmzJ3vROEmCj/QqC02nROFF7PqSoclbmQ
UHA7k2b/3MbId7VIpYaYFaor1m+mv6MJyDSoHJxYNFpHaE30eSzi46bGwgSKrZLu1DN4JgDRNraW
PjfNUoMwftM0k6wOrDvX+GaVEfalvUB6HFLToy26H8APvaTN0/bX5oCJ+ciNqmi0cW670DQA5QzZ
TcFcZhwIPNByvKWcjuBu+eA8wzKA59uySfpAUXpQz53sqfUzSfFWjOsXVmmlglJ+6wXULYwkVOtc
CQZOxZKx965LS9EMIdqFMxfasumnoEQ4NSReQpxBp/p3GRSmpvR8B1JSxeYaPo0zBn/l/cxP+O+2
ZjN0rgQBXLbt4bqRrx9YiKsVp8WRxvzVo4CrWM7NNhKIJjUcHo1SZi9s/pYzWdsrNJWQEiJqp0n/
GtH45/NfKEyWieActIJJ6P9ilPfBbsD9S3MnjFolSMk22iiRa2D7qrAKNvF9CfLjWMYKeHWwreT0
YJIYe14OKaWxFjtHenwNYEBAVnfJM/oASxuKOJuKxP8cKdGuQWTlYlqtFnCgVQ6yAQDe2GDQEaQx
+4WMtSqE4fx5d9TtOERw34ygqcYuVmu865AvoTLawAaWuBLUMDiqh4XwQI4JDEu63ZbRTJEM7K01
W17nSoyjOBA5Q58Y50CpyWAo7UUy4DypArLWBHMr3kmcvbxpomjbH4PqY+EvpDDoiOmbVGnbUwvi
sAJTGX1lJ0Nnh+0NSrk74RpNTNYarzxksY42rs5q5uT8SQLTGqoXPzTRyXc89OaVzEKXczkTgHKF
rHP/t73dojVAU87797N7iIODRLBT1UXP4fYCysXLCN/j7H9gj6mhIvR16zd0sHZZbZ6yqlj/a6n0
JtaHhUqaE2gwkD058t0lAwYtBfmuan4GPU0atGVKdOctnEOzgt2of33iRkWLFSde9mMSl8KAwRhR
yInRkkhbgJ4EmkMkyvPXDiSRpTRyVQnTZsmgKxF7dSwoupyIAH3NPukLclRX29Ch5/LlwuG2PFH6
No57fwCGYZ/GnNbMUNGpWFU4bjnyDKoaz+DCwFr/v3EA3r7dJzRsQ97/+NKFGGAQs2x+VFXCaDy/
EYO2KnY6qr1u1qG3eR4NyjfPRKy5zuTFYUQbUZwqmBYWpOnE+8i4thq11rfPOpodxl3jdIHjpDCj
Xmra811RQk2LVOEBLWhQ8JcGqAf+JwOO814kSIEi8H6nlwlHWxL9AQDQwsZ1swTWIaN2QQt86VaI
xrxLr65OZisxRPP6hGw2ciyLG0mU0DqnsvULJdSrtCV4OLGx6RKZEDpHqJaXlxe32JaHAFI4JR8a
ZsfssD67vPTGxRkKRuFvjX0miXbU3viPsrhuvIoJPSZeSGKM1DXFlVa1CbjSqSRxkaxKml9/ACCc
Jv4puOvcIPuQhHJFO2WZuWcP6QqGQuoVpXNM9DTAw+lrA/nMwKhGK+2AcYsLw84B1OH0llQHhlAq
75F6RhXovXKFNhCUtR3CiDdww3tCYbU2/DgeF4wxsun+gPkIdafRh/g70+w31GuE5Ep2vgubEo7d
9ofUY6LvVeK+Vauynwcqk0BlS9vmaZI2wIAPBgiTIlHPhV5gFt0K0MCtP12XlvHJO4vKp0lAe+wW
932C0UPjIwZjNEMLFTobJR0j+ZVWVIYv73ktVJEw5POwHjRb1n9ndhU064YruZzLhz+IRcw/KvLW
vJxV2SMr2rMd9T42kZqzLuS/t/UW3CYZPGoFYuu3JQGMbuJjJpBDQxDj3BsuFmZldQkWniIyultC
g8HquKTJOCB0oIDgfkqJC+Z+YlVKrB+uhgEDWLlSNUboGsJ3AHis6pyTExq/otixjgGkukZb1JXD
c9s4dgVdUFtVKy7cBkAE7WQG/LO0IT9AAlqVkEz7I4KSMqFtYyh1IMziqLnPowGqc5AXHN7GKEzq
SUDK+8S+wundrw/oMWSJO8B0VuP3H4igRpzqE0eCdBxVgwVZkzyy8m9vriNczikdYGotxbGinsSf
I0BO2C4/DaoXytmJqiFmiArPWCVjL5rWLDVHrkZKIyL5CHuBOXHnTkydHJxn60CAAIe1RvjjH0Kn
IKp5jDnfnhaPb2Bx9TFaxevL66l+FB+9jndLQOV/2RURxxZ1XSWJtiix+tdXasd/7M1XvtrndPj3
pIHEEkXMd6Zh/yd9rozxuqnX0K4jLO4FsPN+W4NU0jj9c/dPHZo4EtOx32PHa3gTVDB/J/vmb4Q+
0w8PCeAyNRl9kS6VoyREAkyUOECobhqm1WkB4i5K5fKktH2V9YUY4jDoovIAL3veoZVQDRhLvred
3cOjjKIQ4rbIaBkK1ZYEgIYAABPg3atTpM/7L2gmXlUl03/TJI2XtGE5Gf30AB7SGlScoVJnQuY8
FejjgWt/TOCuujgmw2iCPOBv8Qv0SU5yMviso5E1mZ0ekMTHbHH6a1bpjx20bRHMBmPUiw811c5/
cVrXYEUNYdkqktloXUiuavbGz2whR3biXtJNSEOmz1oLemFQVPAuxAjXHvQQSdhS+zNXW/rWBinK
qMWPpzb8n8zNtweL/xK6JZgHyxd7E8mrQdiyHMofLxfK8wlau2ahUUj05Tvb3xP66AT37/nNyJEu
SQgcTemq5jUvmOzNwnq1HBDvAQc0VyrU7fYmp2C4yi79KYYIgCNkHOmYhWXSQsvxwTT8Qu2K3DiQ
Yp7byNaxDMgGDC1/Cgd/cksK9myhAYHcvxKPMHu52rcaHpbsniMDa/+cSCz4V9Lg6mgS/wKwb0ak
j0bZmN5+iS9XbF3V9UfuZ2htUEOFs1e/bOE4X2k6ETdH3Wx57Y/KjCWRdvohBfbk4OU1IQQLKXpw
rlDPK7Qvl4IDc/wu6rVNF/RRlUiuWqo2Wx+TCsHe/TmzMJdmem9wYWihGFGYIGpgMs/l+dyB9cyS
L01muBBao6KwCRWh9fjzzQzREJ08Qwotp7BtT5WmTINsNn7+kOm++M5ck2dAtV0SL/oBUPTzGTWs
1jmTkDL+tDp6aQ3Vx2aB061ZLa7O6msMDTsn0kTvMolGP4lzpx0+oopQYxf+s4hzr75HJklX0r63
tT4UKp+GWbl6lu4jTdeOadSwiVhXNXj5TeXHOepjGYwEYA+GX9oR+ap6erTuI5itr2uG7OPnSexH
h7G3GBJDfg0tB+t8SZwbf7unBIDNteA/u0bo68WWNBCAiVoBaWH/rjM5ZgwUSum5Y5mM/v/4Ccl4
G8lY02jc4pS38nFksvOMXrFfkIh0juwK/vUv+EsuhK0atjO/jaDR3YkfvIdgnwoSJhZ+7iqvyfxF
/3n57fIPkosRBbYyOqehXW+0hi1rVuTJceGQo6x5MG7wZyobZ7nvxHvZdiVNPdG1h+UGLuEqRGTP
GfWBTyFMy1XtuxMlm0r8tVBSFaoRSdWVwdVc7xLhr4Kvp8qGWs+u0fDPeGo7SZyg5dKjieVOTusV
TiK8UPSmhciVCcBRoDF7kIVlXpFnTwi3ORWrt7Ao5xwMbmpKczNzR1eZPCD6KZjy2tuhm2Qz+3uw
CWXaoCe+cskzBQWuATNxWjKT6f1QQkaoxpf2vkho5sCJPyQf2eKxWQi9rW/9E7btsF94TTwlVdnk
w9CXgTUmiNtBYq3r5SDC+jfGwetWqP+oUCy33Y28PM+2af+mMHYJgqeWNzvFXQE+/0njljUIuqrL
WKPpAVO/1HdDXxwTl0gRKr0RY/Yru7tjA1Q+nQe4a5hmFS+4qTzXeAvwDR4DfmM3B9Uj6Oddnap3
qznYAR9x4WmZAZ1IjaMIqWdmr+Y+/3Ws8Y75uf8twAdmFwkq+AX6+T2me1UZqH1QxCKqxHjYVPbU
CHq4NFHN6+RkJaz1wXoMJyiXQYlXBQvZStRQX8yYxTCRmSvffOMHvD/UnL/ycPckonuZa1cebpJq
wqC6R05bFiMiaF2ztYaUELHiF+mJr5GDu9aExRVSsEc/qm8cgdnkJA8x2/NPXKGJtEtpry8WbnAE
een4qv1GISBoOi42sT86/qh0hS7n1y0gZUu3RSS8H6lkcEU/HMgMboSAcIEZtFoIYGRLCMjyAiUC
epR/ICZ0qx4qt4ZkNbk8Zj3IB5UrGuPi6+qm92WOBUv4VCe5wPENlcpAdBi45ikfCzDWqxChu5C9
poY29CuvHiLizz+m+sJ8e5uyWqhJ50RuJCBVNaIHSLKodNsdVXK8uO486CJsoAVPHaPwq8kABDZg
I3LipOd21HUPemczrOvwRU/Oboc8TFZBtqLF6VZG1WI3rKwGOI8XTTjJwJNbuqFYhDd6hVUQRqfi
RWlY2NOPnEnMcGlcNejy+dIHNz5/g9pek6NqACujpLVwwibAjqyU/3TpS53SZPI4lsvMxR7PNP/w
sbDO0qRC7/Th5qC1fLpRK9n/KIIAJOygXehWS+k1kdmSS7T5KRhTGrkgXTcNz9SsGbNeuI2Uc9Vz
qu+AKwPWpRYW4zTwkYqrxPwXkZ+Q2ZBdm9nnQxkdXf1APzMzyX5MK6zoL+ZhDhSbpd8mEfPNNctC
U4DLiOa3YNLnFI3TC3r9ZGTFlT96gF4SjFNjP8XFMnuKqGHYbGmJIm5miria+vJTeuPHp4rsBIo6
+Zv9N9BuRjF0nWua9Nc0yS2F2yI/qQymRowu/HFGg8H1S4aly2cIElg9uQYEdiSSSb2X19aYsOGU
DQWgOfIwR6JG22PPGZnL2d9r0N1AwLH2l+wVCKflA/PqE38ltjxHADrYGx8T7KV3Yd7R3LwhwvY6
x0SyF3AnIL7/XQDCjKVJ706gfadkONOs+nUDsOkpYm1plDghpTdueo4OdpEJECXAAsaY4B0CbWRt
3cBAKEH7NkkRI3up3DTOl01N07MbkULTXngHP4HEmBkflatENJA39gE8wAqObMJxq6cXzn5l7R3D
DXQeCeL6xPDjyzEm2XbK0ZxMQBWrf1wI9JJYxM0VbaLd6MSq1NywWYQvrQnwuwlA35b9jXtkHkDm
XeLxXOAUs1M3B5hT4RaZYMCTi2+bocyPfmu3Z+9bN9ny3RSFG8W2/RFrBKh6zW2W3gVfsYC9bcRx
MV+Y/WQNqrskXEmMbqVl2dyUeGXFo1NnJIjT/j/L5EAI9YGNYQEUkYTVWwTvLWQEGYs2JGNJY7Er
WHzPwgyB/DHETodZDy4jG1DXgaP8U1wO3TIm4mmq/SqHxR12J6rt9IJ0FQrq1wAi0nXmCLSqi1qX
DOupNWiBH1bndhC0Cg3D+GEnl8hgfoG97mwgA5IUX7KmFtjemnppWVAk/a2FMyv2kw3X/zixEcrd
0kyJ/VZ+to1IZ6C9XEjaeGnCIQlCjpb6l/qxlH0HrVIzSNp1fMgNztQ9P9vFl/VAXD4LuTJbdLjm
/HtAwOUESdIDGVbXz+Dd7/qGSf1Lk8DiQW1Xgpbh8QQCLvWZDDGWUo7h1rMmTCdQwJD7wtR7bo0u
kACKIYQB6qvRWOsK1NUJAu+RGJGnyv+s+AltDiyroSd3ztpxuQ6oBEYSvk3XQ5vu/CXVA2MaME0H
HZ5FgIibxd8QfVXSdchZJC6h0fMQXIOvI6i8VBh3CKMjLi3tGXKetQVJq+++ftNtiwbeLLA89FCL
0e/dxNvnEShXQ8nEiW9hAsvT5Q7i8rjvSAbGzotusoOv0m5/iHxuDe9sqI6484cRP+sPQ6GCsIgY
LSSL4uGdK4PQTWqqSqNqdAlg/WMXsl0MEpTO4pfBN0w/DXRBlTQnNWcVruXt6LFk++zzB0rQCSgj
4vrKcopCo3+lWpSksTQLpsjUO9xf5TzYZqUb8j7zzFw0f1zP4L6dylPG8Xeyv1qd9VLd+UqCumUa
RSGiLorxM7+P0LRyMsFcoG8oAGkI60LMinPnnsKLb5CWcFV3ZTEVlE+mMPVJownHKGvnb+xavic4
Fup9lT6vydRArMw0eTglIT3TUdxKfQpQKAzpaYi6IwxbtB8Bf1HX+ijKqCrudZmgLmGdIvCpDRsq
ZYKxNXIr2L5Iyley2AU75X3JoQY8SB3Gxg+yXKZR2HudRNg+DYaopiy4jDFnirQMfV8dhDeJvHNB
i+xjU73pUMjt0oWRoJ4G6rz4h9csya4ONPRFobbkvTJ/WfqoTyXwuprEDAqj5dwjhTyaBY/34hLU
wOlwXrWReo7p8KmAXYECzWYtecOFdJrBB1lXl++Z3DdK7qcwIvOem7M9X1t0Vn0f7XJt1OLC4k6t
zDaBUExZR/UtXswiueMLSJ5qp9au331EwkC02PC98ysDc15tNEyn9GY81zaMFYqgvOfvj8QZo7vN
vE2fXsh+fYk3e+30TjeHPPHKGQ3lp/Ibiyf9csx2kGE2zytjf8iQsviNFYilNa5DKpulm1JNnRHq
rgVWWPzPuQFLLGJwdvoHJ/Ki0sGiRrm3IVpip6dbpxXLut9w0RAs+jXWtunvnCjLgQChNoiDXYEn
y2kqNBlhAd2Ibhiqh6melw4CrNvMBRvnt4hxMwuFzqTt11Frm2ZAucz/VL1BCsUfCRtdlbRhhWap
iHjeyQ7VvNSm+YDvHsw2+ltoKxrupZ8BZE68Vqkrav684pFZGd6+4NegwyxoHKE/WaeCU51c8xjq
FCJGpArViKfPaArA3m1fhLExdCsrSXTX/xh4t/56JztaH4L2W3PIjF2520UGTpTJT9mUmQ7NOzhp
fTorjRaKwSHeP8nm3gTRMYFfZZqm5FwkOnrUW2njB0REugavvbApbHz/gfm64+JF3zt7ujjrGQw+
J1TJpl1ljGlmISCUUi8q0taE7Vqb6DZIl4yjvNRs+uNLxRHV66AdZZFUMnp5wYR9+8HHDdSM3liz
lax43KXQ5OrvNDupJz2EM1huOPT1cBn/s3/yZgoqox3uNdVc+rTitwa+7ZGhn2Pwx2oMmxdwn6CZ
JGfW0ry+M2jD+Fq7AiSkAmqXW9TkNp7vr/eBljZ9zGUM0plxCZixNSI7LXcLKy52HRmOW7zQIXlT
6LXDXYry6NoFq1BIKkO4xeTHguFHVgPr/Jxc1jt14CRilxoxEOexcbUGVuzbBYegClY5WWDZ8Yxk
V4DnBfzr4pL/UxMfXoTEqVkL3CHKLcU3ROxUFm3vPE/GkgcW1ks1k4UtpNB1XXz8onkIkP6WNGco
PPPeLSdv6J/RhRMKyn5+FEBgFUh96gWoB25/OEB+TnK+eOo2bLKoX6RokzskUolWhnIPzSqLTvIs
r2tX2GxBDZuAHKMVwBMKmodh1lqH+fGwmsTCP0m9tP4eM06d6kL6D4BYp463VX8hZAtIMw7vHBVU
evpgGmY+B89U0ZX+D3N6Fd9lHUJ5ygYOzSEm7P9P1iq3lVzxLdrjb1aK5FzUiPJeJJvqNuEzxr4s
9STIZzUO36CpNveHCFixnOeHewuXrBjBX/VM11iHIN5HnZH1/waBgBwcaD0YYVOS+JQHBpgOGeUF
CNXWnhM4Sy7NCapGbq7qPE5ivaCfiIsmWs7Ux8UldkaxHiOBxro6Tr9mNTAWiSo0BLJgl82BRGwq
hJsuuUNExAfbBv+faNBU3D/ne1uHAyn6QZe0HeJHUx17fhQfWTflBQIdzDkPGwy46d2esVL9/RDA
dtoKbuvz7hYfqgZ60C6aWy0D0EorBSkJjtg/I0CLF99WxHPGG3t81gFsliRdyCYb43jIyjc6KQhs
M55wy9M/vB41W78R/ne3ZzogRmUM/AGw7254pBWJSfRK+DWTyX8alzUIt7YznFtyMZwODiq4vwwD
f4QW0T2JvL8MGJTVtCmEbLG/kmWxLDCLizHFtT3q33chcc+aseDE4yWLUIWps4ZDMloFOjCkkFqQ
StJN7hX596fHbvwo7uW+6uGXetU29nJ1L/0+rZA2k4atfCLkkaR90PHvs95nxJCooCt+3vPH1Qe5
3f0YBXxphAKWx1i2Pb3by4OzcfgIUg0W9BM3kYnTtMejrlEOts+d/JBy2BZwM3b5vaHHfdK5JGga
lqHVqjy2xgWwouCSw6VtKvj2qivYRdm1ipUYRsvUE9bgm2M4vlIRa9H/k29h/8v/hmQQSeeyV1HQ
yVB4aL+RIcRHEwzh169ziZaSFkMCBpCoGkucuA9IV7z0uHLVliRFjGGq2CpXJ7Y68fih0EN3Uvh8
pJQYXtOJQ0s8N5GId6+uXgPUrxg82fiEseh4+5E0xJpZBO4UMpZOyG1D5aBJDmaIMD+aHklCs5so
Xvjr8pYtIGFUjDiPPtuX0zJB4ZQFBaA56U0cXA1Ym5z4cF0uepukSdQntSn+EgS0eFYlvJ1qYbAx
WOj7TsH1SJNpTMX20QDeHSIW+8iGvnfWqZxbfVcg6oshZ6vc9h9PjdQmyHjzlRVWsCEMomHrozRd
sXMvoLCfLOhsLr3QyWborFKNQad6JbK5T+jVL18aZnvHBBfTNz7IhTaqq3ULzGVbPe1pDWL9olg4
8WlWMxSN2nlgxeXRWe4iARucd2zFPwMqHKJeNhLZVCV5ihwtNQOUTE2e4ZhhRbOvlZEogHTm9c8b
O8+CZqpybt5UMdK2vW2qlARsuJgIl+CGIvOueLI28HMMsQLBD3cLBittEVGxfB0WOey+qIjLyc3Q
Gk6ocmS7cs7URf/Yg9SS4Ki4zjCm1y48KzBxuRY3BqJXkuUegxrN/119pCmoe1OX3hI0ekwWUALj
59mRqEh+ON7J1uhMWPo4soouQK2aPgLIGGbqi+LkGDwageTu//87hicsFRl+qhKrq7Uu5AlAMEbJ
O823EpfJ8YPVx6jX3HfYd24SnpG4UW97KHY4LiJqb1nk6Wc+VZe155zMPnTPR32Zc09JM06z+wHU
NlmfPUXCZAdt1sOeAGRy3W7yyegAauZOAMceVhMa0FoLm7hkIDtwvftWnsj78Jg8kyZTBWetiFMy
/s9BH1Hd8n07MITMgqr1YXZ6/xTzPl2Z8YjffyoUuaYjvvPTHmgCd4YyisDz4nqawwl33LCFgTha
iydRdRWLK6Dgl/OIqprOEtm3u3NtNaJEsx/VKIHxOPbH2LBaqiUAZwr1fTh9ZMT6DpIWTnE8rmtC
t4aq9DBynzGg5FAqUXXDLuIIFbz2E0m69SmR5N35snejDpA4rfTOAQelORoLz7QdDPiM5XIGHRbL
q8uM3ufk5R7NryOm322WVexq+eW9m4vofC0yyoQQ8eIpUltrPWfDrDLK4Nu6iIGGuqRCyRzEe/Jp
CFtX1FKm32qQO34siqf94+KxhZlH/ofPOJOA3Z5tnTPJ5rE6WgNTKhOBEszCR3wwF/b2oGPIztM4
o3Kd84Ev85S/QWkBQc66BWzIjVJeeX4nZJ6H5MmRPNq9sp28NziXYGA8fBVXKlStV4gzEoJg2btO
DQbTVBss0zBT582v6B6kpYQg1n0cw9O1Tewa4/maIF2ZewN/gtN36Gzp/cla5hGu+oMdnkQ8cy81
QYpUfXZ4GS6BtfZuiE3cXkUv5EXAYF3lZi9AEKOs8TlxlOcovWU5c/wlpA33wt2ocC5v6EZnUNYW
w6r20HfhA68+QdSHahHb8jw4J1YiMh2vTv+i2hOXqVgS7jrhHCqSA582n9yHupvrrDUbIiS8Ul45
9zYe/VElUtDaIOxkFznGs1mOmBggWWTbqAB48uyZKA1kAZlvhLE4038GHM4sKhzUUdkJD4Vi2RFD
wKyNsoakl+F0/nFRqc7yWAwWNGXLloi9BlHp0vY6hd6uksbQ+TTpH6frGCNW5ChWvXVk7zkFmgjJ
cKAY120GungYBstMSXblYscor6XaC2tfx/TdATfARMVofF4NZnOHF2L9i9KwxDdkzM84OhL3wusU
iX95pdej6+bvgsuTTcohpKjwFNswnULQLtIub4kKP7iyZlrj5/rv0NLDkIbiWwNiSXKpFLWh5Ihc
4l/9FC/Tm28l2C85bed4vAgvxUPT240xMb9rxsui10Vu3MHrKoD9CCFvOmYGZhnh5wQFe+sG7arb
w1ZMGoiTQQvxjIyoHx6znG7SAGoPeM/i4wwBR0KXNBvZJJj0xpI6nBim41o69mi88CeEOPLPnRzT
bxc0l7Th+oBGyV5l5DRi+tJZq/QeDzr8I4edltr42xy1SN7TeTFv72xbzo2RWG22Erk/N/j5Y5aB
Vo42m/LA0VJvSGMVUNdPMFPioWY+6sE2QKYJ9QWHiHXV+OrNMaw100ZQZ8tXnbV/Yy6ucUbQMUna
sV6DrLv7Wc326ndKr+UaoFnjT58TxcBWbsDGl9poiO88QL3Gfvn5EmveVOzQiGiGflT8jfIp5V3q
4S1UtUiJEbqQfaDM+pGtz7NiCOUtvO0DGV5sid0vStyxWqOnPOX9D/FPK1wCOEJUZ6h13TIfqN3d
/pBzH5umgOn3r2vZOxW4PdgAAF7BGJwgyFdAGU5jhhyk5vYw6w8+ifBs5DRW6cCzQLQARlJ9KRQ5
eEG5ddXUmemiVws9DDNDT4ScEDZxwDTtnhnExv4wybQM9Dbaei9uvuIehn2RjyzHHp+jO+W8sque
uxW4w4JWwXyXrzFhVrIrJRu6Jr7rdJt2MEQozQBFyDUN5naZf5u94ZuFZwhLKqnWhO4LAL2XHYLL
iMKcDblOtDTKGamv7onXNucjnHgWojce+uDlyqrYjt8JjEGSWspWKcVDZh/bWSpB7zOtF93571ym
nw8ujDYtg93AZDuzaXPYLp/q3r11xz2FJdIDBoHJ5ODRn41P43tB+I2a0ogw0d+tBp+wDhQthQOE
OlK6Jpg47+A21Td1EVOsQPLzbVi5PhGQCfB7gr7t5LA5vF5BTwcDS0jeTRajQZ6lfOwK+6Fd80nR
L/lO3OTFlwOOkklfdHbfjkgcyNFbVs6ebWhaee4JFIsnhv2aHT0OvOU8TOHjVeWlVnnJVLRjEceF
9YkWVIPFEHKA+z+ongryGWJLA+BKRkTIfVdBuuD+MrjuYBhoz4n/rIlQ/cJewyEayO/kuj4K/Jo4
+9KT4riWSbOr326JY2hS4Nytde+5Fuio19QfF3I1y0kxFVahOV+1jLDgJSkYXvtJeL0PbYqNmt62
/ziDx5TTZZV/o1XzhwYAG8wr92HuTQvLt0ks8JCKHvelTJHYOnYC1EsdsgLJ+TBieHbGiKe7Vlda
vBL3yPB3THXBE7dsIedd9WrWWU/6iEJAypPm2CYPgcR2ildo641N5bJLlcvu0kr9181K6wN0fmfv
hjl94LfZHP+5zC3M69LAG6SO4bCqmWLzdGwgxkc2UU5/zfysTkBSCJgxZ26IDuavbnGc3IdyXdVS
+s8OArsB+ad76D2BrReFAalmIAg7X3uirH/BnaVcCXiEO6hFLY/zvpOKg3PLfBPkTuojUsDzFnGG
q4CY5G/amclBSNJfBrGuMr6Cvg3I8XfxoAIM1DFWjqbceRpC5wzSt9xMreph71lGM2yIZfxigWIG
GgMiStz6Uf4Vw+JwSYVkP/2OdZLo0T7cIa61Hn9IP41PvsNwZtVpiOlCfHrrGrVM1ZR/P4lzQ4di
CPGvUzwdAZrQ9DwFfftRWIpBcOMNYBfFSqOipu9S0p1IG/Fdt67FIXTz89VGs4StDI2nOMjWvSAK
EgcaG+pwUzXV302/UYT0ls4AKVOxypi7vESUot6lXAHgLmMxd7Nk5I3dR/ubg4HjOHdSXp9zDYc2
3VCbBnlNaoRLzX/IhxXufB3twOcjrF5h5klh17o6DnC5GGs4PQIXja9Cqj8lHiA5Bt4K983Xwyx7
NnyhzmwbJEmQqoO2wE3n5uQnecP0YVlG5mi7FTYob1+RJvDZ6WW3CPZ4N86SjAHitHHsKLpk8LPp
TYhwSEXBsWqhDOUninxEDNsnsc4K23DA80bGM+QP66FInpt5w05X90tRlC0lvQR4S4rxkVlzKPRG
IbuDvN0p9pW0aBAagTDCrBGky1TJwnBBFIEpZbRjeS/4j7er/pCyOqgxLZBxpyDf6V8x66/63Nb+
oa/lu0bRJItyEnMjcWbJyX2vqj7Zvv0Q/KA/Bt2/q47mLMG/hLZOcW5JMldiIukP3i+GBN2GJYqc
k/oFXYwFU4aYvSYdvQ9TGvuh9NVYvKOdplr78ZKi7Y48lxihkM+pZRbqePsfJmLicQYHrRcIWoD4
9N91REc9dnvzNpsPD720sm5nOrv/AqXlTBjGW7tuOXgtF9JatxIOtwa9H0IePMjBKAEfYCO3TKpr
a64kJWDaF5CG1lpm3dSMze4X7WVa1g9GH5X9o72eLOPJXAXOaRALmeZ+05sdibF524zG6jAhQLOD
xfJ/z9QOJZOXql4i1kZl1+oQSdI55Q7DIeVzEjlWycOc8bFj9m8kAxjwJJPIECVYHprr9LVAWR9O
Zz/wZjJSZKxkChXj4S8T2zrZHVd6Cy7xb457byFie+V7roaAXQgpSVRW2lZZLh6DkY/mMFkwtJ5j
54+lpgn1KqYaN2xVZQsD/uHT1eqId0gteT54kUrT9FomG76vi2lwjr48pDtZO1fuTNXHWh99oJjF
Io6uZY1CEY3WGLpNyvhIz+RYPunbUELlfkhknCafovERn+9F1i9zvUh+dEtafewUhB/zNa6gFbrz
JRnppE9zDOoSBKOtYlSPR3D35czfDFLs2tliesZQ1NyWzMgDjNsHLBEeHRFLPqeCwjlkSHQFHXR/
Kx1YqXCjMFgglWgh5YBBZ4RjWujpmJAeKmSQw94snGpIVrLLySdhCPqvu9yFrzOeDUngXH2/tSXJ
8OLknJC5Gc/6NqQSQnjng4fzc4mR1ujSdXtqbqZ2BiKxcpYM9GK4Njo8EIFQCUJTw1he2lHzPD4M
woEPdo7e9Jh0TSWtzgYfB9JnZGc/5/C2RgW9W4taj8s3JdE4ydbiNzs+yssKxCtKMPVNjd5i3uE3
YC5+UaU6l56nZCenJY+UU/s7oNCY7wXSbwoI04JrCUy0XbTtwbDF3gDFJCmTPb7KmOpZ0melTqtU
ty7DtHf9TIYQ7U/rWodDQJNgAb2dJrfF7L7TzvXK9A1WPs4knqYtrAGvexGO41zQcRAQkIsY02oi
p7jaP1P78RMaxgSHLNcVUHCNeEwv+1HD/vPmlQ1gdGlCgNYlgu4DUJnd/EFmV1iBDF28WUU1Dz29
qKPID1HNuE34cqA5i0ANo/pFhQh4PQZEsoyEs4q3nPF3aBRBkPi4fggwv2p97Cjr1JhNjgnHH6qa
+aFcN1Ed3awncsAnoue0RRdXmhhiMbeMle+Mp8ss0zUQUU9WeFVqLE3ZS0rDo/2ODlLXJVC6s7cB
RWfCACSO1y6SzfTN1sUrxQCDi4yu45ICUHkPT9pJJTo2LY1FU/Ixae+4UdZVn5i+vY6z4xjdgPW2
Ez1Jg+Q8JZltzAjM/SBTMNxGpS0gPgBs5LncK9EqwWShoxKCUFkAd82YfIWedVvb7gSV1c5lpzXW
8h3fCGuIHgTMwwj3CiKstNtLfwL1Uv2rIdw+f1iRelHOyE6WFf9NgKbhX4cEQqwhMm9RK4huuxLr
aBvkcSUxJZMuMCkd1SWtcWHtB+sC7yY2N8dCIGwK5PZVOWbHpbi7m0uX7Ycd+lJb0bN+0oe6zJDA
FX+87CZi5vAKJ+PihdY+bI5TTveiB/nQSdD3/xnM5YKxe2NO3vzeWSAjbWOwQ0wOPWyBBwg3lWJR
DX+6q+lq3hOz08KrfOOnYq/VkctQhojpHnT7TTc60851u/mkxNUkjUp03PqYzNyyb1mq0BI+Dn5D
E5M7ik+jA0mC9fX6S7rvvk05U9abtfctP3v+jG0ADHxkY4uCFCCcSHYNcbitMcdT7+wsHcOnBZTQ
uuN4/Vmak8BfYsDPWrP1I300RWoKELJWqoRuEgu1HVWM5zwHu4e0eNZduIkEGk0/zCgx+CtLdgML
Wvif8KGxTYUWQcDE0AZ15gZ0an8JKYDN+WTkjURqic5OKAxjF8s0t2qcu1XpbUIJnM82s8uMaRl+
LzBtd6Z0fOWZAuwFMW7TaZwTRl/yzYrqsAQZMq93y7dptDzQTVj2pX+ivorNE1PlFQ0pA/Thz4G3
DLFL6H72ZDRH3s32Rzqq8TwzkHouETzCbVpdQR0HbJlb5y7r+BInpAE4KyczHpWjU0eVTuf2Z8zn
Wliijc3/jcy6PbS1cWoO+o9tzvDOmmGZWeHfA1TBwGWxa7xGq02XPmpx6ZOdE6Jgq7QcxYlZNzl3
B5BSzrJ6omYNLV6iE7BeZl9i9gHVVDvAYI4x3Oa/lrTukKyBbWvKo0IstO3uSuVxFyq7yNFmb3kP
RcqYi8456uzU1PFbBiojp87LC34XV37C6E9T9Ns9mm9BKBJKfnH1a+z7gN95Qt8lNQtnGPrQPk67
iNZrUIi3w+QTSXa2EylPuhgYjzH+qaFVYL4BllAFNrlfkcCEm7NtH/mFbGd/rror07/zvVZxE1vK
nH0lnyuJcharhvWNPUIP2UNS4YttcHBFzSSe/NLuWu9//j2hlpJDoXWUm8PlXjGwWq9WPVFSUnJk
BzuxnoDaERwNYVLA0brUbR7DoIOa3ZE9pTbyeOeLLQ0tg0X/SvhEVXlW14yTmeNlFJgPG3yQR4Cz
tOu9x513Ra6xY0VDfRGCU9sYHltWVzpfdYcO6o5gfx3icIa+U9cswvJxlLHwgdM2rdBSNsyRKqcU
Y7WLYHC+7wUPD2swj5Brp7e0zrVgdztm8IvAo6zTS1ltaOe2BbWA9ul2lLQo6BqJIrJScAG1oeTS
ML8XhjKxbjpA1J4uEAZC+UlUdbwF3BL/60bee4EAc60ZA4oMpzneBhX1/kA3a9ZELDplmZ0hzdfR
JSqs9nOH4e5z5GXebLPseBee4U08FimZgFJvLsNrDsIS8bSGoJNk722B9LhunnT1Hrj49h9sbvLm
UXkgMQAQ7Jdz7qw7gBEDAc4WlE9ZYsTgOC7MN491bSqVpTEG+CTNAb4TYe+63/QSB6UV3FlhIQAr
1kca60DfwZ83UEFuyBl84bPwK60M42BQqJ6mfxuedmT23CsdtfA6p8NcJzO1ebMtPtDSS66h5G/U
o/WzRY54Hh4vmoW9gGhNQQuSg8k7DtTajm/xzR7qf8n0bLDA5Dd5S65b5mGryGXvf+3AtAxyIgAN
FccOWZ7+augHolD6sqPLT5lJUs3Ro2UMgm/3wQ0J6horT7gKvlofCrrw9mtpS9ZkZfVPrWTEXtt4
Hj2QNW9BPWrMn4gnQShix6IgAwiAvSQ5/06HMu2JClXO/NOsM/gNUaXv7PIQ8ZOf76QI9LB7EYI8
4zpLkGjADwpKuMbbTs1jZcMS+F+yc20xRKgPUc+VhTtJzdRQzEMvNIzWD5GcWjvGbLXbrQ0Tz+I4
9b6bjb1JFbqjnEp8pj9H+ivZBW/nvXffDO4Gyo6o9gOPJIGOiABA9bZhXEv0VZmHNsFnvZIGXSLP
cbBvUP+eKX4Y+21CjBf+QddbAxvxgNcQw+D4aVX2QQALskEF/8BWsZrX8yRIc2RAx0uA4cLgZTc9
9LkJ2k88y6opmXxTstCg+lamMIZ16HTMhbPtvX1M6658vhSWyqsLWOToXyWiALNdIFk8ky0eIHK7
hquKu+ez0L39t8okvVJonI3OI0KR/UIUoo9tshx6bm3Ry0qtE8wOThgxYqdrFinftmcNRCRuEH8T
7eO4H7BOfLcyyboFrKNizaYQkbiMnYy/1Elr+mKEwgrB3Yk8BinDWv4GqVfwQpNq3cEEmmJLWuad
F/fERW832hw0cpmaIDrJIk6m6H5iewYuzbU7OFc1a/R+aOOPTSE1xFKu8xDqzb8gIpI1N6ZLa4I1
gnItAOx0dao8pRlWvftYNrDWUT5v5LT0pLeVxC4XkK3GcdFahgPZveX7mFTcNRINqBmxZvG1HBP/
ov94zIOLGRyPglZnK591KsWBVKmyECnujQsZuHfAlJfeF05q/MpUW7noTH3/6P2/pC/xBevK9IfT
Ox/JUnwQPMPDipQBm5ZFj4UK4PQzKWxsp45QCY70fdk2iKQ7WPXWayMNnEPZTx3UY/X0cYCwfgh8
JwkIYWsl2AEeE6c4+QYikxhReOKACVkCe+lnUAAimb7OI6gWewP2XFLat6kIsn11L/UysaiHC9vN
w05z6uZ5hlFzxJ9Ddq49jWli0E3F3U/slb9hWMR+ebllMHl7+YJfpOuC/Z/j5asY5oZyAy21qi3W
FGQkGCNwOz6z6NfJAs87LidZZ9SjKpvUzpLIvB+MWTmLs62lUTsJCef83EVb1ocD+xgzMHHStAyR
FQOtDjwu7pguRq/q/ennf++6OuKx5FtOsreJiDJdb1QfrsA0tqiw/0Xf95pG2eUNKyl1UKTaTW4O
5PhUpGUqxwdyYv6YOA26US6kx5xepgIe1JxWyHouCz8T2GLVfb/ae2RdjBVSHKcNSGTVcxawzeco
JaXU5vetHEKlJixvBxADMmHeYPc5S1LSX4kHptzsNxXTtLrKydGvcE06+rFZvtj2s3QFUQahqw1z
JJEDqY3XeOugQw3BWQJmRoet1TH5CKqODO95136SDrIg6uPjzNvPKJbR5WlZykD4C7k7tbvlHTYR
0/ZYSDfMHtQEA7lr68+m3N/QOdJVzSaCte/6EW56Ii66CMQGBxudQ5ni9A/Epmm9OdXlnVfzRCDq
i4NnJ49fLNY31gBSaxGBwzUwsr7MpqOpET4PQLJmTxQGfD9R+m3zQZ34/vw3AGutvbDRh7hnqgkd
uf/s5a7iBc/kiDyJSWzRvm419CaToktfn7tip6uqHIhmVN06oeTDifHdNZG5mwj7ezVANJfvNcjs
ascJ8cL8g7OQm4MwM9qL4EU32E24jsT/cRDCGLVQHcKUI3sN9U3rAqUw0KpCLgzFdejxWKBvCyP3
3ZAiqa5iekeceM/sb7UYsiYLnFvz8NCDPEX7W9P7DtOCszTCoRy9kX2T4m9b+ykjcwRN4R5sisqa
77toKLccLb++rgUvDPv/bhnqjkkk93REHL8GU4E5bE14Fajnkfc+jh6BZmsWiuDDhgHjgWFWFTMR
txcMnGwWWk3EpwxQK1fUHcU6ohdLnDJSGShUd5IVxOauMBSvzutCTq0xX9VTOipTKL9tzwGzL81E
ax/jTuMPKs4NK0BUAgXndsHRmskFBdZvuZgNNv9kHGaBbcOg8NbG34rmoyDII3OqAX9pjjreGodj
kICbWgVG80ZufZJ+lPJAFhNkPll6UDrC42a2jOL8XSntAxaqX1pXOMK65Hh9AQ/AluJIAiIfKifT
vPQOMnsSCUJ48wbgL5cpD3CCnZL6HH7veIPTQL3IJGhGa00XRVntCqp4yxp3oCRtWxa/0x4snu/N
pbPmmNXr3syP66W5Eb9Y/NNoKluJxuotAf7/vlHSsDzwpePcib0+P7YJsdX27o+JbkdasicQ2ZHt
qFJWwL6cgmaT5w3y5r5bzk2CobvUAsjJzOmbjrDEZwgVY7pvG/zjxnp5HXRK4WeS1A08JjS/f5YU
utEPbF1SqVheG9Ntzwr6P56Vk59Dsw4K7fuwE9FKduvkYtBvw9XdJPOmwRq9rmRpWp1En+S+0wK/
g+dcsdWKXtqNmmO4k9iPS8DUOj7tjKp82ZBO1L5dbad5Ah7G3kgcU7UkifxQqJEUy1srWb9I6tPb
D4GjSeTiaLk+HDWxt/5FP2eFJDXaXBk3VzwgZdG+LeiYzj4KFioFJYaBkGXVj7EKja+STC+PhFDY
2nrQDVQQa7BCl0IM07PzLDPv4I6Pavl3PRqGQ7he4EhK0bXgwHr10ZuTCumi0cVv5K+w5NfuVG7P
0UgGWVOsJrm08rf7FRdsYcVfgiPq/n9Dk5IR8gkJKlbs4SXNaN3tn4Cu6HbRFeHnSVSCUj7YWwi9
h9QPgQWgQZJgAu5Xy4YlMB8PXEUJ0pSu0twpYall2RLBqpO9qobknZfx+FWMNbdDTz7YULHumUPU
e3+MwtiA/d8Xh74Tn3UFM2ERpJBLhGQi2E4yjQsbwJcO7ybktFZGdwaPcQi03vIGKDrIm09P4/T7
SmSoWUEftXicoMRuAq9txKh78acAFEUO7nZbqjik3H/leH0nq/C0pcuY2TOE+pC1OWIXiwoZ56d2
V8FmPW7KdqGXdG8riu8a8H0pT8jpwUmcWgTu8Ig8Q6q2wfyJ30GX6a+NIFlyS6uv4PCWDhiKUswA
cJQpOaKA11FPW87TJrmAUqagOKfx9bOKlsvIQ83QiKjimvHN3IfTafcucBytIetbRRC9ZI9KVlMk
Yc4epYVdZmpA1A9qjbuPxsTlW/30fNkJfuQnu3BdN7pKdE5EJr7JrZlLEBvvfpOUxPmlcs+YO6xg
08JjSt+Wj5b6z7S/UBPpFdZzid1TEF+DZEBQMXa0OH0DsSk2iAsuawdNaWlyAcHN+qDt+vSTKIQv
XF7RbT8GKupR9/dq/IzoYXZvMZHoR3gfdvaB1YQo6UKYZ7xInHqZ9EkuSLHaKf9axk46Jvsxzfyj
3Ic8xX/lpgcotGkqIQ5L3IlZAzpQz/CcFwC2xR+NiSVvc2t0YMEd/Bz1tr6gNMT2ZcVOB9H2DmYs
F7kdFZEtxOo6tzZGJlJwTZ3sDxIj09HfL9cpLEnEH3dOP7p7oNaef1uUrwhkgLX6hgSKGCW7qOlW
XzCOZ7jLi9KyF7vdLhNM7qazWwxu8fdqZz9A8+8On9qqkaEyCebFQJP7cCKK5co/aI5IdxQSZ5nb
LhHoyiRV1Vwh0/h3ypCPEmTsn5ugvPTArb6WqBll00o61ySZ12BmlqpWBqVVYDvAURekuk928osx
bpeB0U+Q/IW2oUibCevElHdpbb37ZjBtJJCQX34ysVw5s727PwLE3liLSgCW7A0Or9Aak3J850uo
Os4uUc2bmt5j/x5E4pey+rjKMMwlhTnqNN3soPDp5GKfdhAcwWKiWh3PrpFAXtfeWSSr5rWnf4ik
bpDX2AvN9ufMQ2/XJnYeUcAYIboRE5JwbjmY55zaBuJqeUvXoFuU+WDoW5hdTAfmQdmXNhFus+/3
nhSvKnyG+zyTx5lBsWlni+qE1W6TV+F/O6zrDz+r6vFvxrFcyX5kUqgnkMmHHZUeGMyjk+du1kbU
dLabI9zMEgW9L9RVnnWh0Xr4LnZI7NcEXJHobHnLsJ23CureFSSQ6hOpvry6lD9nhrARMv9/7Tmi
Z3lvT24Sfettz2hMkJmzRyOwvLP9xB+fAp1586fImSRR8scjXzuSiWB4nMRrHZx8Zj06+PS95Gru
AN6TG/ZhastRnY8HLGR2tTsF2C7uGeGZCpbDNhTeyxtMO6q4p2pRhxe1+eh7ZWlva2JWUlAyTz8Y
ZvileBEzJ491R92gmhYrO3AMpeQh5EWVQDELp2nzWIXx3zPLGr0TzNJqxnfEN7yqBLV1RS7PpV1p
xxMxBTcFBmq5ezYa6NcMdvG2uNCz5qwITCSTSL1YWWOMv8qisqp4F7htI7nRBdRzET0hYICl86ML
mkJjjoJ6hf7zmVQFGF7aey+UHhqQW1nk2ZAu3X4aIevOwOlnSCzz0fyMVOIdQJlPFtST9/+nuYKk
lvZ+ajBN5tiH9qFr+EgJfLPInFQpixn8c8HN5ZszksrYyQ9JQz7Wf3VkHNx+jeiqcaFc/AwSbCkx
l6QFQ+H4ZnIOLgUAMU+PApMhzqEoKAZxBgMiULL4MzMdSBJWwXS5OHrOFJARgQRsS8B9+ZXTky2L
R8YbCxqxYa9Nz/Mp1KkcWgHrsoGVCJvbqHt5wVHES5eeNRkUB/IQEmdZ/VlXNvCLkxui5tntb5im
ABdjqCW3i0oCS7BYfSY0md/s0BaHrprQn8kd1I4VQinKgNVAwf7piGD6+pq5TnzBSiylWg/oNm1X
9eoaPJdQMx/rD7392EMU1rvNdJL2aRs8jiNyoXw1jxiUJUCvxLb2JAJ96qJYTcW56n8gT/pi4gLx
2rGY6G19DszpktgaLxAkWybkhmDK7En/pq0JUjUdyYvDBOhuGM4eq4jISG4DwcHHWYXVUQx7h7CJ
mJTmqPIrJlE+bm8Uys68VV+Ya85gTHQ6LJaLVqGjuS5Q2sUy5NABloQXkUJ1X0QGjWsq3e5P6qMF
KMpJQjri+xpNxqq1RMqswWeWJy+MV2AhxA0WYhyq4aWMw6QCgtJSLeS7QIOVjqz0wwUwul4pN/OP
G6h8GlMK+O57qO1HnIv8ujHjkZZW4W75LJaE3Ab3QhNCNogRn3jZAYACh3r2z0VY1fxrv5QENJ74
DR2j8FwFFZ2crWsgykkpkDZNk4pm8pVkbSJ80+qFK8Lz8MaSCvfJ1/sp//s7Eo5vROQDgNSfrY4p
ADojuGWenOM4zJTTBqey36eLeh7PbWev6bv2pnKcAZiU4x7DTZQdLxYM50Tr9s1Rg/YSyaqZUTCN
Nd2VpefP1Jg1U1ebxsS7BRbxUUG3Sh2E8k5KwWweHILYwr3Hpw4sO3WVm2ZHVfFCFLbT3igeUk11
WymNfik7fFhqbZo51FYlXoUrHhTHfcT5d4p3LFRMgfsk2o9o68mEI8CA/5Ga/HEO4ZDjkf+HY5dw
+HmXfn5ebdgrK2uAnNTWAfu6Z16KB519HSATGDBdv7eKwr1nsAnRAmYX6OVrkpmu4FQQScRCmdfT
YkOrjRwJvXjUy8fY7kAdP34ioqKFwpms2/KkWRBF8wCqktu0RQBqnQDwVXec2VJJLZ66cHVOEPHA
8j8OqeWXIcLM/gPHex2KAw96rgwAYVSJFO6P3UrzfZgyDHGKdhwgfB6LLYpRRL1ZshsD0R4lbsqu
ryXR6LsqXScZDVaADErHNlzMDO6QjzI6gq4viw92aN7QfhuVdYVEf9ARriipuweDHPSsZEwBGUIl
LLaKlfNbSN20UpjfJCzGD5QgknXjN6jsaxAsGSuscqAciW5Uu3fT/hniDOkrzs2nxQv+iE7crflx
Dkf3A0tf5aQWS6kdq838PyTU5X+oePz6t69nqtlRam7kMRwg6QYyMGlwCgXkimfI3arBQVZO4suF
KEOLzd5JCV5zuDmJC3e04VYGhsvmKBcMqN6i+QM6Oz97ma4QJhTnuRTRwqxmyCigFRCRJzdjWjoL
/O1OIfHogVQcvMeFkeNVxq2kQOp/Ulh+FxzT4YZm7r6YNqsA07YiIxN0yyWk8iQLPEO0IOE9B5DI
GeuRL8evHpBVOt9rUUJdlwjy5y8r9JhsVx9Zb/12b8x5eYPMShgPXovsCRDdMSb6pKmgb5wxBmy3
j7zbS7pgBo2lx5gFRFLr4X1WiiVIjdRIKHIp9O77xVljdjXsSESiTDKWqgg0Aj/q3HUMc6v3rGLG
wvWyKrtqxy7jRM3teF10cYkM2n84DkbYhydqFsHltdnn5S78oL7X9QS5COufBgsTdHkD05Am/GcD
2SSYwCFqZq8PA8ZMgeWhrjtC6owv4qK0aKG3g1wlSsVFs6QfCXaA7Iddpz1k15uqWC/CdkypmSC+
PGX/VhjoLShCT63H+n1pOlhrDBfMX8n3mCrg6CnLf/DdZx2g+aCR2zQtHlsmRQ8o662C5WnX8caW
u0rgsqjzTJChAhhZO9cwI2AukqFUiGcObkHkA01Uc/iPuMM5NQx5jwsohlhO2woPDtndPztJ7+Mx
yxdhaKOgOiWY9/IQBVkKG7OVQj9h728TmmC2zMuwMAL91wf3IWV218tLNkBKyIG2Xbbtp871XSwA
Jra8WW0i0sbuGSNarRRUiHDcWdYBfBLe/Ea6qCaIN6XhCciAp9IZMSRuYSAzfaBuuKP9YSdaflP8
jPyL9YudOR39013JXra0dq2g9Hg0HL5zJVtBMUG/eXi4icMyI72qGTX1yLrG5EBHNLTEJRnSMEHO
6J3KMIi7PYMBIcySwstHQvPSL/yjjhv4tkOnBuyRuWX9FRQAZVRCG/Nptf1TuMOXiHHlTkcWjruP
GXsEwbysQp4ebYwJn2Mg30NpsIhYcPYD9bueeDE3krLBdcHsjNXeAlFfZu+fkkZ1UPjjAdGPDsb2
DMAD/PJgSOsrTFN7mAGsx0gevVIu9ahqeJXi1N6kQwB/6aHWdEVnQyIdN2RUVta4CL6Rc2rC8vKZ
MC/pXn0M/a3Vlnmvm7GvPQRQ5HcQKRXQyXu4FIalIZupMpYZoQEvcF3XIlyoQcxUP37CdJ/ZbfTS
LiDT/xTQJIrcovCAgNGUxJ/whQ8ExdGySOmXaEvtyFEHRJZ/uPk5Z6cmcEyD5QvLRgZbU9+fcCXU
qBZbDtIAUMwdOZJWMaABnGjlkjX92lebg/5pntn3bjYgJP/j+11N3mMyRig+KcetemK5D8AqHYqf
voypD+HhLlGyzMusVRtowavYLV8cx2BDEkpMMuhOlUlICRlpThpiSsJGe/iH/cXSs+g6eQtIIEfJ
wOx6rRuLoiM5v2w0ssffgQDJJ2FPuuHPOsAmqL0+yisaUXKvCbIMhltq8yvcP+iJ1/9wfuJ/RBWt
qDvzLkiboNfB0OeKNekmJJnh/88HXz4CNcjA3YpVn4BIiCXQHhZeAIF7eoxJsGfEY79ChiftaY9f
27LvR8DUY6+drD25wzhgEWUfVl/nhj/skhdCoAl6thR6M2c/yo04xKM+p5ksLeiMr4MCbQ8cdk2g
OBfJoAyHWN6bhdoQkm4k64puvWGdpjv3bDrFLvq5cT1nGUc0+yTgjBSXso1912MlaXNzBIUxlaHY
QQz5QXc3c7xhXlnIk9QhxTve60W/Gpndn3ixEEvL9Qk4+At17C4wmpimd8+G12s81d+NIEhDCJH8
3zWhPS8DJCZXdlhp3l6Dvm85ASvCaixW/m1jpND5IXooImC7XDl7NNx241BU/TqynK7kMD1FUMn6
/WU6Ds/ytDMIaqX3JG9GRFmwcgc2neYx62+7w+ocPa0SqlES/l21pnWyGkvj/hYSIjMM6v5F4HFY
JBo8mfXtZq60qCeAKzi0V4uz0KQ3JE0Pwv+2D0sp97dVHXM6c91nfxc9vgK3YKSKR/G9KqJx/M9u
KVOAePZHIvNUnImFz7RszsJBy6OVlYlVTXDq6RPPT9I6TcV0bJGf48vEvs5EAdXSzlYTP5GNYgnN
XjYtJBAsfO1BW99iNXcDJDtMSoSmdI/EGefiwqW+zedWrMEW3YC4fWLY4pSxJt0kJOQIrNzmR1Yy
nRiVhshj6/LVEzF2x8ZLC9S05HqQFAHg8RuMqZQixdrZOlYWjOazu95vPeLifZn2MJUIuhLE7e6S
Q7ALXM2NuiBUDLTGPEijfZPfi6M0PKaZ/T6mhjhfDx9FJcL2QeMLA2Bk4Lu5wZCHZatiJH6rjYKs
QyuXATORkyhLDt7dadcXDlruChL5RobdbcOzg7czzF8iedppRZfXu0GcLJmUZahWDWDLUetBg9Ix
YcgzYWJ9hM7LTl4Ijus1RD2tJCmLuA2mbeOQSn4NNEjpMwV7NE3kiXuDdcsKkEBXjVeQBQ3PmnWz
lSEuLu3Zn3+b+9gX+sCblCmk7giUjUB4puWEMw5wfr9/L/6/Nq5zHDTE0DuHYh2OiBr2DsQA82f5
nfZedyQ9Ws3Oulzsr5d/InPERpF2sZ3aQaalD4CrSovsZ1E7gi94U1elvO0BQ/UEcOWBbtwhBVRc
oFGvs16Dg3G4vMsQhi8sVit00KgTejUPRzMcKzW8Z+4XPfMDSNTHvvPCvEP188E3jiKN3YqP+FNQ
O2XtP2K36wlL4ifQeja7nOeQIpNyg4n0p7jWbbfgy3ce4Lniid5ZFwwUXqif5+z7gPgqoxnQasAV
cxEYqUvJ8R4rw/J+dw/1hpa4XpO07BGcpCRLwzuA7JdWCurY1LQinm8TtG8RZ5LjI7NEWnkHOBRN
N8r50eOVHV/i4ovkYTTIlldpTjtMqlrf5cPqoHbbxcivZWwKQj2QPo5wyfx6u98PMDwIfLEJW+my
9cQNbJBaBgMb4qAxE4Fy8jMlrSLwL/knXfFNu6K/JIwglFk2kkNUL9DbNs5r1EWV1dniOFylTjdO
IairPnAznRYa67Xh3/0L2Ah2BgLHuwg2a/R+2CK3TsYOB9DK8KxeD9+Oi/1ACXG99vWwcESMRaWf
vT0vFk5F0JxUhgavTGIiwFeGF049+1Z+U3MKQIKVUvvZ5Khq0KAWd+bl73uv/rgDmFLdvaULQV2P
PJUyeKz6AmL8X0zTs6N8aG73ypJcZpV79K2mfI4mMaNGb/ErqlT0YV/VIoRw/MzM7miVvNoJhDhO
RVVz2qRYQk7RBruxl+Y5hYnsU2sgNH/4PPaEN3LxMYinWwYDAckvNQ27dJmRHKv3ETmeUhaFv0LR
+T7lPHrP1p+4S3qHci7Kv7bKZMB0WpOBwWehqvCBYVfA51MDxcEZCSVAA7wr8NbqkADDWunXPy4S
e8Rfpv4GlrDZisJo0q52Kre3K7nN636q9RMyGNtvm76d2yJiqayRHqAHrDT3wvx/VSBVELTF3UgK
hlYPm3+V53hzjM2JIA7SfBtvMLib1R+ostLLsW7Ar2lpqVlU3+kT1qkXqSVvXeQWPUaWDdDzEhc0
M29TqKi+q0InItqeOy0egAEsnypJtjxuqzkIdKxAC0jAfiKMQj08wf4Mui4cqwP1RgrRXxPqZwCV
ocN4DvR+adY6iPt+7Hmp2WAwBUUKS6abU5DOhPPTw9SwL6m9y9AumSNpTjnPzBAdTe6uvumO4U5/
HXek+T37X1mS3D6BRf5dKOola3PYpmqBs4EQgL9q1VI5CSYj3cf6ILviiHmPZL5J0YkSQy/h9cLg
TNRxdQQ6AGfpMlNKVr068YAVJrMsU++Vi8Jed4t0wjX/nYT6p2s5PngqWmm5Fy+9nP8sHnEBhvaO
aVEKtlIWT5c4r7UVI3KG6uznjG6uE1+kxuBww27ZSEu1thK3XYWTY0H9zNf2xgAKVCrBNHtQHFoh
XDKlczpgwxGzxpF3/MoxcB1I320Tw4dJI390nEYpSqH9KY+ySH5hcHa3T4XnnGhKXG8l+VLuFQAj
X2rY+hEXhmNRwP9LwihAVECGul3k24U5PSGAESvQVElnXO77/w8ty1BK+jD2nw/d98vV+2+gs+lG
B1RfuYeNjFpqaLPxmpd9G6u/vJnA+Ho7ATNBLUYwdDtlO8XznCclpDwUX7tohgv4Z7LJUG2ohFVX
xYEMAUNhwCdzjHFkojpr8xp10vUkXJ17IOo3OaYhOTFRbf5A7eLzGsm6ksQvxCAxND3YNY5KFViu
ROToyNULjgczDeZrEdEQE+xvJamqoxhn8LkUOcjisEj/fbjSn0Pm58+CmEgQ2VcR8TD7p4TGuegg
e+vbrBMiTKJxoQQxjUGjK+EFCm7YrkdPjcPrrZE1OcLoLmok0AQzBTFn4MByM0M2PEsc90dxNU4L
LXp2nBV0wQo9Mn0JL5K6Wt6+MdGQt5qQ7FwM7bapfUdNxUSxuNsMPw2DWbc5GZ37GrlvYUNdKQMp
dSrZAHxouiN0r9bdWPVk4xAKfOYNUvl2cnWuSvSc4mJVt7cueaSgk8u4HDpw50gEQK8xzMbNT321
LxizFBp7YP2oX6yRZbsvNglPaZaLvGujayyWXdcld6E4T0/EfJcZ71agpFXNuOz/8BOXNWlJ3tSQ
6y8kXFhch4dfUD8GEMOIHPJ4q7fovtdZw8K0TLb30ejip8Bd9QAW7KjHfYDDngRmc5RaZYd9wDG2
35gZ1qMPOr74HAXrpvfmLrrIUyCgLVbU6bX3EQxsgpNqCvmIiULuYDl4xbiOgRdXYcUO4vrNE+3c
dP58Eml5vEpvhSlp64hXdHvHdZse967cBub5XZS67UYHGQFPesGljzxNJo0mXJ80KLE6ylyc4o1f
USF/RU3D//v0RbuvDHbjhmj0hsXIZqFILKEDn1TW+EJ3Ol9XEIbq4IPrzNKX4d9SK+ErOXoCpRgq
74Rvv7dRfzwDw8cU+u9G/w1FseCHVkNdlSKguBRNcXX5EhjzIs72tw0YKZg7J2AEEkNodb2YlrzL
fgomFIbpCA2Pd7udW4cLiRjVzDeS3Ca4Ii76A8+amebNCRS9LoyYOLNoyv4k9G+HhYZoHcvNzpcz
gJLjZpGFClZCVqZMYKQ04oNvpsTEdrRr2GPGMzHG/UXKalziiHS/wqJZjgO1ZrYv3ffUerpFgIy3
O2PomDACOjtwNGSY5GQ5eIVnEn7EHq1SriFEifnDLhF+zIqDxhm7a+rYdexT8FWGjcGhFCUvCJsT
IEDJQlGRsnf4xc78CbNkOORC190tDmr4rp+Drrmlb7UBqQ22mKQuAd57kzQt0c3eJDzaO1vKps0k
yn1MQZm4uDLYzF9upN8VeXUyEALLy2KhZshqGYudu5S5QuOwgQckoVZ4yTdSqrf0GuiwOqKZgjdf
eVHRVShGUZm1VBvkCfY2TADeE+kY8wDt7ABA8Vhc2dGzh5PuJN2xZVTgrpWRWKaTYXE00otFb3Us
KUf890b06hOHiEoD8YvwwQhlDY4YK+RKowTMEcX8aH75g3wdhKqg9iD0gej+EkQkTO7oqB9zz3kf
yxoS0m+xzA5DwP54/8H1MV75NZcm/NdyoFTOYj8xrvu05dkFl6sD0gASYFuS6q/9OVw3ElBtZCY6
T5HL4KhteOM9SOXg14Zv7tbM5BRpZGIbHw9lrbLlFiVnwPZBMjoFOQZ5orr4N1QjtmYMjeH5pfhA
QaKCiOXgDlISD8mjU8lA4rpiuoCs4EPiz39ZrUXU/WxuOewgtLmkmTsB18pq3InqiJrvGoTJpsjO
B3H+LUtwdYjXfFC3AWncaI2CqDHM8Jje8sijopxzMBTW74X9fbxnNnUASbhQKS+nDAm7RM0TLDHk
om17ctHK+RQNIIo3FKTYTZzr1so0g9cB9JA/FyhAI/jfY7yNVo5YZZsSe5erQGR1MkTRBBUaOpHL
doCFm8NCrCKxgLox5dlr0X0uzfW3fIXr9M3hBxMD9BgRTcec2ybEnGpbtWp1BMfFnjESqB0Cfp+I
6N8GRGBAkaoz5v13Y8iPGJjquUTvZVmOiZfvBOeP8Y8AVtawmmO+jAgDQTBmuuITzmt2KvwwMBOW
FeQOzycG7/hUAG8ewDS84NKYZXFbZqUjNoNlmwvVfaf4bQD35Pvr4+3DdAcToLoy0GmIP+3bv4y7
qWol4qXwW88gOhCG8eRWJI8dJ/C6NvdtLBVwGxHrHpXVfu3U6mcvOyke6NkkAiIaz9vIvBzVm9Nm
8Ft4nUltmhH7OYvvb1/obxJjlk/ow1fJq4BxOuyGeYNWaGf0zyvHryaVRFCca/3QfJeYdO/FFtWF
+rWmbSVC8DhUazdvQ2xHXt7hBf2bsZtABwEQyHZi14GqC6Z0YBvWehCIanXEgzojBwr0AP7Z5EHO
4qkfCjxiXn05HbuFmeYoN1S0cSzFeyXh0gYvn7Q0s0cQO3fIqr8Auwr9cuZTw0KpZ9uPASfH5sql
Wh7hfQKWcNx056I5zJK+5mSkOZKKYp9B2IYc3cXsuNPUfn2SIJa/IG42IcHeC4nfAhZLS8QZAdEf
6yPc1/psz+2JvjOH6jWgZ/DGmYu8m+hmirsS/WUyYfD/59dA74XMpr4oqBp/4bL/I1LVp7XMSgGZ
BGd52SlP+ZQBhPTX8ES0J8k2/dRnwe4Tr26LC5Sjz0H285jFaKUgI7J6+JSzWOb+po1oc5MqGwFA
WImiPuEg2SW4WdIbmmNpCeaI2I2HP6uB5j5ebtjZgWP75mVyxyVbro1mydicsTrmOtWkMTrPuz9K
vuRE21l0ugnlWZGOM6dazKEU2asFPE4ahoByvuBV58E32WuB+ge5QFpGqDnwBl0GuPy2bnWo+n4Q
/fJa049owC190qgIN9LX843HuUHhoGduc2UiQntKIoYaL1nUC4t6WTximBN6/hMLwkMN9cHTPMDz
B3+VpW76t4yoOyfniC6cpCjFHXY99KLOC9n56IJhU7WmdIdrNAq4qROA9aZO6trz2vSANpCFR3hP
bGTUsoi6C+6M8ebKd3vdzCT1UJNQqCh5PbQQx5GG5d/sra1qREzkh8F9lXByLKtHYh2DyS6D1XBt
6sqwBaxu3+pacFAvTI4Avg2zdiHZRKGXyOSNzpIdhGa7Aok8zuvhxkY1zAjAWyNXbWVH773H0zAB
xeR3d6Qa82fEjTXzZCx4TblMkKmIroSjjLkmn9gc3YdsNyV4ycvpLtzbbmla8rPiCIyde0gCo5Ff
qcPTzOGxKHdriaHhg469mjKRhOAP+6eMTMlurRLnzHA0UY0FwfKUWJWQQp87gctDxViS/Bi79Sdf
5gCn+gWpSMHEUaipOW3MQrVGa9tyAVNisMEAz/GiifSRlayaGmEtuB2rkvcJD04WVSAXpDhdN9Oa
XfxN60DyljlCNdJcl2rV+VD/OyNjRLO08LMsUayfUeVvd8vpkdwJSSaTxDjzo6UKH+5uUQ2p0Q7V
JHmpmILTpGj5DFwgY4L1YdISPoQTf7vdgQnVlk3oAwamcjzYSurL9FV5xNRWHF3EtO5wYJa9KS/u
FtM+wbMfsuTFLPYj+qhj6ABT/Fhhi20oG2Dn0qKCCgKOpUajdrN1srP20UUJ4PbAjK2QGKJrTy7H
Yu7+K4L8Kgdqjitbwqa+Ey7Efp40OJ0+8xWbuPOKVGVIPNGcWhfbGFClO+a2lbTwxqwIioBmSok/
u3ZbBpUPV1mkGwEKJArzNjQZo0F8q5/m7j/DdBr8R7NQNDluxzMrBv17m63FKQYDW3lSqwdxOiS6
qKgpxWowPuJ5ZrrCPHxFVeWmS82b1RTmgG4LWQuMG7JIz5R/zq2OwpAbrTIGOCoLtX0jf+MCujN9
aiw9zcR/vRiAAqFdhrUZ29vzyJR1ldwZkQ63vCMGg1bhKI8MAdOvWOc2LcY1AEunb1jk/QKHWbh+
IIHF7ZDxhT3Jry/AP8GfxpzcCfxf39rine9DtBf16YHLaJ7cfnt/vAZj4iJAneF0e76MNFfltvYX
rYCdoGAkES85rai/XzmRe1mUBob5tiUR9ZIBJRtoD/Cpo/PuMDJVkMbw7+BXBvW4D2+YBYmMRT3p
Yw+l0UnsiZiVRS5VxCwCQjSCdDmYxWzc+QzgLKLzVHF5fkW5UMLJ1dlwS7CdnWMMt10xY8QUM4fV
LrpITqIfjw0U0KpDRMwL8Mp2M4NuOOlESJ0iTa7KJmi2z9BqhkofpfUMvfHjH/TGFAsCOx2rw4Zt
y1eBdVpjdI9U9Dhg9Moeye0GQ/bCfXCwejX+k0QcBqMkXD+MXpxbIP3YGTr9V6mYLVZHSL3LJkcH
nLdGI/1oWU1HI//PfG1DBcWSfLRV1kZpPnNwNospxARdc+rfavoI/md/XzGVdQFknTepr8l8qkww
RERPO2LzDDilFggBx5VIhp/5QG/JkEmxphLfHVIQAzJcMp8T19DMqLgqRDmNxtgI7tCS27nrK9fX
SYH+YSZQgOrsRG7rp1CervoBw3Qu49KH59HRaLhu3sscA+thE3lExcg9mZswWzhq4jW6YyJckfdH
KqDh1XXB6pRHD89ngL+yswqZj1Q1j3o4LMPwaKblY9AvXndgGLwBkgn3AVNaIW3waYuHJtm5qVUh
66aRYVeFdtX7fz2zPpflSC3atEc8lLPrHnwhf5EH6IsPMaqFS2eq9OxfhEBvbZYNpRgDx9CAmsIs
0BVkictPp7+mhqYikvJl2SC4D43B8PvG/vrMz+c3IbZebxZ6y/BFClddQRv5k+fW/bSV330zEDhr
baweP0RI58+6kHk3F3lDMwWyy8bpUDyABOSfrA91EdQ7K0EcVa18txcV1e1feI8HFeHgYcrNPHgN
ltBA3cIXBKxApA2d6+WIWFWWm9vz0V42fWUnFebyihA2yqYeYzZY14yIUl52i998wOz0nH287sl3
qR9UiVfesK/VTjWAY1k3SqfWPw0UGdyd1F5aTu5YqDQFM1Bm0ovCGjpyJIh6mldFsen9QV8bpzz8
M6sxuK0QwVS63UPayXsg0CIP9qh9tGdEN9O1Km8jZQoV1SNzyI4WmSKB/7D0ojexbGwRIYh6MGvR
0EC1L/r/tF2qZfdVU8grFeFGGImRIJeGEaIARmaH7/Ut53TRNSAbLbG09Zfio7Xma1bTexvj1TNN
7weGdNi/4Yl97A9EIo9LHNQ8Kf5qhr5qoUR6kAWBccqF+Fl+lOtjQyeo1/IrN0Q7gijvd+u8K31f
aYtgQUWadl+b6sYmrA8qp1I8GWOOQ/8HQEglCV85Wb5w/3z9RTRSx0N0fMaJ/XxN7a3o7Fn+Jtl7
EE0upxYMswenaXkiOO0t6Y1lPyTFtRrPWbAv2JtoJbZ5U1wC4z9kx+ZdeYZOQ0PZ7flp3zJsDwyd
0yBRfKVXq6/cTAgJnP29O+tTpKIHtZWOeAhSXvX6EzhEnAoOyImGmFMipJHFN/JEDJMxiwjiNM7k
k/rmUVuC5UKDm2QktZoDUE7B6HqDvtnvN1PTzYJ0dqv5cxvVUdpsFRRBIoo3M9V4z8kEXxZTChaN
idSAUcN/c6XnVxfLS2pczVUgIcWCFvFsmV36UytNn5wwlqlEnVia4C3mQQO7jBPvIWPQWWsb7Q3z
B+5JRzu7xKdW/k2gFsj2jOWYnTK+X9yhWWhNdkzmO2a5MYk9i+PbKSd4Tty1qt4WmB1EQF9ROTTM
9ayujlqBYYQoJEEv+LljIwyryPdQV4vYwWHaZlF7+RKZURj9eg8FxGSfFJwX6019yuNN0erLxL8M
8pLmXl+bMPV5tP17XfUMKQXswzMQ0Z2xwAbp6NGttdZGq3UxOeWubH69w4trOw0msdtZCxdkJIc+
cZVv06OmftcRujGcevpr9kzCJApOLwNauwZl1cOUFhZPau6/gwfmpSbNaqgKp+2Vob4o/0dJN3WE
GSHy7pWczHFQkekxviqVnWjusWIcjwojAbxfRVFLVl6pIPKrRgdNOpLa2K+1Nc2mAVJnPWk2ww+N
Vn+PG0w9bj6CaNwAS7sKt3vJzFSWlpa8mfzZZeEkEzmnh/n5VRC81GT2hMDx/5okYcx1ClgLCE5c
+8oqApwK/FTvfe8ONfb2wjNglPCHFxK46g9vl2FqqPiyemImWt7bITxd6hUqVzR5JeiV6BZoWrey
W71GceUIFiYRUWxHTsoH0IinKIDs8tX5C66sCAcw2rABCc+CfrOEkswn97l9gBFuOqWWCG8Pxsum
vFrHdUqiVXCRUyxIbFgSC2bBHVPogtAzMd34n0IEdZ0Mklt4fslYD6xbn8d6WqciACS9LSrAR5eG
ZQy7m/EUckhztIJhWiEqyYiMdDHqWO/Ubuib0CsvK7SkT8aaYS7Y1UAwj9pnzY0oIsnLTXi3hWnJ
hAGfYtastBv6HOvg9dpG7CABy6TB681QNxzYEoXwvE2tc7lmzaEB6UIO5xVo/rGJCNy+APFGbTPK
iWrnIq6SYlP1b5PMmdDhdsmvRwLDehYXcj3IIJ/WogR0hHrJlRRYxRhmzIyzZT7XaoD7+pR/zG3d
lsTMbEgU9jXzOyDh6jOLD1VnBgOqYN+2KI3ET6h3RBMILiKJiNQYepGiLvv9wrp4Dn6Tjr78mcf9
r+4MMbiZPpHvVIliucwCRrissp6l/F2NQQnLa80qzWZ4iD5AHSLu9z31pIxVOlZKn+ZGHmErtgNW
fIhbotE5dOWan+EV5Dv68MP15HHBs/3S5MNktiJbk+7vUtLdRHES9s3lX0fPLf5FhQFc+c4Odj3f
8tad/t+tMT+DPA8ftZuVPdtcraFUuG7Cc9y8mqutHI4YVW7R0tKd1kJTvsAL5mDR/QWNFRUC/IUW
FIeJHRbkbGzBJXaa31DtZBjzbn85ocKstRx4NZkskWjLWejrGkg86ufwTyDfDe3fpUpex+pGbcT0
p3GT46Nil/B1DVc9Q6AvpLZ/rK5mVir2lDykJnnfg8yx4IDdunwtCtnrVsf0KNVgC40ECCCQ20tM
YBTUiBBKYDcBWgY89fUjxdKGw0uYyO+e4T4E3Yq+hNHfNZVkEh2+BlX9Wv6Sf5GIr1VAC4n3gpZq
OxeTh8HWY0Ymp1tFkjuen5EeG8AOAX8FVbohUueTr1wTyRWhTUs+nxIsoRJcXv91naXDYRtdpr9y
Bl2Cq9BiaKFDGgVg9a9q4Ji8YpV+JYob3mKO+uQwwcte5o2KeoshXAM2Y2MypCFsgRB3oNEkT7/z
DbCLUfKGcFzqmZOLtyZidOb8ScONL4jBwMO5eQSkFP6D9tqVrT33OP4ZOJ6dENEG4BsUj4gA8Z1z
rpZUPsXPJ13V0fnnz+SlNL9eoTrHcdp6YZfFv/TBTGcjpKNaHAPwAyImCnH5nJFX9QjB6YXXGxnh
6L+pDw0Mr8Xrp8zuUPahvLaIqa676D0xe95TLY1byPoT2UZFCVRdaiyt1f2UgsWMHo/w5zmojujU
UKiuTlErUIBnc+YuTVEQSj+kSrBSd4oi0Xt2Dzb1yLcG7QZjCNmDFWM6vjg9tnpE2xjGpbpZParv
gO16h2dKJrxSjbehexktMoPYAOunJXgmr02DinzHvpSuSXBQx4Nu/qPDhE/VaGGJexIgQWDBut1a
noqE1/B+khIy2fPrAjy3uUez+ZIuERterjiZx9luzN8GS3ri2xxpF7HasagIq1kCfBK7G+H1XPLB
V13kIR7DU7O4PCKIITZxJbH94hhSjHToeZ8dIt4teC2Uv6k/X5IfWIaxPi2Go+cR6rmHiVx10Er7
lrnoWtADfWQ1vbCCEi1yD4U/eFprq9uP883zBfu7ht7arkzZEQWnuH8nHkwYEg29+O2oHIUUKx6p
rD1WPQRlD9PhorBMDARsa4Ay44j1cv2CCejP1pNzMFBTEagW7vDk6/BwO2YYfs7ZFJAWTLq4a0bd
3qwSV6SaHNGk/sXMMTpFZTFCQfuWctrNsngKnSQE2ch6TK/ay8c1v90iUfPoN1p/rRqR3Kt65kml
GuAUZlZyQhkYSnUGfRNgP7CuwFwPM3LC1fxnXxK3pQt5FtmZXEdw7gjlq1ILx7E1Qt1IjWE6bbBn
iQmgmVmhZyxdEQmFD2mSTm6hgiSPaWVfNvmm7kOYZbY2Wc8hvCFuaRF75KPKTgRkD2o5mvo1X5wF
nDiIw1tCVG5vtjStffqG5pGS7zI8XAoUfcjg28Moi7D6ooUYO92xaKSlzF2xw6DTS8o2gSCV2mhs
FT4s37AZTQxiquCPi/obJpHquFEbqtw0BV6yU93j+Cdf1XEkMu69Ewtr1ipg/Y9uGvuNr0/1q+ax
Aohn7lj5E8LqfBRBTMTe07aTBhLbgp4JTKr5RPrpE+qbHOBvNut6SmhVi75f/DhNeSTL/6ww494/
mRZP3c09vq70gLTNfCKKowWYfzE4bV4KpxhHma3jvi016wPhLD79D7PW3EnUnu6d4ahLsztPUVMu
QGP24+fVIHp3u94lqUfTnM4bVcPBX+6/yCyFEX3syPlt0WwTz08siKCM/pUOhZy+fKVIfiAqdWAF
kX6S5d7sdgprle8N72ZEeJTe0sNL+5ma54inw8m4GfLB1k5t2YywELdzvsUAXIcLjDTwJ7o73CQd
y2WJU2IXg7bDnmVHHA51PKf9FTfYVIGhBiA0RmBH9V/A6GGzIN5RQWcSo4MzGoxF3yjzov8g5hR4
r7FKRjoWB9SXIktMUmeS3pM1hfwoL48D65g8DTZkE6LBAfxmGxeJHslfCrZbc1AKtfkQoVr9Q0c4
orjGj61zdT/uFhOo/Zp3rSDOjyfnYtu+vnn8e1XRyoWBKf71ih+inGhIt3sn4yKk/IKF6qs70pek
H95AcfAnBFSYZkK5gPDKPd0IKiGFMph5oH/cKef/o1ueN8S1besQ9QnJOQ+QNfu7mt3IkvKYn61p
1JJ4tTXyhD3fN5oFP6dx7z7eqH5LmKa4z+t4kqCqBF10kXbaUNFY5hrCVHcoHa0+sKdMMXW3Sx0d
y8pBsBCsFNpMt54rJkmzkI01YWTdPys1Ov03QI/vl4w/13iPEv2D6OYssQidlWHnlNreUiJ7wZy5
ub1G+QFzWYzn6RTSWarq658CKzFQYq2YgyqClXfZVgoqgqIhRpIFnw29xxEPBg5wnD5/0beLy8JL
CGRrf8hq0Z3j3bp2ZDcdgqfos0x15E8rsd9Xqj+iSLrv+78UJc1VnRnr8/TwKV78nWxAFR8a+xHO
Yty2I9Nf5BwV3Eu2RqdCiMJrHakUlsCwf+IGC/SKBgTf0bvjD+RhqeQJfrB9deyZyaJ0Oir3WnFy
GdQuTqqWS8K76RWbXPg/DqNSrjKY2RT18UtolkTyjopqwdNoJPPOlXBi2cnE3IL41TBTfeNFGLBI
lcwiXCT8yK2IVfGWnNb/tHhO2/8o7eBkx5QxHllD7EWYTVySPurGmU+2k0OIFG5aCHKaldsBHCa8
/OTXU1z6xQuiP+FVVRBhpUhzixkut99T3aFaqbwNR7I/dQHrm85o3jrxxSz1otJ631rFbWc2mvbq
9a0usyf1/x9PnS9Ukwc+D60+vEvfsYPzCRvgY29hKa1ws8JWN2YOWfylTMYQgbGeq7lSPWWvnXPE
Mhk9Ex7Hs8CdzaLaRAxFsyzMCXLa7nWnwE8Yj2Rxq7i+kaygaO/nPU4w99HNkuvaIBxY0WD1dPqT
frTHL2Si8VsCGFJ2Pjo1iDLv3Zop/+WAo5Bj5YSBmL8yylX8zMELXnQfzJNowuMjbu1kHIgaN8BA
EnC3iOq3AAnTiXoshiDhWvmA5r+FT2R6Zl91Xh8cr0fReDS+l20m7qVy0XmIc1wzTjRcg1C9rKnE
ulR0i5JBRMl46tO52egJc53+Js6QOch7OOP2epY+zSG9x/0APGXLotCA1Cen0D4HXVXKOWvjDxft
J5VnpmtUNVvkTbLuHgoXtOSM4DkXO/I2tz9cEUJHyLeDsiqLkCNsVZeQygPdaW82+qGnsPQBbnCt
lLWH8Yskt85zPpyixI0oPQ59c9Ekw+/NDcEtuOEPuLA03smhxMUP2MBu7VZ1y7IJH8VNKwZozTwi
qgRTxNxJRMo6BnRVDF7dhqMLGMtSHOJszF9nr5TcjzjyOBP+rlOdQJ6NCSVQe3jTcBuSNfZ72fKu
ZZxi/a0BOtFhVyc2yskusZLIHejKxEA8dflmX3FCDrwmzeDDmmpxPUkWd1hIOYouGfa8KozHgmSR
l8H7DR9CuC7ujevaJ7/HqADTW2gkAtaaPYPrWDMcrgQSkzjrGgzmLgenj9HAasAuw3H07k5ZZ/gK
tiYNv9tYuBIqfWn3Eq7Q2L5HHb+/l18H+fE90lt+2IpWWjFI1xrx0lWhU8FvNw29Y3/Hgoq4jvV9
FAVWBrP6v7SFH+SRc7EX4y1hyMEFB44vDmhgJM9+qzffvCq1TEgZr/1O+c3hDtYsLf5do98v2LCA
YPPEui3JQZInhDl2LcWVTICe58gvLdnZWZH0339LADPae3pF/gfIfSGFnpmebQ8essDfteJwwAG2
+yo2v5piOoZU6m4IdLxvbw3o32z7uzP40Q/zMUcqT9FwxJLYVV/MqZUVw0DCe8tMAPWpleUxofcH
wiFlWtoYnuc4iaXHQOkWRmSTN0y9+14fcJSzoDaYWt6jpSNAIEgPn75CqBgyokA5G77p2OkYwJxz
VIdh3nT6mfXYd5jNnSVQS4q5iFbieVTwy38WTQSnegwc+xWc9QFDXYjfgkgEFp+VQ/7939SL+TDh
dFXMO/bDV/Gx5oUcRHtcHFUXLLb5LJO2hN1FQUZPZocJ+ydDrk4Dm/KhGEQk7iRboFqgHVO7fjrk
mDMV81ZHRELJx1nfvT/BJU/tObLns5jkWO+o6R4TXoChMe/pZcNmhS5mRznWTzuaQnpluH8t5X34
+4SuJ7tqpUPXo87z86CMKU3pZDg1OjRB612AHMVVyIQ8jaD5Ye2bleUpSqVTZXTWGL/gi499efTb
4VaGOZy3XOCV2adC+opcaBZnu1VxcBS3OgSU0XK+9zbgEpEfqECE9IT6n/HBcZNMkSpbSasZOmpq
LKvlqie6NhiL2g4ixS9rhz+6IDbzDblXGo67N5TjkAo30oI6eSgyXa02/idhzyocBFepmyTYApFk
N2JXzXzn+J7P4xD4z0ew3+Uj/4nUuPpvc9+O8bCWCU3ylqpaNcOC8PoXFUlisAnGCw5kvZxJ+JP2
12Dk4PCidFlus+3czZoYPC1Zia4CK7N8GuTb2H8rwURqCW1u8YjJl93QVEdL3oJwLuNrQYq/QYqZ
mgOQAPP5NvgmdAJMtMo1OE8MiW+gnSbRfmAU7G1z0V+zOcKcYFHtZBl1IP88eyar01y7R/76HR3Z
iuAJ7vbJMPFf97PrpPJOEipZ30k7eFGi85MFTM2L21b3iONwN1ARTMRF9xYuUoromHeFUU0DGU2g
MNaqFWWnO/7QrguDdAlFZR0q4kLonL/6WeznAEJk0ZZRXMy5pbCWLe7Xyh9azPA+QLXBexgfqB2a
URivdUJ6eeJZE4ldEN4tHwXmDmlEGO2UnRyqxzkoZbG2aHDVytsKhCSsHgQLzqR1Px3EkOGsimPm
BmsUQYzTGd88ngEjGBasMH9yO9Paz6rbJNBFB78nKbTHy/RnC8jYDKQQP/gsmgeyAHL3/pbgygX8
8CNO9OA42wsBy1cIwNaydzyLi1a4WRGRjAAS0wjU3ciKUwTx+qb9SsPv81VhW2GOpPgV+ILTG9t1
e4ydxWMM8fAJO8emlA50BzRI8IbwFr9hUG8EMJkZuDuv93TmfvkouadN5DJV1Yo61teyg9Fwc+Nx
gXFV8LqV9ZGQBPkMb4BHOe/qEdTUuNnrnMwc+0Hb5KrzwPsBJxPo64ok5+8Ds4IxX9vxigNvz8h8
MmdBtN9geMPSv/tr397ZNHwRr16MO6KXpL5f6Mk3WWyhX0TemZNvA9jnrCFgFkw2vR93wNWiKHWC
34WiTgAuZ30/k7alxmsWW4IdzlK4E1dN0Kb7nC1w9JiOvddvUGogRjIOVNzDEAMjEJ6XCzbZ3nCh
oQhyudILkMpG3gAkJvi5FKIbG0T8ag5H9mwkJ7Xs70g0voIzNmR7YYScm00QxDnInSTPLf4U7eDz
DAAWZWiShoj4wQw/GdPIVuH6jHvZd09L1/Awc0iF5ntnE8FwB4qbmkY24p/WtjRZfhIvBL333uVo
j/KqCa74hHonpdiT1+6fV9ziuLlsC076dwsTHCKMAp2ODbnyoS/drYRhG0I9KogvMQABsJqRQP9b
uJhqZR3LMWlu5l9FL0alo43vEMNMHsfp1FmO9QKIi8131u47Ojzsge0O0GjSpbqpupBmKN4ejyv5
7e6MeMbFxP65hZpeGTKajvRnw/v1QqalQdqNmoNLQA1z0L8sdzxeBvpmRfnRIK/1uRidMyMAmFJh
sv4PvjcznCsjm3MiR5QKeR9ov3NPf7DMLrUYEm02nHZCo+3WC+FTQ++YhtrU/MBCPqUeUex9VNZh
yZpoHdPZ2wlYutqREgs6dqW3AM5oqkdxjeLkvNefdpmtnsnM9PKAIcw8Nb6KWWhT0LSJvUE2m4dR
SiJn3YfdJO3QVCRKWD3yRkrNeNTDd4oVQ0lojt3zwj4ME4TilFyH8lE9UYRyZyM0rjEDbC/eD4HB
mocK1f8wneGt59BDS75sVhUKrnvuqGKDONepq+p8WgmPGoSd2Xi3qdhaAjwxZUmNVO0cOypD7hl4
hclPmjLE1ePxwu4dWnvtmtdG+RXeN/WDVF2WF7MqUARb+vkKjj5TAwdHyZtR1ZZdXUunhNTHOOL6
7AdTT7SPXWqfXTp7/bVubMYpqeWRQQlmxlcCw1ug0X8iv2LCMKyWQJK3Y/yEIh9ZCuaf9iSDxNWO
O7kTxh8loA7Bi9ZSGjotwxj4tZr0P0xC4JQlAgQWvy/vAy6hYKOxL2kdcDs2v5OhQNXxa+tO38Gv
RVI3BY2q0Dm6IUzMNHlx1xU+AAFvr/cZif5oHfzYqiS70ngGHe7myLR8kvoF2iOfanVf9gOHQIgC
FYgOkz0T258njmlwC5HgmeAor6UBlwBj2HEUptQSAT/ZB4xNn3quRdD2u/MQHGffX8QtP+WtsFVe
5E0QOsMp6eGvFpuQ1v2Gte68gTr1BKfOjThIpdlp6F4pWgBBlbTm2xf5yp6VD/Nf4sIjgjOfc04A
CU7Eg4/ALfwDSXiM+/R4d0Wf5FR/QsoyqtAeuFYMN240hLEzaT1BLy8dK8BTfGDw6M2Orl+yIL3m
RgLdb/hjobvfW2uVl9PWYdVMbcWRpnnp+Ylk6TL1fzZfPvSnIPSpLLTxVyxo0qMUfoklwySZC5Xd
bXUFLx4b5Qq5jogKt+cPIwktt7g05+SpF6IAo2M2W1as9ppOaSg9EMTmBZ9g0pVeMzqUSXCe7gHZ
6pVcYEDysdyCJnb6ubdBnWik0oCzr4klpkFOSSNJhRkYgK5U5NF9d55HgmJUSc+WaXoggWfNr3eu
MrePGHaeN6w8E0VOXo39mZ1ab8zTshrH/qvUF93GJxVlv7gklXGv1KO2DLNTOvVhnyXza3uRnZMq
CjRacalFvSsjjk1F6Ux8zt1KA9p8jIWNZIJvRkZ0qRvuAR++g+N52OCasPVWQnpI169KKBMpv0Jg
iHdOws31dga9/twh1opFTaKyvmsHVg1RDq5pea8M44ONsZBN22oDMqwSUFo8yZBx5xJmRHyPNb/Y
ymJC7QpQWY6XF8c4lofKdyvbVCOdKpG4HIw5FvgbY22i/3cZArItjM7r+LCffa8L3pu95oskA25E
90sCe8U/SpXgPdN7rljOtxYH2cjpXOhkeBEX1d2G1oXyHb/wvtySzCmiWIU4NKWnqrbCDOAw3pFt
al3V68ripVlrP0v1c9hFjIh3zwyUBtyjE6+5fJACfk0SFDcSx/cO9rejc73yy1s2+Kfdfpd4sX7u
ISM40ang8aNZmNBGnky1smeeScKVxd/toDoCvwDA6YmKs0jaICNmjExi4q74hiADfGMRdvQtrTzu
kYFeuG2fjAalJLCYZPygEI5MVzhMB3bKLONyONrVVpr+YtvFZwT8ZWw4L1vZ52a19+2LiOqkv6TS
VDAtipWCIPoNLTwZHXfYM/toLkkgBo6rgbd/cMkq+yhD+EEXcEKfEt9fd77hcTfVVqd4kNxcui+8
azVHDY8xfJcuwx5wYh5YTUFy2xTNL9Q/yFDmwdIoGIT4yl3WflAjrqUsuKvl/H252Gpn+M2bFT1+
jDckA14r4OaYNOZoDJ7JWQR58T9Y2ck+Fu68/B3gbVX6qWqvDLzTaOYmn2nSDINodA7Oni/9lDNb
SU8Egi1h+KuDXY1LqjRFZqUqaicc+N4u/ML3+9pJo8Z2GZn3a0Fac4oNRxZmEru9CjQzRywAMRj7
CG/CRerD8JgkSBoCJFPYoxEGVS89NV2Uo42CSj+IhGOgmNRWkwt/QJSsdVIsXTiCOoy9nzfE3m4Z
MGJJLnmx66GFDR6/A4KdoCMoe/leMIkByPnOdJ1z2BL7yauMVZyWA1r3wzynVRCiy6A9Sw5GRT+x
oBOiL+v1tituKo1IUJyOaacyeN//s8K4CJ9poFlQYRTK2Tw89NitTtikgcesvZQaoYy2lnEjhwQS
8rnIq0fzwfPqh2Jy8Ey57j5eqgCCa0sdqg54Gi9YO7tfsaAS3g/Ywc/1vG/EIJHcOTZXO6kKZz9r
AzcztIUBYZNar9VJkwb4AUD5hy9mpsppJ6WlPbnkvBXHu3kgwd6j4o9BDkl1PsRd+4bjPdX0ivBJ
vYpeZPWgC0zjSSGTUtWnGSE2Zh/hl3NbDKZkPq/Kx75kKjVDWQNQZxlQY7r4489EQEFmZUPbjlMQ
027PBQDZoPHCUW6lJZjZ8pL1fKJ25CeLrksy1skHsrn/5+xyqhCD6QxQQeGhjXz2kgteaMOPiqiI
ww12o/Zk/JGuIUKX4F5HUT3sMbJVuqeHrAQpZJJp9lzP6R9n/jmXIUBEqipKc9Am4jbNHdG+KEGX
wFHuV2tamgVX8Oe5RW40mNxh9NC+BLS1Im75yq55i52kQbJAtm6sbp4Mw2A6e3Y/3dMRVihhAETS
Ray1jdTJyRc8FlZBhba99bpJACBZkFi/C/pMDfXQA7nTJOpS5tOE4LqJwPX/Tds+FnkE5gSft6Kf
r4YX9GnhHhjQBNS3TR0bmrzLXmMQP93dyabzMLwYt9fXPvG4zCOsqtD2wElzvMK8jMJ4NA9iuxsF
K4dzXhu46VCrEB6hGa31Jc2ADuy209J/KicY7EPnaItua5cdK50JPTf1mNSGrIfimRWGZ/O83DbF
ezcX9mefxGtEq5jkxd5lKvcKOl0am2EK5I6O1gSnt5akXDjGF0HO4Y/P+TVpwmKz8wVUwDHaelAq
1z9ys4qKFXAbwriGx/XFXURhvlmEl4o9XLXpUQCndLaL8PWmsenPE+m7JqZJ5D4idvSSwOcTylgK
KBwzjlQuRUqMwlnsAMq0nUXRIH9QYTRQ6l8tVGlp4n5lhYRXPNC/gREFcc4HWE8GuOnO8qgTpgZu
6+pAPWG3ZpGrlvoDUd97pdWNVsxkvOGm/4jtMbDrNq/x4jRISsyNqi6hFPoKWm32VC6prFoc1iaS
2t9qlc6okDociTlysgzomTq1CEXBSxAG7N6YGqiwzqWShownPnCQmjXr/H6WzGWxl4jv2p+MnDPE
PU/9G7LKVajRmybS0FZWq3e1yAFNPjLHxDIwlxP2dX2C90uSaQcYMVzsqQsr7e/aoHNkoQRKlxhx
EFWg+DiPtau3g5ivFP4U7gr6DVBJoqXXlmhlc2r84JJcheYBqPpXNlP/BO18lkOeatSVYbHEZxvM
X4V3XRCMHs7M8+F7Hfv1k7kajjz7jl2xq0NfAweQyd7FcSUkn46YSMnuqU/IfiSlsMfYO9SM9bjj
cLLVWgbiT7A5J2nX0d0mCMrO/UNJd0qd7FORW8X9blQVemVpc0V7iajcs0ppXczsFd4je228OZQa
Zq2wbQWqwVFayGuWEwBTqTHZvEx+O6WZgQSX1RUTU3Y3xLOnVDlY8WIeovp/MjSUHOmnyFS7U0rR
tVsCOurC6YqFDEGKnAxIpYjwFoK4c7ISvcS1HnbRpBEMexpzX/9xIeouSjwymZcd77kBhODiGQz1
NPZmVGdKzbidGfQsWwVt02kSXvNBXa/1tMe5UOGYNCLSq0l5Sbm+zmrD+jLGCGtuvmNCDt48dOC6
gZ5OB3GhHESJgCk5m8JH+eTDwXY5ZtemZeSjrCp2fNxsufJAL0GXW1Kv4ui3jz2jsnmq5boEzqyr
l9ly7xLNKWqHLI5HOtTyXvOijxPjwohIUtNMXs88macYDwhpKZZVMW4xmadHLIfFAr3kUOz39Gcg
eDZ6eDzM4IhFNkuQ6oUvav/ZlCEqRpTrMxH/Ron90jXdk40N+hf1f/o00X0hyy/LexxKSmlDe7M0
t/yjXUYO2Rp+yEwmepkBEm35PCmPXQ29VWaagJQ3sc7s/SgLy0BaIIKMFLq7Hb1dNgfjIDaji/Yl
20rGqJnm3f9vioEHdCJ1mfTKRIfiT3wKyJCmm8Czjxh4nngoaaJWg6ImFScO6PrZrt0KQyk8A5kv
DQaZtnpNeGBwA74qjTJbhS9Llgp+76gY3NzZXvm2O0uRMyOp/w+JbuypDaWg7mWvJBSl5M7Ygkdu
VF53dOm39YPcnEKj5+wUypzNMbf6Ri2fYiIQwGNosEUFbR1sG7vdPPDim1SbW4AcfYAfXwyY54UH
LoidxwyrtenIZNK4N6apWlo5+wo93wm+HalibMZzYG64jQ6ES5sanViplWhaMpP4SGBnZvTqZFTM
BUWGRRtJeNU2icjfJH8NVv3B/9rexM33csjNq1yqbdMgdEem1ReJ1ATVQks8wBN+p0fondu1/rpx
UdHEwWR/+ud9r1L1Dc88XkyAIkbzMcUFLVYVgn2GNXLaK8vCAIt5O9pC5J3yIGCU8Z7T25SwsvXG
uPSuso9XYHRe1tZA1EWxtUSZW3LFGFWA4uy1SMBeBah8a+tRPwZHjCllAfHyk9tOrz1YxIMTSR/6
aTEHl8lCTERnBmBLbWF9biDDUFR3+lShIEnnmj4u9kp6VRpj2r8qldO6/pdL/oEdwA/f5chLU2To
32yGQBUYloJOrdpgbB526Keob0BmJY2m3V+vwIb9c7kFeKn0umCAjcB2ZgVZ8aIl8BCstTIeT0Y/
kqLpUnBqucvlhBUgiaK+Y+vojb30mEUCtWWDrLkWQg1UUzPcODmemdJcD6Q1EjQeKuR/5IBw0fTl
jnzpZe34KC1m0gyhb9ThJQ7GM9JeRX544Wl/VQzUxA9j97/GHHSV4QtPk/8p86jhKyqN62puI1KM
yoEEWOx5XoK2TogYD9dAXixsIe/iU2Ecjm/1xlPoZLIOsa9rnpbyut1TG7HLOiTo8gkYImQHTKmc
P6wu3axhb5UyT00ONAwYyPFF29zWtQC2E9nc1Uox5TkhhhL4oU/UZOhuxptLNUli41FCt41P3/d/
i13RjKR853qVssC1lN0qaWTQWqnz4a62JeXQZe2XgtbXt9+m0gBEJBl3xs/xJiry4EwiIHKSOEZO
jOemBLtwIQNN1LTt7boExxCYwMfvjDTkX6BENchjcveutY07yvLrj0f8get0MiOJ2sYZQkNPcnaL
adsBODH2AIxttjD27nPr9bc6acsv/mhOz3yuzRBEDQFQP9y94NOhjR+LrgedbmJh3zTHj60X0e3i
dA/eJFyC9wlZ5l6t6ugZVuF+dQBrEaZN0gwyLiO+/zuJmD7p/d0zMXZz6HskBMh9rEn86edJb4PH
TN4M0eEL1EmUL/SzAWaRjThirDFG/MaxKirHGioLM925j0G8Xg1W8/iahseGLN3iWFCibWx6c7De
+V84f+cxsVrkDYt2+mk0JtMpaVFaA/KD6ciVXVmIM4s3aroljKrmUG8xT2JngU5J2ST/mdvlHH8a
VpqhRSwW+trMQiA0OdQWGPAuMmj2jJo/5s/nmddpbxPogDAa1E6x+x5MJzjm4ZeX793bxMO/BSoT
ZooGjbt18U3QHF7Fcm8R0RS6oTSJj7Imn9e4FCLAG+NoEQX+ovpDfU2sZ0K4Ao4VUOV7fLtIZORI
JZX1rIblKTqopPxt7btpwE1budDyCYMnnNXtltsYdNHmcUUslpSDi1AlcgXfm6uOHImZhDlEm0WS
+aYnBsq+byDQVYH+ImxGbVCj5gz0e7j8tT01XEL7j4BiUpm4FC8yT+AfAbQphhA7wR+4mxeYAihj
vPUgaqIN/81m2bvKpl/00vdaLSUyH4/TcwBYdxYR+6QQUUgLU/8fJsUdAHRTlmHmoyc75NyC06C0
XZCiHSa4T0F3ndHC40BqUhr89jTQ8QcEK0/EMiEs6n31yYe/EWaFyYYlTVlXD+cBZcxe3scDaHLc
achmVor4s7ezkDqVctzNFGegluqmDcccnHtLfHTQQBXPjGsJp3ASlkB4VLcZwJuKS5AO5nN9/nJA
DvIRH4+gXrr73fcsxK5Z2x08+ZYK5R07d/ZgRGOEa7eqT+uUSY7YRUIWwOQUgtb0FBhy3JOuIAak
hsdnO3ZYD1q94trWxPDfjJvDCVXADQM/4VSfKcecFM5tHbtQ5MzY6HuSyD9KRIvT7Ous8pQC5quq
Lt+OMgNWyIOj4dNv7DD2HMGkJoyIryF0UyPXQPzF/a9jZY1coeLHURoTDUWTYogVTysHE7wtNkre
aXNqsn3XaZ017TBYJ7kqvLqlsvpd35MvrE9cHbJrjcKM2l5ensq6GhpLM8nXM0WbIIoFH08+VZnY
2EK8HRjnhAg+oUxH9nQD+x92gfLL8ZoDsFj3I7R8pyGZRKFJ0U03mTATEnUI1RLZwfxi1RP3HFW3
mY1vokkw98CQNBQitjiQBxBszjQ75DUFXSLgtQ/sulwvCCUHDQCbPL6eV5V+2Yh5oUiRYIsFjxWn
G3opgSUvJtgcPsv89XVB9ed5mHLHhD9mUzO4x3AU1UBP2SJSRHQvhFZWq7zcurKx4f4erDTTOkxZ
axLXw+a1/O1fFmTp4zW4rjl8ZVv6b8p2RsJGMVosVebIdP+ueR/xi7r9i6QPDMoClDYsTyq55ElX
ypFk4ui49MzUmUd+xtO/CeWblVSCy7qyhKpZUVdq7pT1e7fN3Xs4u055U2kB1igHjtN705HiPSAa
xmDgYSMOUxAk6wPbN7w4m/lFfdbZZVUYPVHVWcPftv2dPZXMLaecn2oex0P8YlY3KsGUrtgfskPU
0xslDxnsrqb+SbFX1YVjvF/GU5UpmsydI9Huj43rXhIo95R5H6rvOIdgOlwoMQjGw+CerBZ0Nccc
JpIxsO3iEx7MnYkCra89dW2U3St/SPd2cpdlg8D7I6bW98zxZZtMTt2BSQHWl1wEAKwXTIYdwG4Z
gQ+9VMyVElO8CJbNs5PgvizoUL1qwrdFHw2HGQPC8Kf3bslUIYIY0UcpnKHRypnkb4RIUB64uP6s
q/WXt+NmNtAdkhLMrLzHM/OAD6R+Wweg10z+C3a9PYg0N/5WEyZ2cSl2QeH5hdFXV+xTuxaiNtUk
Ml46zREPqdxla3h8n7OMpj5nknJH4t4X4E/SQt3w8U7UQXswgpDcIRBpe1tbMwdmRxZoFPWn6gLz
i9Tk+aYQbQQmLIHv6a9hrkQA1oOU48TZ1bYnyjw02iSU3GtHBmacl4GnxHaVwSUQeI9oEvMKbKTr
gTBo0WGuzQ67JUfrlO+kQg6cAnZK9sxvCKfIQ6vBCLKFa2yzcPu3u7r/WCmhD1hpzcAzGHvCsvFG
OayOwHgR+Op0mj4BI4ijngdcFVdgBTB+acxUYVEdD/HQzaiuYO3wAkknAuHVi+8VqoeYiznGddnR
BTJgGC+SOYzPm7sVbDxdjoTg2NJYCOpf7qz7ZNUActopukXuRW4dpLXyqlmcqosmuFcFthVd6GMi
pTLzEdpSzbMcNNVfRm1s9jTTtHfreTu5vBLcuny9Q05y4tIl5bjdJeN0Q5ZCbn9w6UuqqNWFUWlz
1gkZrSF1P41zjyijLsYNxvLNMlJihDxYHRZ6tmqDrDnmRQ3FIZD7QX/vZE+VNA0GCrzE+FRbYbKq
lCMkBb03+HhsZx7LhoS3AjrhHYkB7ZB9fRgrtNcRyDj+BJnVCKQJb9Y8WiP4pC6TtcX7pugZNUIl
ZYMtZXNOfNzrU3Gsq5nc08D9pLKrXRSqSytOmil4WgqfpFY9kCx9Ef1EWAlf80Vr5yIvZL4o9+GG
9k3Q/ZlDd4MEuGyA14gsOpMQY7optG5ni6Qg6YTpAECOY+N00A0C0/PV3JC6cuhonanoN2F5qEDR
JRoOTSEN/3GALtqZGHS4NoY9YJxMqjb58ZQjeIvZPmEhBdWQsTBND4KSriG6Gs0bY5UnJW4jq7+4
Uov65AZZSr60CTkOwilD4bCLKyV/HDp49TdKJNqnTzg5YihWcA1JNb7EIBUTtqsS81OCxYxQtKzY
Ix6m0QkLxyFAzIEHvK/tewzLX4L83nYwfYmSVCqhp6iDZ6yzmidsljlPecXbXs2gj7+tZLPbt6lY
ihOf85d0z/h1j+T4comIOOEDJwHYzv4hah3pWUV8q6Y1Y2upCUoPGOUaiO+tCjSnsVzvrpIAR/s8
6akS5oxkC8Sp8tO0pXKXZPDv28wkeWlkk7DaWU4S/YGA7E1EoLg3MagJp4sS2laDMU3Nbz19im3w
7cAZR6Xu28TdEKVXpcL8nsfm+QqzZd13+i6IoF2Tezy2OeucVGZjLQIPDtcKwya/TkPsJUWKAOH0
OQXPZPLEyGjjpIwah7tyeJiKx36lvDPlfctOp0ssADgJcQu6PSrZjCKsnCINEvqxTBYENn1rDJWO
Z0mH3IsXeFKOp35uhW7FlqA8iLvt2o+OpvFAK0Qlw2loT9cLY1DU+/Cu2lT6xlyjkWzmA7w5mPNL
XgmH4nWekgl2xaoieckFKhnid69HG/dgL/gPu+44O0K/iI0gH2uMNCUvGdXb38yOtK6ibzzAUHB7
gFrTpwfcMQxFgM0P/POJAIlv3oX1WVbe5cRpcmVPioflGQ/CBHXQs98UKdHG5QYxSTNYhPMtvhVo
S//EKQHYc6nqyYAjrvRWHMldWTaF9FyF4dcdGXDxwy/p+IEdvUqPjF4OoLV9sTqRhtVCwf6XXROy
lMTYF2mIsTA+9gIPkTzM1ZQA7ithU5F+wuvw9NDA6crZIIVMDtuWp7Y7beCzRuyUYnYIgr3t1yCx
y0WuEy71dRne/UQBZbjzzXxLg6GSfA==
`pragma protect end_protected

// 
