// Copyright (C) 2022, Advanced Micro Devices, Inc. All rights reserved.
// SPDX-License-Identifier: MIT
// ==============================================================
// Version: 2022.1.0
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module testEnc_process_r (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        p_read,
        p_read1,
        p_read2,
        p_read3,
        p_read4,
        p_read5,
        p_read6,
        p_read7,
        p_read8,
        p_read9,
        p_read10,
        p_read11,
        p_read12,
        plaintext,
        ap_return
);

parameter    ap_ST_fsm_pp0_stage0 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [127:0] p_read;
input  [127:0] p_read1;
input  [127:0] p_read2;
input  [127:0] p_read3;
input  [127:0] p_read4;
input  [127:0] p_read5;
input  [127:0] p_read6;
input  [127:0] p_read7;
input  [127:0] p_read8;
input  [127:0] p_read9;
input  [127:0] p_read10;
input  [127:0] p_read11;
input  [127:0] p_read12;
input  [127:0] plaintext;
output  [127:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;

(* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg    ap_enable_reg_pp0_iter5;
reg    ap_enable_reg_pp0_iter6;
reg    ap_enable_reg_pp0_iter7;
reg    ap_enable_reg_pp0_iter8;
reg    ap_enable_reg_pp0_iter9;
reg    ap_enable_reg_pp0_iter10;
reg    ap_enable_reg_pp0_iter11;
reg    ap_enable_reg_pp0_iter12;
reg    ap_enable_reg_pp0_iter13;
reg    ap_enable_reg_pp0_iter14;
reg    ap_enable_reg_pp0_iter15;
reg    ap_enable_reg_pp0_iter16;
reg    ap_enable_reg_pp0_iter17;
reg    ap_enable_reg_pp0_iter18;
reg    ap_enable_reg_pp0_iter19;
reg    ap_enable_reg_pp0_iter20;
reg    ap_enable_reg_pp0_iter21;
reg    ap_enable_reg_pp0_iter22;
reg    ap_enable_reg_pp0_iter23;
reg    ap_idle_pp0;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_state4_pp0_stage0_iter3;
wire    ap_block_state5_pp0_stage0_iter4;
wire    ap_block_state6_pp0_stage0_iter5;
wire    ap_block_state7_pp0_stage0_iter6;
wire    ap_block_state8_pp0_stage0_iter7;
wire    ap_block_state9_pp0_stage0_iter8;
wire    ap_block_state10_pp0_stage0_iter9;
wire    ap_block_state11_pp0_stage0_iter10;
wire    ap_block_state12_pp0_stage0_iter11;
wire    ap_block_state13_pp0_stage0_iter12;
wire    ap_block_state14_pp0_stage0_iter13;
wire    ap_block_state15_pp0_stage0_iter14;
wire    ap_block_state16_pp0_stage0_iter15;
wire    ap_block_state17_pp0_stage0_iter16;
wire    ap_block_state18_pp0_stage0_iter17;
wire    ap_block_state19_pp0_stage0_iter18;
wire    ap_block_state20_pp0_stage0_iter19;
wire    ap_block_state21_pp0_stage0_iter20;
wire    ap_block_state22_pp0_stage0_iter21;
wire    ap_block_state23_pp0_stage0_iter22;
wire    ap_block_state24_pp0_stage0_iter23;
wire    ap_block_pp0_stage0_subdone;
wire   [7:0] cipher_0_ssbox_address0;
reg    cipher_0_ssbox_ce0;
wire   [7:0] cipher_0_ssbox_q0;
wire   [7:0] cipher_0_ssbox_address1;
reg    cipher_0_ssbox_ce1;
wire   [7:0] cipher_0_ssbox_q1;
wire   [7:0] cipher_0_ssbox_address2;
reg    cipher_0_ssbox_ce2;
wire   [7:0] cipher_0_ssbox_q2;
wire   [7:0] cipher_0_ssbox_address3;
reg    cipher_0_ssbox_ce3;
wire   [7:0] cipher_0_ssbox_q3;
wire   [7:0] cipher_0_ssbox_address4;
reg    cipher_0_ssbox_ce4;
wire   [7:0] cipher_0_ssbox_q4;
wire   [7:0] cipher_0_ssbox_address5;
reg    cipher_0_ssbox_ce5;
wire   [7:0] cipher_0_ssbox_q5;
wire   [7:0] cipher_0_ssbox_address6;
reg    cipher_0_ssbox_ce6;
wire   [7:0] cipher_0_ssbox_q6;
wire   [7:0] cipher_0_ssbox_address7;
reg    cipher_0_ssbox_ce7;
wire   [7:0] cipher_0_ssbox_q7;
wire   [7:0] cipher_0_ssbox_address8;
reg    cipher_0_ssbox_ce8;
wire   [7:0] cipher_0_ssbox_q8;
wire   [7:0] cipher_0_ssbox_address9;
reg    cipher_0_ssbox_ce9;
wire   [7:0] cipher_0_ssbox_q9;
wire   [7:0] cipher_0_ssbox_address10;
reg    cipher_0_ssbox_ce10;
wire   [7:0] cipher_0_ssbox_q10;
wire   [7:0] cipher_0_ssbox_address11;
reg    cipher_0_ssbox_ce11;
wire   [7:0] cipher_0_ssbox_q11;
wire   [7:0] cipher_0_ssbox_address12;
reg    cipher_0_ssbox_ce12;
wire   [7:0] cipher_0_ssbox_q12;
wire   [7:0] cipher_0_ssbox_address13;
reg    cipher_0_ssbox_ce13;
wire   [7:0] cipher_0_ssbox_q13;
wire   [7:0] cipher_0_ssbox_address14;
reg    cipher_0_ssbox_ce14;
wire   [7:0] cipher_0_ssbox_q14;
wire   [7:0] cipher_0_ssbox_address15;
reg    cipher_0_ssbox_ce15;
wire   [7:0] cipher_0_ssbox_q15;
wire   [7:0] cipher_0_ssbox_address16;
reg    cipher_0_ssbox_ce16;
wire   [7:0] cipher_0_ssbox_q16;
wire   [7:0] cipher_0_ssbox_address17;
reg    cipher_0_ssbox_ce17;
wire   [7:0] cipher_0_ssbox_q17;
wire   [7:0] cipher_0_ssbox_address18;
reg    cipher_0_ssbox_ce18;
wire   [7:0] cipher_0_ssbox_q18;
wire   [7:0] cipher_0_ssbox_address19;
reg    cipher_0_ssbox_ce19;
wire   [7:0] cipher_0_ssbox_q19;
wire   [7:0] cipher_0_ssbox_address20;
reg    cipher_0_ssbox_ce20;
wire   [7:0] cipher_0_ssbox_q20;
wire   [7:0] cipher_0_ssbox_address21;
reg    cipher_0_ssbox_ce21;
wire   [7:0] cipher_0_ssbox_q21;
wire   [7:0] cipher_0_ssbox_address22;
reg    cipher_0_ssbox_ce22;
wire   [7:0] cipher_0_ssbox_q22;
wire   [7:0] cipher_0_ssbox_address23;
reg    cipher_0_ssbox_ce23;
wire   [7:0] cipher_0_ssbox_q23;
wire   [7:0] cipher_0_ssbox_address24;
reg    cipher_0_ssbox_ce24;
wire   [7:0] cipher_0_ssbox_q24;
wire   [7:0] cipher_0_ssbox_address25;
reg    cipher_0_ssbox_ce25;
wire   [7:0] cipher_0_ssbox_q25;
wire   [7:0] cipher_0_ssbox_address26;
reg    cipher_0_ssbox_ce26;
wire   [7:0] cipher_0_ssbox_q26;
wire   [7:0] cipher_0_ssbox_address27;
reg    cipher_0_ssbox_ce27;
wire   [7:0] cipher_0_ssbox_q27;
wire   [7:0] cipher_0_ssbox_address28;
reg    cipher_0_ssbox_ce28;
wire   [7:0] cipher_0_ssbox_q28;
wire   [7:0] cipher_0_ssbox_address29;
reg    cipher_0_ssbox_ce29;
wire   [7:0] cipher_0_ssbox_q29;
wire   [7:0] cipher_0_ssbox_address30;
reg    cipher_0_ssbox_ce30;
wire   [7:0] cipher_0_ssbox_q30;
wire   [7:0] cipher_0_ssbox_address31;
reg    cipher_0_ssbox_ce31;
wire   [7:0] cipher_0_ssbox_q31;
wire   [7:0] cipher_0_ssbox_address32;
reg    cipher_0_ssbox_ce32;
wire   [7:0] cipher_0_ssbox_q32;
wire   [7:0] cipher_0_ssbox_address33;
reg    cipher_0_ssbox_ce33;
wire   [7:0] cipher_0_ssbox_q33;
wire   [7:0] cipher_0_ssbox_address34;
reg    cipher_0_ssbox_ce34;
wire   [7:0] cipher_0_ssbox_q34;
wire   [7:0] cipher_0_ssbox_address35;
reg    cipher_0_ssbox_ce35;
wire   [7:0] cipher_0_ssbox_q35;
wire   [7:0] cipher_0_ssbox_address36;
reg    cipher_0_ssbox_ce36;
wire   [7:0] cipher_0_ssbox_q36;
wire   [7:0] cipher_0_ssbox_address37;
reg    cipher_0_ssbox_ce37;
wire   [7:0] cipher_0_ssbox_q37;
wire   [7:0] cipher_0_ssbox_address38;
reg    cipher_0_ssbox_ce38;
wire   [7:0] cipher_0_ssbox_q38;
wire   [7:0] cipher_0_ssbox_address39;
reg    cipher_0_ssbox_ce39;
wire   [7:0] cipher_0_ssbox_q39;
wire   [7:0] cipher_0_ssbox_address40;
reg    cipher_0_ssbox_ce40;
wire   [7:0] cipher_0_ssbox_q40;
wire   [7:0] cipher_0_ssbox_address41;
reg    cipher_0_ssbox_ce41;
wire   [7:0] cipher_0_ssbox_q41;
wire   [7:0] cipher_0_ssbox_address42;
reg    cipher_0_ssbox_ce42;
wire   [7:0] cipher_0_ssbox_q42;
wire   [7:0] cipher_0_ssbox_address43;
reg    cipher_0_ssbox_ce43;
wire   [7:0] cipher_0_ssbox_q43;
wire   [7:0] cipher_0_ssbox_address44;
reg    cipher_0_ssbox_ce44;
wire   [7:0] cipher_0_ssbox_q44;
wire   [7:0] cipher_0_ssbox_address45;
reg    cipher_0_ssbox_ce45;
wire   [7:0] cipher_0_ssbox_q45;
wire   [7:0] cipher_0_ssbox_address46;
reg    cipher_0_ssbox_ce46;
wire   [7:0] cipher_0_ssbox_q46;
wire   [7:0] cipher_0_ssbox_address47;
reg    cipher_0_ssbox_ce47;
wire   [7:0] cipher_0_ssbox_q47;
wire   [7:0] cipher_0_ssbox_address48;
reg    cipher_0_ssbox_ce48;
wire   [7:0] cipher_0_ssbox_q48;
wire   [7:0] cipher_0_ssbox_address49;
reg    cipher_0_ssbox_ce49;
wire   [7:0] cipher_0_ssbox_q49;
wire   [7:0] cipher_0_ssbox_address50;
reg    cipher_0_ssbox_ce50;
wire   [7:0] cipher_0_ssbox_q50;
wire   [7:0] cipher_0_ssbox_address51;
reg    cipher_0_ssbox_ce51;
wire   [7:0] cipher_0_ssbox_q51;
wire   [7:0] cipher_0_ssbox_address52;
reg    cipher_0_ssbox_ce52;
wire   [7:0] cipher_0_ssbox_q52;
wire   [7:0] cipher_0_ssbox_address53;
reg    cipher_0_ssbox_ce53;
wire   [7:0] cipher_0_ssbox_q53;
wire   [7:0] cipher_0_ssbox_address54;
reg    cipher_0_ssbox_ce54;
wire   [7:0] cipher_0_ssbox_q54;
wire   [7:0] cipher_0_ssbox_address55;
reg    cipher_0_ssbox_ce55;
wire   [7:0] cipher_0_ssbox_q55;
wire   [7:0] cipher_0_ssbox_address56;
reg    cipher_0_ssbox_ce56;
wire   [7:0] cipher_0_ssbox_q56;
wire   [7:0] cipher_0_ssbox_address57;
reg    cipher_0_ssbox_ce57;
wire   [7:0] cipher_0_ssbox_q57;
wire   [7:0] cipher_0_ssbox_address58;
reg    cipher_0_ssbox_ce58;
wire   [7:0] cipher_0_ssbox_q58;
wire   [7:0] cipher_0_ssbox_address59;
reg    cipher_0_ssbox_ce59;
wire   [7:0] cipher_0_ssbox_q59;
wire   [7:0] cipher_0_ssbox_address60;
reg    cipher_0_ssbox_ce60;
wire   [7:0] cipher_0_ssbox_q60;
wire   [7:0] cipher_0_ssbox_address61;
reg    cipher_0_ssbox_ce61;
wire   [7:0] cipher_0_ssbox_q61;
wire   [7:0] cipher_0_ssbox_address62;
reg    cipher_0_ssbox_ce62;
wire   [7:0] cipher_0_ssbox_q62;
wire   [7:0] cipher_0_ssbox_address63;
reg    cipher_0_ssbox_ce63;
wire   [7:0] cipher_0_ssbox_q63;
wire   [7:0] cipher_0_ssbox_address64;
reg    cipher_0_ssbox_ce64;
wire   [7:0] cipher_0_ssbox_q64;
wire   [7:0] cipher_0_ssbox_address65;
reg    cipher_0_ssbox_ce65;
wire   [7:0] cipher_0_ssbox_q65;
wire   [7:0] cipher_0_ssbox_address66;
reg    cipher_0_ssbox_ce66;
wire   [7:0] cipher_0_ssbox_q66;
wire   [7:0] cipher_0_ssbox_address67;
reg    cipher_0_ssbox_ce67;
wire   [7:0] cipher_0_ssbox_q67;
wire   [7:0] cipher_0_ssbox_address68;
reg    cipher_0_ssbox_ce68;
wire   [7:0] cipher_0_ssbox_q68;
wire   [7:0] cipher_0_ssbox_address69;
reg    cipher_0_ssbox_ce69;
wire   [7:0] cipher_0_ssbox_q69;
wire   [7:0] cipher_0_ssbox_address70;
reg    cipher_0_ssbox_ce70;
wire   [7:0] cipher_0_ssbox_q70;
wire   [7:0] cipher_0_ssbox_address71;
reg    cipher_0_ssbox_ce71;
wire   [7:0] cipher_0_ssbox_q71;
wire   [7:0] cipher_0_ssbox_address72;
reg    cipher_0_ssbox_ce72;
wire   [7:0] cipher_0_ssbox_q72;
wire   [7:0] cipher_0_ssbox_address73;
reg    cipher_0_ssbox_ce73;
wire   [7:0] cipher_0_ssbox_q73;
wire   [7:0] cipher_0_ssbox_address74;
reg    cipher_0_ssbox_ce74;
wire   [7:0] cipher_0_ssbox_q74;
wire   [7:0] cipher_0_ssbox_address75;
reg    cipher_0_ssbox_ce75;
wire   [7:0] cipher_0_ssbox_q75;
wire   [7:0] cipher_0_ssbox_address76;
reg    cipher_0_ssbox_ce76;
wire   [7:0] cipher_0_ssbox_q76;
wire   [7:0] cipher_0_ssbox_address77;
reg    cipher_0_ssbox_ce77;
wire   [7:0] cipher_0_ssbox_q77;
wire   [7:0] cipher_0_ssbox_address78;
reg    cipher_0_ssbox_ce78;
wire   [7:0] cipher_0_ssbox_q78;
wire   [7:0] cipher_0_ssbox_address79;
reg    cipher_0_ssbox_ce79;
wire   [7:0] cipher_0_ssbox_q79;
wire   [7:0] cipher_0_ssbox_address80;
reg    cipher_0_ssbox_ce80;
wire   [7:0] cipher_0_ssbox_q80;
wire   [7:0] cipher_0_ssbox_address81;
reg    cipher_0_ssbox_ce81;
wire   [7:0] cipher_0_ssbox_q81;
wire   [7:0] cipher_0_ssbox_address82;
reg    cipher_0_ssbox_ce82;
wire   [7:0] cipher_0_ssbox_q82;
wire   [7:0] cipher_0_ssbox_address83;
reg    cipher_0_ssbox_ce83;
wire   [7:0] cipher_0_ssbox_q83;
wire   [7:0] cipher_0_ssbox_address84;
reg    cipher_0_ssbox_ce84;
wire   [7:0] cipher_0_ssbox_q84;
wire   [7:0] cipher_0_ssbox_address85;
reg    cipher_0_ssbox_ce85;
wire   [7:0] cipher_0_ssbox_q85;
wire   [7:0] cipher_0_ssbox_address86;
reg    cipher_0_ssbox_ce86;
wire   [7:0] cipher_0_ssbox_q86;
wire   [7:0] cipher_0_ssbox_address87;
reg    cipher_0_ssbox_ce87;
wire   [7:0] cipher_0_ssbox_q87;
wire   [7:0] cipher_0_ssbox_address88;
reg    cipher_0_ssbox_ce88;
wire   [7:0] cipher_0_ssbox_q88;
wire   [7:0] cipher_0_ssbox_address89;
reg    cipher_0_ssbox_ce89;
wire   [7:0] cipher_0_ssbox_q89;
wire   [7:0] cipher_0_ssbox_address90;
reg    cipher_0_ssbox_ce90;
wire   [7:0] cipher_0_ssbox_q90;
wire   [7:0] cipher_0_ssbox_address91;
reg    cipher_0_ssbox_ce91;
wire   [7:0] cipher_0_ssbox_q91;
wire   [7:0] cipher_0_ssbox_address92;
reg    cipher_0_ssbox_ce92;
wire   [7:0] cipher_0_ssbox_q92;
wire   [7:0] cipher_0_ssbox_address93;
reg    cipher_0_ssbox_ce93;
wire   [7:0] cipher_0_ssbox_q93;
wire   [7:0] cipher_0_ssbox_address94;
reg    cipher_0_ssbox_ce94;
wire   [7:0] cipher_0_ssbox_q94;
wire   [7:0] cipher_0_ssbox_address95;
reg    cipher_0_ssbox_ce95;
wire   [7:0] cipher_0_ssbox_q95;
wire   [7:0] cipher_0_ssbox_address96;
reg    cipher_0_ssbox_ce96;
wire   [7:0] cipher_0_ssbox_q96;
wire   [7:0] cipher_0_ssbox_address97;
reg    cipher_0_ssbox_ce97;
wire   [7:0] cipher_0_ssbox_q97;
wire   [7:0] cipher_0_ssbox_address98;
reg    cipher_0_ssbox_ce98;
wire   [7:0] cipher_0_ssbox_q98;
wire   [7:0] cipher_0_ssbox_address99;
reg    cipher_0_ssbox_ce99;
wire   [7:0] cipher_0_ssbox_q99;
wire   [7:0] cipher_0_ssbox_address100;
reg    cipher_0_ssbox_ce100;
wire   [7:0] cipher_0_ssbox_q100;
wire   [7:0] cipher_0_ssbox_address101;
reg    cipher_0_ssbox_ce101;
wire   [7:0] cipher_0_ssbox_q101;
wire   [7:0] cipher_0_ssbox_address102;
reg    cipher_0_ssbox_ce102;
wire   [7:0] cipher_0_ssbox_q102;
wire   [7:0] cipher_0_ssbox_address103;
reg    cipher_0_ssbox_ce103;
wire   [7:0] cipher_0_ssbox_q103;
wire   [7:0] cipher_0_ssbox_address104;
reg    cipher_0_ssbox_ce104;
wire   [7:0] cipher_0_ssbox_q104;
wire   [7:0] cipher_0_ssbox_address105;
reg    cipher_0_ssbox_ce105;
wire   [7:0] cipher_0_ssbox_q105;
wire   [7:0] cipher_0_ssbox_address106;
reg    cipher_0_ssbox_ce106;
wire   [7:0] cipher_0_ssbox_q106;
wire   [7:0] cipher_0_ssbox_address107;
reg    cipher_0_ssbox_ce107;
wire   [7:0] cipher_0_ssbox_q107;
wire   [7:0] cipher_0_ssbox_address108;
reg    cipher_0_ssbox_ce108;
wire   [7:0] cipher_0_ssbox_q108;
wire   [7:0] cipher_0_ssbox_address109;
reg    cipher_0_ssbox_ce109;
wire   [7:0] cipher_0_ssbox_q109;
wire   [7:0] cipher_0_ssbox_address110;
reg    cipher_0_ssbox_ce110;
wire   [7:0] cipher_0_ssbox_q110;
wire   [7:0] cipher_0_ssbox_address111;
reg    cipher_0_ssbox_ce111;
wire   [7:0] cipher_0_ssbox_q111;
wire   [7:0] cipher_0_ssbox_address112;
reg    cipher_0_ssbox_ce112;
wire   [7:0] cipher_0_ssbox_q112;
wire   [7:0] cipher_0_ssbox_address113;
reg    cipher_0_ssbox_ce113;
wire   [7:0] cipher_0_ssbox_q113;
wire   [7:0] cipher_0_ssbox_address114;
reg    cipher_0_ssbox_ce114;
wire   [7:0] cipher_0_ssbox_q114;
wire   [7:0] cipher_0_ssbox_address115;
reg    cipher_0_ssbox_ce115;
wire   [7:0] cipher_0_ssbox_q115;
wire   [7:0] cipher_0_ssbox_address116;
reg    cipher_0_ssbox_ce116;
wire   [7:0] cipher_0_ssbox_q116;
wire   [7:0] cipher_0_ssbox_address117;
reg    cipher_0_ssbox_ce117;
wire   [7:0] cipher_0_ssbox_q117;
wire   [7:0] cipher_0_ssbox_address118;
reg    cipher_0_ssbox_ce118;
wire   [7:0] cipher_0_ssbox_q118;
wire   [7:0] cipher_0_ssbox_address119;
reg    cipher_0_ssbox_ce119;
wire   [7:0] cipher_0_ssbox_q119;
wire   [7:0] cipher_0_ssbox_address120;
reg    cipher_0_ssbox_ce120;
wire   [7:0] cipher_0_ssbox_q120;
wire   [7:0] cipher_0_ssbox_address121;
reg    cipher_0_ssbox_ce121;
wire   [7:0] cipher_0_ssbox_q121;
wire   [7:0] cipher_0_ssbox_address122;
reg    cipher_0_ssbox_ce122;
wire   [7:0] cipher_0_ssbox_q122;
wire   [7:0] cipher_0_ssbox_address123;
reg    cipher_0_ssbox_ce123;
wire   [7:0] cipher_0_ssbox_q123;
wire   [7:0] cipher_0_ssbox_address124;
reg    cipher_0_ssbox_ce124;
wire   [7:0] cipher_0_ssbox_q124;
wire   [7:0] cipher_0_ssbox_address125;
reg    cipher_0_ssbox_ce125;
wire   [7:0] cipher_0_ssbox_q125;
wire   [7:0] cipher_0_ssbox_address126;
reg    cipher_0_ssbox_ce126;
wire   [7:0] cipher_0_ssbox_q126;
wire   [7:0] cipher_0_ssbox_address127;
reg    cipher_0_ssbox_ce127;
wire   [7:0] cipher_0_ssbox_q127;
wire   [7:0] cipher_0_ssbox_address128;
reg    cipher_0_ssbox_ce128;
wire   [7:0] cipher_0_ssbox_q128;
wire   [7:0] cipher_0_ssbox_address129;
reg    cipher_0_ssbox_ce129;
wire   [7:0] cipher_0_ssbox_q129;
wire   [7:0] cipher_0_ssbox_address130;
reg    cipher_0_ssbox_ce130;
wire   [7:0] cipher_0_ssbox_q130;
wire   [7:0] cipher_0_ssbox_address131;
reg    cipher_0_ssbox_ce131;
wire   [7:0] cipher_0_ssbox_q131;
wire   [7:0] cipher_0_ssbox_address132;
reg    cipher_0_ssbox_ce132;
wire   [7:0] cipher_0_ssbox_q132;
wire   [7:0] cipher_0_ssbox_address133;
reg    cipher_0_ssbox_ce133;
wire   [7:0] cipher_0_ssbox_q133;
wire   [7:0] cipher_0_ssbox_address134;
reg    cipher_0_ssbox_ce134;
wire   [7:0] cipher_0_ssbox_q134;
wire   [7:0] cipher_0_ssbox_address135;
reg    cipher_0_ssbox_ce135;
wire   [7:0] cipher_0_ssbox_q135;
wire   [7:0] cipher_0_ssbox_address136;
reg    cipher_0_ssbox_ce136;
wire   [7:0] cipher_0_ssbox_q136;
wire   [7:0] cipher_0_ssbox_address137;
reg    cipher_0_ssbox_ce137;
wire   [7:0] cipher_0_ssbox_q137;
wire   [7:0] cipher_0_ssbox_address138;
reg    cipher_0_ssbox_ce138;
wire   [7:0] cipher_0_ssbox_q138;
wire   [7:0] cipher_0_ssbox_address139;
reg    cipher_0_ssbox_ce139;
wire   [7:0] cipher_0_ssbox_q139;
wire   [7:0] cipher_0_ssbox_address140;
reg    cipher_0_ssbox_ce140;
wire   [7:0] cipher_0_ssbox_q140;
wire   [7:0] cipher_0_ssbox_address141;
reg    cipher_0_ssbox_ce141;
wire   [7:0] cipher_0_ssbox_q141;
wire   [7:0] cipher_0_ssbox_address142;
reg    cipher_0_ssbox_ce142;
wire   [7:0] cipher_0_ssbox_q142;
wire   [7:0] cipher_0_ssbox_address143;
reg    cipher_0_ssbox_ce143;
wire   [7:0] cipher_0_ssbox_q143;
wire   [7:0] cipher_0_ssbox_address144;
reg    cipher_0_ssbox_ce144;
wire   [7:0] cipher_0_ssbox_q144;
wire   [7:0] cipher_0_ssbox_address145;
reg    cipher_0_ssbox_ce145;
wire   [7:0] cipher_0_ssbox_q145;
wire   [7:0] cipher_0_ssbox_address146;
reg    cipher_0_ssbox_ce146;
wire   [7:0] cipher_0_ssbox_q146;
wire   [7:0] cipher_0_ssbox_address147;
reg    cipher_0_ssbox_ce147;
wire   [7:0] cipher_0_ssbox_q147;
wire   [7:0] cipher_0_ssbox_address148;
reg    cipher_0_ssbox_ce148;
wire   [7:0] cipher_0_ssbox_q148;
wire   [7:0] cipher_0_ssbox_address149;
reg    cipher_0_ssbox_ce149;
wire   [7:0] cipher_0_ssbox_q149;
wire   [7:0] cipher_0_ssbox_address150;
reg    cipher_0_ssbox_ce150;
wire   [7:0] cipher_0_ssbox_q150;
wire   [7:0] cipher_0_ssbox_address151;
reg    cipher_0_ssbox_ce151;
wire   [7:0] cipher_0_ssbox_q151;
wire   [7:0] cipher_0_ssbox_address152;
reg    cipher_0_ssbox_ce152;
wire   [7:0] cipher_0_ssbox_q152;
wire   [7:0] cipher_0_ssbox_address153;
reg    cipher_0_ssbox_ce153;
wire   [7:0] cipher_0_ssbox_q153;
wire   [7:0] cipher_0_ssbox_address154;
reg    cipher_0_ssbox_ce154;
wire   [7:0] cipher_0_ssbox_q154;
wire   [7:0] cipher_0_ssbox_address155;
reg    cipher_0_ssbox_ce155;
wire   [7:0] cipher_0_ssbox_q155;
wire   [7:0] cipher_0_ssbox_address156;
reg    cipher_0_ssbox_ce156;
wire   [7:0] cipher_0_ssbox_q156;
wire   [7:0] cipher_0_ssbox_address157;
reg    cipher_0_ssbox_ce157;
wire   [7:0] cipher_0_ssbox_q157;
wire   [7:0] cipher_0_ssbox_address158;
reg    cipher_0_ssbox_ce158;
wire   [7:0] cipher_0_ssbox_q158;
wire   [7:0] cipher_0_ssbox_address159;
reg    cipher_0_ssbox_ce159;
wire   [7:0] cipher_0_ssbox_q159;
wire   [7:0] cipher_0_ssbox_address160;
reg    cipher_0_ssbox_ce160;
wire   [7:0] cipher_0_ssbox_q160;
wire   [7:0] cipher_0_ssbox_address161;
reg    cipher_0_ssbox_ce161;
wire   [7:0] cipher_0_ssbox_q161;
wire   [7:0] cipher_0_ssbox_address162;
reg    cipher_0_ssbox_ce162;
wire   [7:0] cipher_0_ssbox_q162;
wire   [7:0] cipher_0_ssbox_address163;
reg    cipher_0_ssbox_ce163;
wire   [7:0] cipher_0_ssbox_q163;
wire   [7:0] cipher_0_ssbox_address164;
reg    cipher_0_ssbox_ce164;
wire   [7:0] cipher_0_ssbox_q164;
wire   [7:0] cipher_0_ssbox_address165;
reg    cipher_0_ssbox_ce165;
wire   [7:0] cipher_0_ssbox_q165;
wire   [7:0] cipher_0_ssbox_address166;
reg    cipher_0_ssbox_ce166;
wire   [7:0] cipher_0_ssbox_q166;
wire   [7:0] cipher_0_ssbox_address167;
reg    cipher_0_ssbox_ce167;
wire   [7:0] cipher_0_ssbox_q167;
wire   [7:0] cipher_0_ssbox_address168;
reg    cipher_0_ssbox_ce168;
wire   [7:0] cipher_0_ssbox_q168;
wire   [7:0] cipher_0_ssbox_address169;
reg    cipher_0_ssbox_ce169;
wire   [7:0] cipher_0_ssbox_q169;
wire   [7:0] cipher_0_ssbox_address170;
reg    cipher_0_ssbox_ce170;
wire   [7:0] cipher_0_ssbox_q170;
wire   [7:0] cipher_0_ssbox_address171;
reg    cipher_0_ssbox_ce171;
wire   [7:0] cipher_0_ssbox_q171;
wire   [7:0] cipher_0_ssbox_address172;
reg    cipher_0_ssbox_ce172;
wire   [7:0] cipher_0_ssbox_q172;
wire   [7:0] cipher_0_ssbox_address173;
reg    cipher_0_ssbox_ce173;
wire   [7:0] cipher_0_ssbox_q173;
wire   [7:0] cipher_0_ssbox_address174;
reg    cipher_0_ssbox_ce174;
wire   [7:0] cipher_0_ssbox_q174;
wire   [7:0] cipher_0_ssbox_address175;
reg    cipher_0_ssbox_ce175;
wire   [7:0] cipher_0_ssbox_q175;
wire   [7:0] cipher_0_ssbox_address176;
reg    cipher_0_ssbox_ce176;
wire   [7:0] cipher_0_ssbox_q176;
wire   [7:0] cipher_0_ssbox_address177;
reg    cipher_0_ssbox_ce177;
wire   [7:0] cipher_0_ssbox_q177;
wire   [7:0] cipher_0_ssbox_address178;
reg    cipher_0_ssbox_ce178;
wire   [7:0] cipher_0_ssbox_q178;
wire   [7:0] cipher_0_ssbox_address179;
reg    cipher_0_ssbox_ce179;
wire   [7:0] cipher_0_ssbox_q179;
wire   [7:0] cipher_0_ssbox_address180;
reg    cipher_0_ssbox_ce180;
wire   [7:0] cipher_0_ssbox_q180;
wire   [7:0] cipher_0_ssbox_address181;
reg    cipher_0_ssbox_ce181;
wire   [7:0] cipher_0_ssbox_q181;
wire   [7:0] cipher_0_ssbox_address182;
reg    cipher_0_ssbox_ce182;
wire   [7:0] cipher_0_ssbox_q182;
wire   [7:0] cipher_0_ssbox_address183;
reg    cipher_0_ssbox_ce183;
wire   [7:0] cipher_0_ssbox_q183;
wire   [7:0] cipher_0_ssbox_address184;
reg    cipher_0_ssbox_ce184;
wire   [7:0] cipher_0_ssbox_q184;
wire   [7:0] cipher_0_ssbox_address185;
reg    cipher_0_ssbox_ce185;
wire   [7:0] cipher_0_ssbox_q185;
wire   [7:0] cipher_0_ssbox_address186;
reg    cipher_0_ssbox_ce186;
wire   [7:0] cipher_0_ssbox_q186;
wire   [7:0] cipher_0_ssbox_address187;
reg    cipher_0_ssbox_ce187;
wire   [7:0] cipher_0_ssbox_q187;
wire   [7:0] cipher_0_ssbox_address188;
reg    cipher_0_ssbox_ce188;
wire   [7:0] cipher_0_ssbox_q188;
wire   [7:0] cipher_0_ssbox_address189;
reg    cipher_0_ssbox_ce189;
wire   [7:0] cipher_0_ssbox_q189;
wire   [7:0] cipher_0_ssbox_address190;
reg    cipher_0_ssbox_ce190;
wire   [7:0] cipher_0_ssbox_q190;
wire   [7:0] cipher_0_ssbox_address191;
reg    cipher_0_ssbox_ce191;
wire   [7:0] cipher_0_ssbox_q191;
wire   [7:0] cipher_0_p16box_address0;
reg    cipher_0_p16box_ce0;
wire   [15:0] cipher_0_p16box_q0;
wire   [7:0] cipher_0_p16box_address1;
reg    cipher_0_p16box_ce1;
wire   [15:0] cipher_0_p16box_q1;
wire   [7:0] cipher_0_p16box_address2;
reg    cipher_0_p16box_ce2;
wire   [15:0] cipher_0_p16box_q2;
wire   [7:0] cipher_0_p16box_address3;
reg    cipher_0_p16box_ce3;
wire   [15:0] cipher_0_p16box_q3;
wire   [7:0] cipher_0_p16box_address4;
reg    cipher_0_p16box_ce4;
wire   [15:0] cipher_0_p16box_q4;
wire   [7:0] cipher_0_p16box_address5;
reg    cipher_0_p16box_ce5;
wire   [15:0] cipher_0_p16box_q5;
wire   [7:0] cipher_0_p16box_address6;
reg    cipher_0_p16box_ce6;
wire   [15:0] cipher_0_p16box_q6;
wire   [7:0] cipher_0_p16box_address7;
reg    cipher_0_p16box_ce7;
wire   [15:0] cipher_0_p16box_q7;
wire   [7:0] cipher_0_p16box_address8;
reg    cipher_0_p16box_ce8;
wire   [15:0] cipher_0_p16box_q8;
wire   [7:0] cipher_0_p16box_address9;
reg    cipher_0_p16box_ce9;
wire   [15:0] cipher_0_p16box_q9;
wire   [7:0] cipher_0_p16box_address10;
reg    cipher_0_p16box_ce10;
wire   [15:0] cipher_0_p16box_q10;
wire   [7:0] cipher_0_p16box_address11;
reg    cipher_0_p16box_ce11;
wire   [15:0] cipher_0_p16box_q11;
wire   [7:0] cipher_0_p16box_address12;
reg    cipher_0_p16box_ce12;
wire   [15:0] cipher_0_p16box_q12;
wire   [7:0] cipher_0_p16box_address13;
reg    cipher_0_p16box_ce13;
wire   [15:0] cipher_0_p16box_q13;
wire   [7:0] cipher_0_p16box_address14;
reg    cipher_0_p16box_ce14;
wire   [15:0] cipher_0_p16box_q14;
wire   [7:0] cipher_0_p16box_address15;
reg    cipher_0_p16box_ce15;
wire   [15:0] cipher_0_p16box_q15;
wire   [7:0] cipher_0_p16box_address16;
reg    cipher_0_p16box_ce16;
wire   [15:0] cipher_0_p16box_q16;
wire   [7:0] cipher_0_p16box_address17;
reg    cipher_0_p16box_ce17;
wire   [15:0] cipher_0_p16box_q17;
wire   [7:0] cipher_0_p16box_address18;
reg    cipher_0_p16box_ce18;
wire   [15:0] cipher_0_p16box_q18;
wire   [7:0] cipher_0_p16box_address19;
reg    cipher_0_p16box_ce19;
wire   [15:0] cipher_0_p16box_q19;
wire   [7:0] cipher_0_p16box_address20;
reg    cipher_0_p16box_ce20;
wire   [15:0] cipher_0_p16box_q20;
wire   [7:0] cipher_0_p16box_address21;
reg    cipher_0_p16box_ce21;
wire   [15:0] cipher_0_p16box_q21;
wire   [7:0] cipher_0_p16box_address22;
reg    cipher_0_p16box_ce22;
wire   [15:0] cipher_0_p16box_q22;
wire   [7:0] cipher_0_p16box_address23;
reg    cipher_0_p16box_ce23;
wire   [15:0] cipher_0_p16box_q23;
wire   [7:0] cipher_0_p16box_address24;
reg    cipher_0_p16box_ce24;
wire   [15:0] cipher_0_p16box_q24;
wire   [7:0] cipher_0_p16box_address25;
reg    cipher_0_p16box_ce25;
wire   [15:0] cipher_0_p16box_q25;
wire   [7:0] cipher_0_p16box_address26;
reg    cipher_0_p16box_ce26;
wire   [15:0] cipher_0_p16box_q26;
wire   [7:0] cipher_0_p16box_address27;
reg    cipher_0_p16box_ce27;
wire   [15:0] cipher_0_p16box_q27;
wire   [7:0] cipher_0_p16box_address28;
reg    cipher_0_p16box_ce28;
wire   [15:0] cipher_0_p16box_q28;
wire   [7:0] cipher_0_p16box_address29;
reg    cipher_0_p16box_ce29;
wire   [15:0] cipher_0_p16box_q29;
wire   [7:0] cipher_0_p16box_address30;
reg    cipher_0_p16box_ce30;
wire   [15:0] cipher_0_p16box_q30;
wire   [7:0] cipher_0_p16box_address31;
reg    cipher_0_p16box_ce31;
wire   [15:0] cipher_0_p16box_q31;
wire   [7:0] cipher_0_p16box_address32;
reg    cipher_0_p16box_ce32;
wire   [15:0] cipher_0_p16box_q32;
wire   [7:0] cipher_0_p16box_address33;
reg    cipher_0_p16box_ce33;
wire   [15:0] cipher_0_p16box_q33;
wire   [7:0] cipher_0_p16box_address34;
reg    cipher_0_p16box_ce34;
wire   [15:0] cipher_0_p16box_q34;
wire   [7:0] cipher_0_p16box_address35;
reg    cipher_0_p16box_ce35;
wire   [15:0] cipher_0_p16box_q35;
wire   [7:0] cipher_0_p16box_address36;
reg    cipher_0_p16box_ce36;
wire   [15:0] cipher_0_p16box_q36;
wire   [7:0] cipher_0_p16box_address37;
reg    cipher_0_p16box_ce37;
wire   [15:0] cipher_0_p16box_q37;
wire   [7:0] cipher_0_p16box_address38;
reg    cipher_0_p16box_ce38;
wire   [15:0] cipher_0_p16box_q38;
wire   [7:0] cipher_0_p16box_address39;
reg    cipher_0_p16box_ce39;
wire   [15:0] cipher_0_p16box_q39;
wire   [7:0] cipher_0_p16box_address40;
reg    cipher_0_p16box_ce40;
wire   [15:0] cipher_0_p16box_q40;
wire   [7:0] cipher_0_p16box_address41;
reg    cipher_0_p16box_ce41;
wire   [15:0] cipher_0_p16box_q41;
wire   [7:0] cipher_0_p16box_address42;
reg    cipher_0_p16box_ce42;
wire   [15:0] cipher_0_p16box_q42;
wire   [7:0] cipher_0_p16box_address43;
reg    cipher_0_p16box_ce43;
wire   [15:0] cipher_0_p16box_q43;
wire   [7:0] cipher_0_p16box_address44;
reg    cipher_0_p16box_ce44;
wire   [15:0] cipher_0_p16box_q44;
wire   [7:0] cipher_0_p16box_address45;
reg    cipher_0_p16box_ce45;
wire   [15:0] cipher_0_p16box_q45;
wire   [7:0] cipher_0_p16box_address46;
reg    cipher_0_p16box_ce46;
wire   [15:0] cipher_0_p16box_q46;
wire   [7:0] cipher_0_p16box_address47;
reg    cipher_0_p16box_ce47;
wire   [15:0] cipher_0_p16box_q47;
wire   [7:0] cipher_0_p16box_address48;
reg    cipher_0_p16box_ce48;
wire   [15:0] cipher_0_p16box_q48;
wire   [7:0] cipher_0_p16box_address49;
reg    cipher_0_p16box_ce49;
wire   [15:0] cipher_0_p16box_q49;
wire   [7:0] cipher_0_p16box_address50;
reg    cipher_0_p16box_ce50;
wire   [15:0] cipher_0_p16box_q50;
wire   [7:0] cipher_0_p16box_address51;
reg    cipher_0_p16box_ce51;
wire   [15:0] cipher_0_p16box_q51;
wire   [7:0] cipher_0_p16box_address52;
reg    cipher_0_p16box_ce52;
wire   [15:0] cipher_0_p16box_q52;
wire   [7:0] cipher_0_p16box_address53;
reg    cipher_0_p16box_ce53;
wire   [15:0] cipher_0_p16box_q53;
wire   [7:0] cipher_0_p16box_address54;
reg    cipher_0_p16box_ce54;
wire   [15:0] cipher_0_p16box_q54;
wire   [7:0] cipher_0_p16box_address55;
reg    cipher_0_p16box_ce55;
wire   [15:0] cipher_0_p16box_q55;
wire   [7:0] cipher_0_p16box_address56;
reg    cipher_0_p16box_ce56;
wire   [15:0] cipher_0_p16box_q56;
wire   [7:0] cipher_0_p16box_address57;
reg    cipher_0_p16box_ce57;
wire   [15:0] cipher_0_p16box_q57;
wire   [7:0] cipher_0_p16box_address58;
reg    cipher_0_p16box_ce58;
wire   [15:0] cipher_0_p16box_q58;
wire   [7:0] cipher_0_p16box_address59;
reg    cipher_0_p16box_ce59;
wire   [15:0] cipher_0_p16box_q59;
wire   [7:0] cipher_0_p16box_address60;
reg    cipher_0_p16box_ce60;
wire   [15:0] cipher_0_p16box_q60;
wire   [7:0] cipher_0_p16box_address61;
reg    cipher_0_p16box_ce61;
wire   [15:0] cipher_0_p16box_q61;
wire   [7:0] cipher_0_p16box_address62;
reg    cipher_0_p16box_ce62;
wire   [15:0] cipher_0_p16box_q62;
wire   [7:0] cipher_0_p16box_address63;
reg    cipher_0_p16box_ce63;
wire   [15:0] cipher_0_p16box_q63;
wire   [7:0] cipher_0_p16box_address64;
reg    cipher_0_p16box_ce64;
wire   [15:0] cipher_0_p16box_q64;
wire   [7:0] cipher_0_p16box_address65;
reg    cipher_0_p16box_ce65;
wire   [15:0] cipher_0_p16box_q65;
wire   [7:0] cipher_0_p16box_address66;
reg    cipher_0_p16box_ce66;
wire   [15:0] cipher_0_p16box_q66;
wire   [7:0] cipher_0_p16box_address67;
reg    cipher_0_p16box_ce67;
wire   [15:0] cipher_0_p16box_q67;
wire   [7:0] cipher_0_p16box_address68;
reg    cipher_0_p16box_ce68;
wire   [15:0] cipher_0_p16box_q68;
wire   [7:0] cipher_0_p16box_address69;
reg    cipher_0_p16box_ce69;
wire   [15:0] cipher_0_p16box_q69;
wire   [7:0] cipher_0_p16box_address70;
reg    cipher_0_p16box_ce70;
wire   [15:0] cipher_0_p16box_q70;
wire   [7:0] cipher_0_p16box_address71;
reg    cipher_0_p16box_ce71;
wire   [15:0] cipher_0_p16box_q71;
wire   [7:0] cipher_0_p16box_address72;
reg    cipher_0_p16box_ce72;
wire   [15:0] cipher_0_p16box_q72;
wire   [7:0] cipher_0_p16box_address73;
reg    cipher_0_p16box_ce73;
wire   [15:0] cipher_0_p16box_q73;
wire   [7:0] cipher_0_p16box_address74;
reg    cipher_0_p16box_ce74;
wire   [15:0] cipher_0_p16box_q74;
wire   [7:0] cipher_0_p16box_address75;
reg    cipher_0_p16box_ce75;
wire   [15:0] cipher_0_p16box_q75;
wire   [7:0] cipher_0_p16box_address76;
reg    cipher_0_p16box_ce76;
wire   [15:0] cipher_0_p16box_q76;
wire   [7:0] cipher_0_p16box_address77;
reg    cipher_0_p16box_ce77;
wire   [15:0] cipher_0_p16box_q77;
wire   [7:0] cipher_0_p16box_address78;
reg    cipher_0_p16box_ce78;
wire   [15:0] cipher_0_p16box_q78;
wire   [7:0] cipher_0_p16box_address79;
reg    cipher_0_p16box_ce79;
wire   [15:0] cipher_0_p16box_q79;
wire   [7:0] cipher_0_p16box_address80;
reg    cipher_0_p16box_ce80;
wire   [15:0] cipher_0_p16box_q80;
wire   [7:0] cipher_0_p16box_address81;
reg    cipher_0_p16box_ce81;
wire   [15:0] cipher_0_p16box_q81;
wire   [7:0] cipher_0_p16box_address82;
reg    cipher_0_p16box_ce82;
wire   [15:0] cipher_0_p16box_q82;
wire   [7:0] cipher_0_p16box_address83;
reg    cipher_0_p16box_ce83;
wire   [15:0] cipher_0_p16box_q83;
wire   [7:0] cipher_0_p16box_address84;
reg    cipher_0_p16box_ce84;
wire   [15:0] cipher_0_p16box_q84;
wire   [7:0] cipher_0_p16box_address85;
reg    cipher_0_p16box_ce85;
wire   [15:0] cipher_0_p16box_q85;
wire   [7:0] cipher_0_p16box_address86;
reg    cipher_0_p16box_ce86;
wire   [15:0] cipher_0_p16box_q86;
wire   [7:0] cipher_0_p16box_address87;
reg    cipher_0_p16box_ce87;
wire   [15:0] cipher_0_p16box_q87;
wire   [7:0] cipher_0_p16box_address88;
reg    cipher_0_p16box_ce88;
wire   [15:0] cipher_0_p16box_q88;
wire   [7:0] cipher_0_p16box_address89;
reg    cipher_0_p16box_ce89;
wire   [15:0] cipher_0_p16box_q89;
wire   [7:0] cipher_0_p16box_address90;
reg    cipher_0_p16box_ce90;
wire   [15:0] cipher_0_p16box_q90;
wire   [7:0] cipher_0_p16box_address91;
reg    cipher_0_p16box_ce91;
wire   [15:0] cipher_0_p16box_q91;
wire   [7:0] cipher_0_p16box_address92;
reg    cipher_0_p16box_ce92;
wire   [15:0] cipher_0_p16box_q92;
wire   [7:0] cipher_0_p16box_address93;
reg    cipher_0_p16box_ce93;
wire   [15:0] cipher_0_p16box_q93;
wire   [7:0] cipher_0_p16box_address94;
reg    cipher_0_p16box_ce94;
wire   [15:0] cipher_0_p16box_q94;
wire   [7:0] cipher_0_p16box_address95;
reg    cipher_0_p16box_ce95;
wire   [15:0] cipher_0_p16box_q95;
wire   [7:0] cipher_0_p16box_address96;
reg    cipher_0_p16box_ce96;
wire   [15:0] cipher_0_p16box_q96;
wire   [7:0] cipher_0_p16box_address97;
reg    cipher_0_p16box_ce97;
wire   [15:0] cipher_0_p16box_q97;
wire   [7:0] cipher_0_p16box_address98;
reg    cipher_0_p16box_ce98;
wire   [15:0] cipher_0_p16box_q98;
wire   [7:0] cipher_0_p16box_address99;
reg    cipher_0_p16box_ce99;
wire   [15:0] cipher_0_p16box_q99;
wire   [7:0] cipher_0_p16box_address100;
reg    cipher_0_p16box_ce100;
wire   [15:0] cipher_0_p16box_q100;
wire   [7:0] cipher_0_p16box_address101;
reg    cipher_0_p16box_ce101;
wire   [15:0] cipher_0_p16box_q101;
wire   [7:0] cipher_0_p16box_address102;
reg    cipher_0_p16box_ce102;
wire   [15:0] cipher_0_p16box_q102;
wire   [7:0] cipher_0_p16box_address103;
reg    cipher_0_p16box_ce103;
wire   [15:0] cipher_0_p16box_q103;
wire   [7:0] cipher_0_p16box_address104;
reg    cipher_0_p16box_ce104;
wire   [15:0] cipher_0_p16box_q104;
wire   [7:0] cipher_0_p16box_address105;
reg    cipher_0_p16box_ce105;
wire   [15:0] cipher_0_p16box_q105;
wire   [7:0] cipher_0_p16box_address106;
reg    cipher_0_p16box_ce106;
wire   [15:0] cipher_0_p16box_q106;
wire   [7:0] cipher_0_p16box_address107;
reg    cipher_0_p16box_ce107;
wire   [15:0] cipher_0_p16box_q107;
wire   [7:0] cipher_0_p16box_address108;
reg    cipher_0_p16box_ce108;
wire   [15:0] cipher_0_p16box_q108;
wire   [7:0] cipher_0_p16box_address109;
reg    cipher_0_p16box_ce109;
wire   [15:0] cipher_0_p16box_q109;
wire   [7:0] cipher_0_p16box_address110;
reg    cipher_0_p16box_ce110;
wire   [15:0] cipher_0_p16box_q110;
wire   [7:0] cipher_0_p16box_address111;
reg    cipher_0_p16box_ce111;
wire   [15:0] cipher_0_p16box_q111;
wire   [7:0] cipher_0_p16box_address112;
reg    cipher_0_p16box_ce112;
wire   [15:0] cipher_0_p16box_q112;
wire   [7:0] cipher_0_p16box_address113;
reg    cipher_0_p16box_ce113;
wire   [15:0] cipher_0_p16box_q113;
wire   [7:0] cipher_0_p16box_address114;
reg    cipher_0_p16box_ce114;
wire   [15:0] cipher_0_p16box_q114;
wire   [7:0] cipher_0_p16box_address115;
reg    cipher_0_p16box_ce115;
wire   [15:0] cipher_0_p16box_q115;
wire   [7:0] cipher_0_p16box_address116;
reg    cipher_0_p16box_ce116;
wire   [15:0] cipher_0_p16box_q116;
wire   [7:0] cipher_0_p16box_address117;
reg    cipher_0_p16box_ce117;
wire   [15:0] cipher_0_p16box_q117;
wire   [7:0] cipher_0_p16box_address118;
reg    cipher_0_p16box_ce118;
wire   [15:0] cipher_0_p16box_q118;
wire   [7:0] cipher_0_p16box_address119;
reg    cipher_0_p16box_ce119;
wire   [15:0] cipher_0_p16box_q119;
wire   [7:0] cipher_0_p16box_address120;
reg    cipher_0_p16box_ce120;
wire   [15:0] cipher_0_p16box_q120;
wire   [7:0] cipher_0_p16box_address121;
reg    cipher_0_p16box_ce121;
wire   [15:0] cipher_0_p16box_q121;
wire   [7:0] cipher_0_p16box_address122;
reg    cipher_0_p16box_ce122;
wire   [15:0] cipher_0_p16box_q122;
wire   [7:0] cipher_0_p16box_address123;
reg    cipher_0_p16box_ce123;
wire   [15:0] cipher_0_p16box_q123;
wire   [7:0] cipher_0_p16box_address124;
reg    cipher_0_p16box_ce124;
wire   [15:0] cipher_0_p16box_q124;
wire   [7:0] cipher_0_p16box_address125;
reg    cipher_0_p16box_ce125;
wire   [15:0] cipher_0_p16box_q125;
wire   [7:0] cipher_0_p16box_address126;
reg    cipher_0_p16box_ce126;
wire   [15:0] cipher_0_p16box_q126;
wire   [7:0] cipher_0_p16box_address127;
reg    cipher_0_p16box_ce127;
wire   [15:0] cipher_0_p16box_q127;
wire   [7:0] cipher_0_p16box_address128;
reg    cipher_0_p16box_ce128;
wire   [15:0] cipher_0_p16box_q128;
wire   [7:0] cipher_0_p16box_address129;
reg    cipher_0_p16box_ce129;
wire   [15:0] cipher_0_p16box_q129;
wire   [7:0] cipher_0_p16box_address130;
reg    cipher_0_p16box_ce130;
wire   [15:0] cipher_0_p16box_q130;
wire   [7:0] cipher_0_p16box_address131;
reg    cipher_0_p16box_ce131;
wire   [15:0] cipher_0_p16box_q131;
wire   [7:0] cipher_0_p16box_address132;
reg    cipher_0_p16box_ce132;
wire   [15:0] cipher_0_p16box_q132;
wire   [7:0] cipher_0_p16box_address133;
reg    cipher_0_p16box_ce133;
wire   [15:0] cipher_0_p16box_q133;
wire   [7:0] cipher_0_p16box_address134;
reg    cipher_0_p16box_ce134;
wire   [15:0] cipher_0_p16box_q134;
wire   [7:0] cipher_0_p16box_address135;
reg    cipher_0_p16box_ce135;
wire   [15:0] cipher_0_p16box_q135;
wire   [7:0] cipher_0_p16box_address136;
reg    cipher_0_p16box_ce136;
wire   [15:0] cipher_0_p16box_q136;
wire   [7:0] cipher_0_p16box_address137;
reg    cipher_0_p16box_ce137;
wire   [15:0] cipher_0_p16box_q137;
wire   [7:0] cipher_0_p16box_address138;
reg    cipher_0_p16box_ce138;
wire   [15:0] cipher_0_p16box_q138;
wire   [7:0] cipher_0_p16box_address139;
reg    cipher_0_p16box_ce139;
wire   [15:0] cipher_0_p16box_q139;
wire   [7:0] cipher_0_p16box_address140;
reg    cipher_0_p16box_ce140;
wire   [15:0] cipher_0_p16box_q140;
wire   [7:0] cipher_0_p16box_address141;
reg    cipher_0_p16box_ce141;
wire   [15:0] cipher_0_p16box_q141;
wire   [7:0] cipher_0_p16box_address142;
reg    cipher_0_p16box_ce142;
wire   [15:0] cipher_0_p16box_q142;
wire   [7:0] cipher_0_p16box_address143;
reg    cipher_0_p16box_ce143;
wire   [15:0] cipher_0_p16box_q143;
wire   [7:0] cipher_0_p16box_address144;
reg    cipher_0_p16box_ce144;
wire   [15:0] cipher_0_p16box_q144;
wire   [7:0] cipher_0_p16box_address145;
reg    cipher_0_p16box_ce145;
wire   [15:0] cipher_0_p16box_q145;
wire   [7:0] cipher_0_p16box_address146;
reg    cipher_0_p16box_ce146;
wire   [15:0] cipher_0_p16box_q146;
wire   [7:0] cipher_0_p16box_address147;
reg    cipher_0_p16box_ce147;
wire   [15:0] cipher_0_p16box_q147;
wire   [7:0] cipher_0_p16box_address148;
reg    cipher_0_p16box_ce148;
wire   [15:0] cipher_0_p16box_q148;
wire   [7:0] cipher_0_p16box_address149;
reg    cipher_0_p16box_ce149;
wire   [15:0] cipher_0_p16box_q149;
wire   [7:0] cipher_0_p16box_address150;
reg    cipher_0_p16box_ce150;
wire   [15:0] cipher_0_p16box_q150;
wire   [7:0] cipher_0_p16box_address151;
reg    cipher_0_p16box_ce151;
wire   [15:0] cipher_0_p16box_q151;
wire   [7:0] cipher_0_p16box_address152;
reg    cipher_0_p16box_ce152;
wire   [15:0] cipher_0_p16box_q152;
wire   [7:0] cipher_0_p16box_address153;
reg    cipher_0_p16box_ce153;
wire   [15:0] cipher_0_p16box_q153;
wire   [7:0] cipher_0_p16box_address154;
reg    cipher_0_p16box_ce154;
wire   [15:0] cipher_0_p16box_q154;
wire   [7:0] cipher_0_p16box_address155;
reg    cipher_0_p16box_ce155;
wire   [15:0] cipher_0_p16box_q155;
wire   [7:0] cipher_0_p16box_address156;
reg    cipher_0_p16box_ce156;
wire   [15:0] cipher_0_p16box_q156;
wire   [7:0] cipher_0_p16box_address157;
reg    cipher_0_p16box_ce157;
wire   [15:0] cipher_0_p16box_q157;
wire   [7:0] cipher_0_p16box_address158;
reg    cipher_0_p16box_ce158;
wire   [15:0] cipher_0_p16box_q158;
wire   [7:0] cipher_0_p16box_address159;
reg    cipher_0_p16box_ce159;
wire   [15:0] cipher_0_p16box_q159;
wire   [7:0] cipher_0_p16box_address160;
reg    cipher_0_p16box_ce160;
wire   [15:0] cipher_0_p16box_q160;
wire   [7:0] cipher_0_p16box_address161;
reg    cipher_0_p16box_ce161;
wire   [15:0] cipher_0_p16box_q161;
wire   [7:0] cipher_0_p16box_address162;
reg    cipher_0_p16box_ce162;
wire   [15:0] cipher_0_p16box_q162;
wire   [7:0] cipher_0_p16box_address163;
reg    cipher_0_p16box_ce163;
wire   [15:0] cipher_0_p16box_q163;
wire   [7:0] cipher_0_p16box_address164;
reg    cipher_0_p16box_ce164;
wire   [15:0] cipher_0_p16box_q164;
wire   [7:0] cipher_0_p16box_address165;
reg    cipher_0_p16box_ce165;
wire   [15:0] cipher_0_p16box_q165;
wire   [7:0] cipher_0_p16box_address166;
reg    cipher_0_p16box_ce166;
wire   [15:0] cipher_0_p16box_q166;
wire   [7:0] cipher_0_p16box_address167;
reg    cipher_0_p16box_ce167;
wire   [15:0] cipher_0_p16box_q167;
wire   [7:0] cipher_0_p16box_address168;
reg    cipher_0_p16box_ce168;
wire   [15:0] cipher_0_p16box_q168;
wire   [7:0] cipher_0_p16box_address169;
reg    cipher_0_p16box_ce169;
wire   [15:0] cipher_0_p16box_q169;
wire   [7:0] cipher_0_p16box_address170;
reg    cipher_0_p16box_ce170;
wire   [15:0] cipher_0_p16box_q170;
wire   [7:0] cipher_0_p16box_address171;
reg    cipher_0_p16box_ce171;
wire   [15:0] cipher_0_p16box_q171;
wire   [7:0] cipher_0_p16box_address172;
reg    cipher_0_p16box_ce172;
wire   [15:0] cipher_0_p16box_q172;
wire   [7:0] cipher_0_p16box_address173;
reg    cipher_0_p16box_ce173;
wire   [15:0] cipher_0_p16box_q173;
wire   [7:0] cipher_0_p16box_address174;
reg    cipher_0_p16box_ce174;
wire   [15:0] cipher_0_p16box_q174;
wire   [7:0] cipher_0_p16box_address175;
reg    cipher_0_p16box_ce175;
wire   [15:0] cipher_0_p16box_q175;
reg   [127:0] p_read_1_reg_14078;
wire    ap_block_pp0_stage0_11001;
reg   [127:0] p_read_1_reg_14078_pp0_iter1_reg;
reg   [127:0] p_read_1_reg_14078_pp0_iter2_reg;
reg   [127:0] p_read_1_reg_14078_pp0_iter3_reg;
reg   [127:0] p_read_1_reg_14078_pp0_iter4_reg;
reg   [127:0] p_read_1_reg_14078_pp0_iter5_reg;
reg   [127:0] p_read_1_reg_14078_pp0_iter6_reg;
reg   [127:0] p_read_1_reg_14078_pp0_iter7_reg;
reg   [127:0] p_read_1_reg_14078_pp0_iter8_reg;
reg   [127:0] p_read_1_reg_14078_pp0_iter9_reg;
reg   [127:0] p_read_1_reg_14078_pp0_iter10_reg;
reg   [127:0] p_read_1_reg_14078_pp0_iter11_reg;
reg   [127:0] p_read_1_reg_14078_pp0_iter12_reg;
reg   [127:0] p_read_1_reg_14078_pp0_iter13_reg;
reg   [127:0] p_read_1_reg_14078_pp0_iter14_reg;
reg   [127:0] p_read_1_reg_14078_pp0_iter15_reg;
reg   [127:0] p_read_1_reg_14078_pp0_iter16_reg;
reg   [127:0] p_read_1_reg_14078_pp0_iter17_reg;
reg   [127:0] p_read_1_reg_14078_pp0_iter18_reg;
reg   [127:0] p_read_1_reg_14078_pp0_iter19_reg;
reg   [127:0] p_read_1_reg_14078_pp0_iter20_reg;
reg   [127:0] p_read_1_reg_14078_pp0_iter21_reg;
reg   [127:0] p_read_1_reg_14078_pp0_iter22_reg;
reg   [127:0] p_read_2_reg_14083;
reg   [127:0] p_read_2_reg_14083_pp0_iter1_reg;
reg   [127:0] p_read_2_reg_14083_pp0_iter2_reg;
reg   [127:0] p_read_2_reg_14083_pp0_iter3_reg;
reg   [127:0] p_read_2_reg_14083_pp0_iter4_reg;
reg   [127:0] p_read_2_reg_14083_pp0_iter5_reg;
reg   [127:0] p_read_2_reg_14083_pp0_iter6_reg;
reg   [127:0] p_read_2_reg_14083_pp0_iter7_reg;
reg   [127:0] p_read_2_reg_14083_pp0_iter8_reg;
reg   [127:0] p_read_2_reg_14083_pp0_iter9_reg;
reg   [127:0] p_read_2_reg_14083_pp0_iter10_reg;
reg   [127:0] p_read_2_reg_14083_pp0_iter11_reg;
reg   [127:0] p_read_2_reg_14083_pp0_iter12_reg;
reg   [127:0] p_read_2_reg_14083_pp0_iter13_reg;
reg   [127:0] p_read_2_reg_14083_pp0_iter14_reg;
reg   [127:0] p_read_2_reg_14083_pp0_iter15_reg;
reg   [127:0] p_read_2_reg_14083_pp0_iter16_reg;
reg   [127:0] p_read_2_reg_14083_pp0_iter17_reg;
reg   [127:0] p_read_2_reg_14083_pp0_iter18_reg;
reg   [127:0] p_read_2_reg_14083_pp0_iter19_reg;
reg   [127:0] p_read_2_reg_14083_pp0_iter20_reg;
reg   [127:0] p_read_2_reg_14083_pp0_iter21_reg;
reg   [127:0] p_read_3_reg_14088;
reg   [127:0] p_read_3_reg_14088_pp0_iter1_reg;
reg   [127:0] p_read_3_reg_14088_pp0_iter2_reg;
reg   [127:0] p_read_3_reg_14088_pp0_iter3_reg;
reg   [127:0] p_read_3_reg_14088_pp0_iter4_reg;
reg   [127:0] p_read_3_reg_14088_pp0_iter5_reg;
reg   [127:0] p_read_3_reg_14088_pp0_iter6_reg;
reg   [127:0] p_read_3_reg_14088_pp0_iter7_reg;
reg   [127:0] p_read_3_reg_14088_pp0_iter8_reg;
reg   [127:0] p_read_3_reg_14088_pp0_iter9_reg;
reg   [127:0] p_read_3_reg_14088_pp0_iter10_reg;
reg   [127:0] p_read_3_reg_14088_pp0_iter11_reg;
reg   [127:0] p_read_3_reg_14088_pp0_iter12_reg;
reg   [127:0] p_read_3_reg_14088_pp0_iter13_reg;
reg   [127:0] p_read_3_reg_14088_pp0_iter14_reg;
reg   [127:0] p_read_3_reg_14088_pp0_iter15_reg;
reg   [127:0] p_read_3_reg_14088_pp0_iter16_reg;
reg   [127:0] p_read_3_reg_14088_pp0_iter17_reg;
reg   [127:0] p_read_3_reg_14088_pp0_iter18_reg;
reg   [127:0] p_read_3_reg_14088_pp0_iter19_reg;
reg   [127:0] p_read_4_reg_14093;
reg   [127:0] p_read_4_reg_14093_pp0_iter1_reg;
reg   [127:0] p_read_4_reg_14093_pp0_iter2_reg;
reg   [127:0] p_read_4_reg_14093_pp0_iter3_reg;
reg   [127:0] p_read_4_reg_14093_pp0_iter4_reg;
reg   [127:0] p_read_4_reg_14093_pp0_iter5_reg;
reg   [127:0] p_read_4_reg_14093_pp0_iter6_reg;
reg   [127:0] p_read_4_reg_14093_pp0_iter7_reg;
reg   [127:0] p_read_4_reg_14093_pp0_iter8_reg;
reg   [127:0] p_read_4_reg_14093_pp0_iter9_reg;
reg   [127:0] p_read_4_reg_14093_pp0_iter10_reg;
reg   [127:0] p_read_4_reg_14093_pp0_iter11_reg;
reg   [127:0] p_read_4_reg_14093_pp0_iter12_reg;
reg   [127:0] p_read_4_reg_14093_pp0_iter13_reg;
reg   [127:0] p_read_4_reg_14093_pp0_iter14_reg;
reg   [127:0] p_read_4_reg_14093_pp0_iter15_reg;
reg   [127:0] p_read_4_reg_14093_pp0_iter16_reg;
reg   [127:0] p_read_4_reg_14093_pp0_iter17_reg;
reg   [127:0] p_read_5_reg_14098;
reg   [127:0] p_read_5_reg_14098_pp0_iter1_reg;
reg   [127:0] p_read_5_reg_14098_pp0_iter2_reg;
reg   [127:0] p_read_5_reg_14098_pp0_iter3_reg;
reg   [127:0] p_read_5_reg_14098_pp0_iter4_reg;
reg   [127:0] p_read_5_reg_14098_pp0_iter5_reg;
reg   [127:0] p_read_5_reg_14098_pp0_iter6_reg;
reg   [127:0] p_read_5_reg_14098_pp0_iter7_reg;
reg   [127:0] p_read_5_reg_14098_pp0_iter8_reg;
reg   [127:0] p_read_5_reg_14098_pp0_iter9_reg;
reg   [127:0] p_read_5_reg_14098_pp0_iter10_reg;
reg   [127:0] p_read_5_reg_14098_pp0_iter11_reg;
reg   [127:0] p_read_5_reg_14098_pp0_iter12_reg;
reg   [127:0] p_read_5_reg_14098_pp0_iter13_reg;
reg   [127:0] p_read_5_reg_14098_pp0_iter14_reg;
reg   [127:0] p_read_5_reg_14098_pp0_iter15_reg;
reg   [127:0] p_read_6_reg_14103;
reg   [127:0] p_read_6_reg_14103_pp0_iter1_reg;
reg   [127:0] p_read_6_reg_14103_pp0_iter2_reg;
reg   [127:0] p_read_6_reg_14103_pp0_iter3_reg;
reg   [127:0] p_read_6_reg_14103_pp0_iter4_reg;
reg   [127:0] p_read_6_reg_14103_pp0_iter5_reg;
reg   [127:0] p_read_6_reg_14103_pp0_iter6_reg;
reg   [127:0] p_read_6_reg_14103_pp0_iter7_reg;
reg   [127:0] p_read_6_reg_14103_pp0_iter8_reg;
reg   [127:0] p_read_6_reg_14103_pp0_iter9_reg;
reg   [127:0] p_read_6_reg_14103_pp0_iter10_reg;
reg   [127:0] p_read_6_reg_14103_pp0_iter11_reg;
reg   [127:0] p_read_6_reg_14103_pp0_iter12_reg;
reg   [127:0] p_read_6_reg_14103_pp0_iter13_reg;
reg   [127:0] p_read_7_reg_14108;
reg   [127:0] p_read_7_reg_14108_pp0_iter1_reg;
reg   [127:0] p_read_7_reg_14108_pp0_iter2_reg;
reg   [127:0] p_read_7_reg_14108_pp0_iter3_reg;
reg   [127:0] p_read_7_reg_14108_pp0_iter4_reg;
reg   [127:0] p_read_7_reg_14108_pp0_iter5_reg;
reg   [127:0] p_read_7_reg_14108_pp0_iter6_reg;
reg   [127:0] p_read_7_reg_14108_pp0_iter7_reg;
reg   [127:0] p_read_7_reg_14108_pp0_iter8_reg;
reg   [127:0] p_read_7_reg_14108_pp0_iter9_reg;
reg   [127:0] p_read_7_reg_14108_pp0_iter10_reg;
reg   [127:0] p_read_7_reg_14108_pp0_iter11_reg;
reg   [127:0] p_read_8_reg_14113;
reg   [127:0] p_read_8_reg_14113_pp0_iter1_reg;
reg   [127:0] p_read_8_reg_14113_pp0_iter2_reg;
reg   [127:0] p_read_8_reg_14113_pp0_iter3_reg;
reg   [127:0] p_read_8_reg_14113_pp0_iter4_reg;
reg   [127:0] p_read_8_reg_14113_pp0_iter5_reg;
reg   [127:0] p_read_8_reg_14113_pp0_iter6_reg;
reg   [127:0] p_read_8_reg_14113_pp0_iter7_reg;
reg   [127:0] p_read_8_reg_14113_pp0_iter8_reg;
reg   [127:0] p_read_8_reg_14113_pp0_iter9_reg;
reg   [127:0] p_read_9_reg_14118;
reg   [127:0] p_read_9_reg_14118_pp0_iter1_reg;
reg   [127:0] p_read_9_reg_14118_pp0_iter2_reg;
reg   [127:0] p_read_9_reg_14118_pp0_iter3_reg;
reg   [127:0] p_read_9_reg_14118_pp0_iter4_reg;
reg   [127:0] p_read_9_reg_14118_pp0_iter5_reg;
reg   [127:0] p_read_9_reg_14118_pp0_iter6_reg;
reg   [127:0] p_read_9_reg_14118_pp0_iter7_reg;
reg   [127:0] p_read_10_reg_14123;
reg   [127:0] p_read_10_reg_14123_pp0_iter1_reg;
reg   [127:0] p_read_10_reg_14123_pp0_iter2_reg;
reg   [127:0] p_read_10_reg_14123_pp0_iter3_reg;
reg   [127:0] p_read_10_reg_14123_pp0_iter4_reg;
reg   [127:0] p_read_10_reg_14123_pp0_iter5_reg;
reg   [127:0] p_read_11_reg_14128;
reg   [127:0] p_read_11_reg_14128_pp0_iter1_reg;
reg   [127:0] p_read_11_reg_14128_pp0_iter2_reg;
reg   [127:0] p_read_11_reg_14128_pp0_iter3_reg;
reg   [127:0] p_read_12_reg_14133;
reg   [127:0] p_read_12_reg_14133_pp0_iter1_reg;
reg   [7:0] tmp_V_reg_14218;
reg   [7:0] tmp_1_V_12_reg_14224;
reg   [7:0] tmp_2_1_V_12_reg_14230;
reg   [7:0] tmp_V_7_reg_14236;
reg   [7:0] tmp_V_4_reg_14242;
reg   [7:0] tmp_V_1_reg_14248;
reg   [7:0] tmp_2_2_V_12_reg_14254;
reg   [7:0] tmp_V_11_reg_14260;
reg   [7:0] tmp_V_8_reg_14266;
reg   [7:0] tmp_V_5_reg_14272;
reg   [7:0] tmp_V_2_reg_14278;
reg   [7:0] tmp_V_15_reg_14284;
reg   [7:0] tmp_V_12_reg_14290;
reg   [7:0] tmp_V_9_reg_14296;
reg   [7:0] tmp_V_6_reg_14302;
reg   [7:0] tmp_3_V_12_reg_14308;
reg   [7:0] tmp_V_16_reg_14474;
reg   [7:0] tmp_1_V_13_reg_14480;
reg   [7:0] tmp_2_1_V_13_reg_14486;
reg   [7:0] tmp_V_23_reg_14492;
reg   [7:0] tmp_V_20_reg_14498;
reg   [7:0] tmp_V_17_reg_14504;
reg   [7:0] tmp_2_2_V_13_reg_14510;
reg   [7:0] tmp_V_27_reg_14516;
reg   [7:0] tmp_V_24_reg_14522;
reg   [7:0] tmp_V_21_reg_14528;
reg   [7:0] tmp_V_18_reg_14534;
reg   [7:0] tmp_V_31_reg_14540;
reg   [7:0] tmp_V_28_reg_14546;
reg   [7:0] tmp_V_25_reg_14552;
reg   [7:0] tmp_V_22_reg_14558;
reg   [7:0] tmp_3_V_13_reg_14564;
reg   [7:0] tmp_V_32_reg_14730;
reg   [7:0] tmp_1_V_14_reg_14736;
reg   [7:0] tmp_2_1_V_14_reg_14742;
reg   [7:0] tmp_V_39_reg_14748;
reg   [7:0] tmp_V_36_reg_14754;
reg   [7:0] tmp_V_33_reg_14760;
reg   [7:0] tmp_2_2_V_14_reg_14766;
reg   [7:0] tmp_V_43_reg_14772;
reg   [7:0] tmp_V_40_reg_14778;
reg   [7:0] tmp_V_37_reg_14784;
reg   [7:0] tmp_V_34_reg_14790;
reg   [7:0] tmp_V_47_reg_14796;
reg   [7:0] tmp_V_44_reg_14802;
reg   [7:0] tmp_V_41_reg_14808;
reg   [7:0] tmp_V_38_reg_14814;
reg   [7:0] tmp_3_V_14_reg_14820;
reg   [7:0] tmp_V_48_reg_14986;
reg   [7:0] tmp_1_V_15_reg_14992;
reg   [7:0] tmp_2_1_V_15_reg_14998;
reg   [7:0] tmp_V_55_reg_15004;
reg   [7:0] tmp_V_52_reg_15010;
reg   [7:0] tmp_V_49_reg_15016;
reg   [7:0] tmp_2_2_V_15_reg_15022;
reg   [7:0] tmp_V_59_reg_15028;
reg   [7:0] tmp_V_56_reg_15034;
reg   [7:0] tmp_V_53_reg_15040;
reg   [7:0] tmp_V_50_reg_15046;
reg   [7:0] tmp_V_63_reg_15052;
reg   [7:0] tmp_V_60_reg_15058;
reg   [7:0] tmp_V_57_reg_15064;
reg   [7:0] tmp_V_54_reg_15070;
reg   [7:0] tmp_3_V_15_reg_15076;
reg   [7:0] tmp_V_64_reg_15242;
reg   [7:0] tmp_1_V_16_reg_15248;
reg   [7:0] tmp_2_1_V_16_reg_15254;
reg   [7:0] tmp_V_71_reg_15260;
reg   [7:0] tmp_V_68_reg_15266;
reg   [7:0] tmp_V_65_reg_15272;
reg   [7:0] tmp_2_2_V_16_reg_15278;
reg   [7:0] tmp_V_75_reg_15284;
reg   [7:0] tmp_V_72_reg_15290;
reg   [7:0] tmp_V_69_reg_15296;
reg   [7:0] tmp_V_66_reg_15302;
reg   [7:0] tmp_V_79_reg_15308;
reg   [7:0] tmp_V_76_reg_15314;
reg   [7:0] tmp_V_73_reg_15320;
reg   [7:0] tmp_V_70_reg_15326;
reg   [7:0] tmp_3_V_16_reg_15332;
reg   [7:0] tmp_V_80_reg_15498;
reg   [7:0] tmp_1_V_17_reg_15504;
reg   [7:0] tmp_2_1_V_17_reg_15510;
reg   [7:0] tmp_V_87_reg_15516;
reg   [7:0] tmp_V_84_reg_15522;
reg   [7:0] tmp_V_81_reg_15528;
reg   [7:0] tmp_2_2_V_17_reg_15534;
reg   [7:0] tmp_V_91_reg_15540;
reg   [7:0] tmp_V_88_reg_15546;
reg   [7:0] tmp_V_85_reg_15552;
reg   [7:0] tmp_V_82_reg_15558;
reg   [7:0] tmp_V_95_reg_15564;
reg   [7:0] tmp_V_92_reg_15570;
reg   [7:0] tmp_V_89_reg_15576;
reg   [7:0] tmp_V_86_reg_15582;
reg   [7:0] tmp_3_V_17_reg_15588;
reg   [7:0] tmp_V_96_reg_15754;
reg   [7:0] tmp_1_V_18_reg_15760;
reg   [7:0] tmp_2_1_V_18_reg_15766;
reg   [7:0] tmp_V_103_reg_15772;
reg   [7:0] tmp_V_100_reg_15778;
reg   [7:0] tmp_V_97_reg_15784;
reg   [7:0] tmp_2_2_V_18_reg_15790;
reg   [7:0] tmp_V_107_reg_15796;
reg   [7:0] tmp_V_104_reg_15802;
reg   [7:0] tmp_V_101_reg_15808;
reg   [7:0] tmp_V_98_reg_15814;
reg   [7:0] tmp_V_111_reg_15820;
reg   [7:0] tmp_V_108_reg_15826;
reg   [7:0] tmp_V_105_reg_15832;
reg   [7:0] tmp_V_102_reg_15838;
reg   [7:0] tmp_3_V_18_reg_15844;
reg   [7:0] tmp_V_112_reg_16010;
reg   [7:0] tmp_1_V_19_reg_16016;
reg   [7:0] tmp_2_1_V_19_reg_16022;
reg   [7:0] tmp_V_119_reg_16028;
reg   [7:0] tmp_V_116_reg_16034;
reg   [7:0] tmp_V_113_reg_16040;
reg   [7:0] tmp_2_2_V_19_reg_16046;
reg   [7:0] tmp_V_123_reg_16052;
reg   [7:0] tmp_V_120_reg_16058;
reg   [7:0] tmp_V_117_reg_16064;
reg   [7:0] tmp_V_114_reg_16070;
reg   [7:0] tmp_V_127_reg_16076;
reg   [7:0] tmp_V_124_reg_16082;
reg   [7:0] tmp_V_121_reg_16088;
reg   [7:0] tmp_V_118_reg_16094;
reg   [7:0] tmp_3_V_19_reg_16100;
reg   [7:0] tmp_V_128_reg_16266;
reg   [7:0] tmp_1_V_20_reg_16272;
reg   [7:0] tmp_2_1_V_20_reg_16278;
reg   [7:0] tmp_V_135_reg_16284;
reg   [7:0] tmp_V_132_reg_16290;
reg   [7:0] tmp_V_129_reg_16296;
reg   [7:0] tmp_2_2_V_20_reg_16302;
reg   [7:0] tmp_V_139_reg_16308;
reg   [7:0] tmp_V_136_reg_16314;
reg   [7:0] tmp_V_133_reg_16320;
reg   [7:0] tmp_V_130_reg_16326;
reg   [7:0] tmp_V_143_reg_16332;
reg   [7:0] tmp_V_140_reg_16338;
reg   [7:0] tmp_V_137_reg_16344;
reg   [7:0] tmp_V_134_reg_16350;
reg   [7:0] tmp_3_V_20_reg_16356;
reg   [7:0] tmp_V_144_reg_16522;
reg   [7:0] tmp_1_V_21_reg_16528;
reg   [7:0] tmp_2_1_V_21_reg_16534;
reg   [7:0] tmp_V_151_reg_16540;
reg   [7:0] tmp_V_148_reg_16546;
reg   [7:0] tmp_V_145_reg_16552;
reg   [7:0] tmp_2_2_V_21_reg_16558;
reg   [7:0] tmp_V_155_reg_16564;
reg   [7:0] tmp_V_152_reg_16570;
reg   [7:0] tmp_V_149_reg_16576;
reg   [7:0] tmp_V_146_reg_16582;
reg   [7:0] tmp_V_159_reg_16588;
reg   [7:0] tmp_V_156_reg_16594;
reg   [7:0] tmp_V_153_reg_16600;
reg   [7:0] tmp_V_150_reg_16606;
reg   [7:0] tmp_3_V_21_reg_16612;
reg   [7:0] tmp_V_160_reg_16778;
reg   [7:0] tmp_1_V_22_reg_16784;
reg   [7:0] tmp_2_1_V_22_reg_16790;
reg   [7:0] tmp_V_167_reg_16796;
reg   [7:0] tmp_V_164_reg_16802;
reg   [7:0] tmp_V_161_reg_16808;
reg   [7:0] tmp_2_2_V_22_reg_16814;
reg   [7:0] tmp_V_171_reg_16820;
reg   [7:0] tmp_V_168_reg_16826;
reg   [7:0] tmp_V_165_reg_16832;
reg   [7:0] tmp_V_162_reg_16838;
reg   [7:0] tmp_V_175_reg_16844;
reg   [7:0] tmp_V_172_reg_16850;
reg   [7:0] tmp_V_169_reg_16856;
reg   [7:0] tmp_V_166_reg_16862;
reg   [7:0] tmp_3_V_22_reg_16868;
wire   [63:0] zext_ln708_fu_4622_p1;
wire    ap_block_pp0_stage0;
wire   [63:0] zext_ln708_4_fu_4637_p1;
wire   [63:0] zext_ln708_5_fu_4652_p1;
wire   [63:0] zext_ln708_6_fu_4667_p1;
wire   [63:0] zext_ln708_7_fu_4682_p1;
wire   [63:0] zext_ln708_8_fu_4697_p1;
wire   [63:0] zext_ln708_9_fu_4712_p1;
wire   [63:0] zext_ln708_10_fu_4727_p1;
wire   [63:0] zext_ln708_11_fu_4742_p1;
wire   [63:0] zext_ln708_12_fu_4757_p1;
wire   [63:0] zext_ln708_13_fu_4772_p1;
wire   [63:0] zext_ln708_14_fu_4787_p1;
wire   [63:0] zext_ln708_15_fu_4802_p1;
wire   [63:0] zext_ln708_16_fu_4817_p1;
wire   [63:0] zext_ln708_17_fu_4832_p1;
wire   [63:0] zext_ln708_18_fu_4847_p1;
wire   [63:0] zext_ln587_fu_4852_p1;
wire   [63:0] zext_ln587_1_fu_4857_p1;
wire   [63:0] zext_ln587_2_fu_4862_p1;
wire   [63:0] zext_ln587_3_fu_4867_p1;
wire   [63:0] zext_ln587_4_fu_4872_p1;
wire   [63:0] zext_ln587_5_fu_4877_p1;
wire   [63:0] zext_ln587_6_fu_4882_p1;
wire   [63:0] zext_ln587_7_fu_4887_p1;
wire   [63:0] zext_ln587_8_fu_4892_p1;
wire   [63:0] zext_ln587_9_fu_4897_p1;
wire   [63:0] zext_ln587_10_fu_4902_p1;
wire   [63:0] zext_ln587_11_fu_4907_p1;
wire   [63:0] zext_ln587_12_fu_4912_p1;
wire   [63:0] zext_ln587_13_fu_4917_p1;
wire   [63:0] zext_ln587_14_fu_4922_p1;
wire   [63:0] zext_ln587_15_fu_4927_p1;
wire   [63:0] zext_ln708_19_fu_5457_p1;
wire   [63:0] zext_ln708_20_fu_5472_p1;
wire   [63:0] zext_ln708_21_fu_5487_p1;
wire   [63:0] zext_ln708_22_fu_5502_p1;
wire   [63:0] zext_ln708_23_fu_5517_p1;
wire   [63:0] zext_ln708_24_fu_5532_p1;
wire   [63:0] zext_ln708_25_fu_5547_p1;
wire   [63:0] zext_ln708_26_fu_5562_p1;
wire   [63:0] zext_ln708_27_fu_5577_p1;
wire   [63:0] zext_ln708_28_fu_5592_p1;
wire   [63:0] zext_ln708_29_fu_5607_p1;
wire   [63:0] zext_ln708_30_fu_5622_p1;
wire   [63:0] zext_ln708_31_fu_5637_p1;
wire   [63:0] zext_ln708_32_fu_5652_p1;
wire   [63:0] zext_ln708_33_fu_5667_p1;
wire   [63:0] zext_ln708_34_fu_5682_p1;
wire   [63:0] zext_ln587_16_fu_5687_p1;
wire   [63:0] zext_ln587_17_fu_5692_p1;
wire   [63:0] zext_ln587_18_fu_5697_p1;
wire   [63:0] zext_ln587_19_fu_5702_p1;
wire   [63:0] zext_ln587_20_fu_5707_p1;
wire   [63:0] zext_ln587_21_fu_5712_p1;
wire   [63:0] zext_ln587_22_fu_5717_p1;
wire   [63:0] zext_ln587_23_fu_5722_p1;
wire   [63:0] zext_ln587_24_fu_5727_p1;
wire   [63:0] zext_ln587_25_fu_5732_p1;
wire   [63:0] zext_ln587_26_fu_5737_p1;
wire   [63:0] zext_ln587_27_fu_5742_p1;
wire   [63:0] zext_ln587_28_fu_5747_p1;
wire   [63:0] zext_ln587_29_fu_5752_p1;
wire   [63:0] zext_ln587_30_fu_5757_p1;
wire   [63:0] zext_ln587_31_fu_5762_p1;
wire   [63:0] zext_ln708_35_fu_6292_p1;
wire   [63:0] zext_ln708_36_fu_6307_p1;
wire   [63:0] zext_ln708_37_fu_6322_p1;
wire   [63:0] zext_ln708_38_fu_6337_p1;
wire   [63:0] zext_ln708_39_fu_6352_p1;
wire   [63:0] zext_ln708_40_fu_6367_p1;
wire   [63:0] zext_ln708_41_fu_6382_p1;
wire   [63:0] zext_ln708_42_fu_6397_p1;
wire   [63:0] zext_ln708_43_fu_6412_p1;
wire   [63:0] zext_ln708_44_fu_6427_p1;
wire   [63:0] zext_ln708_45_fu_6442_p1;
wire   [63:0] zext_ln708_46_fu_6457_p1;
wire   [63:0] zext_ln708_47_fu_6472_p1;
wire   [63:0] zext_ln708_48_fu_6487_p1;
wire   [63:0] zext_ln708_49_fu_6502_p1;
wire   [63:0] zext_ln708_50_fu_6517_p1;
wire   [63:0] zext_ln587_32_fu_6522_p1;
wire   [63:0] zext_ln587_33_fu_6527_p1;
wire   [63:0] zext_ln587_34_fu_6532_p1;
wire   [63:0] zext_ln587_35_fu_6537_p1;
wire   [63:0] zext_ln587_36_fu_6542_p1;
wire   [63:0] zext_ln587_37_fu_6547_p1;
wire   [63:0] zext_ln587_38_fu_6552_p1;
wire   [63:0] zext_ln587_39_fu_6557_p1;
wire   [63:0] zext_ln587_40_fu_6562_p1;
wire   [63:0] zext_ln587_41_fu_6567_p1;
wire   [63:0] zext_ln587_42_fu_6572_p1;
wire   [63:0] zext_ln587_43_fu_6577_p1;
wire   [63:0] zext_ln587_44_fu_6582_p1;
wire   [63:0] zext_ln587_45_fu_6587_p1;
wire   [63:0] zext_ln587_46_fu_6592_p1;
wire   [63:0] zext_ln587_47_fu_6597_p1;
wire   [63:0] zext_ln708_51_fu_7127_p1;
wire   [63:0] zext_ln708_52_fu_7142_p1;
wire   [63:0] zext_ln708_53_fu_7157_p1;
wire   [63:0] zext_ln708_54_fu_7172_p1;
wire   [63:0] zext_ln708_55_fu_7187_p1;
wire   [63:0] zext_ln708_56_fu_7202_p1;
wire   [63:0] zext_ln708_57_fu_7217_p1;
wire   [63:0] zext_ln708_58_fu_7232_p1;
wire   [63:0] zext_ln708_59_fu_7247_p1;
wire   [63:0] zext_ln708_60_fu_7262_p1;
wire   [63:0] zext_ln708_61_fu_7277_p1;
wire   [63:0] zext_ln708_62_fu_7292_p1;
wire   [63:0] zext_ln708_63_fu_7307_p1;
wire   [63:0] zext_ln708_64_fu_7322_p1;
wire   [63:0] zext_ln708_65_fu_7337_p1;
wire   [63:0] zext_ln708_66_fu_7352_p1;
wire   [63:0] zext_ln587_48_fu_7357_p1;
wire   [63:0] zext_ln587_49_fu_7362_p1;
wire   [63:0] zext_ln587_50_fu_7367_p1;
wire   [63:0] zext_ln587_51_fu_7372_p1;
wire   [63:0] zext_ln587_52_fu_7377_p1;
wire   [63:0] zext_ln587_53_fu_7382_p1;
wire   [63:0] zext_ln587_54_fu_7387_p1;
wire   [63:0] zext_ln587_55_fu_7392_p1;
wire   [63:0] zext_ln587_56_fu_7397_p1;
wire   [63:0] zext_ln587_57_fu_7402_p1;
wire   [63:0] zext_ln587_58_fu_7407_p1;
wire   [63:0] zext_ln587_59_fu_7412_p1;
wire   [63:0] zext_ln587_60_fu_7417_p1;
wire   [63:0] zext_ln587_61_fu_7422_p1;
wire   [63:0] zext_ln587_62_fu_7427_p1;
wire   [63:0] zext_ln587_63_fu_7432_p1;
wire   [63:0] zext_ln708_67_fu_7962_p1;
wire   [63:0] zext_ln708_68_fu_7977_p1;
wire   [63:0] zext_ln708_69_fu_7992_p1;
wire   [63:0] zext_ln708_70_fu_8007_p1;
wire   [63:0] zext_ln708_71_fu_8022_p1;
wire   [63:0] zext_ln708_72_fu_8037_p1;
wire   [63:0] zext_ln708_73_fu_8052_p1;
wire   [63:0] zext_ln708_74_fu_8067_p1;
wire   [63:0] zext_ln708_75_fu_8082_p1;
wire   [63:0] zext_ln708_76_fu_8097_p1;
wire   [63:0] zext_ln708_77_fu_8112_p1;
wire   [63:0] zext_ln708_78_fu_8127_p1;
wire   [63:0] zext_ln708_79_fu_8142_p1;
wire   [63:0] zext_ln708_80_fu_8157_p1;
wire   [63:0] zext_ln708_81_fu_8172_p1;
wire   [63:0] zext_ln708_82_fu_8187_p1;
wire   [63:0] zext_ln587_64_fu_8192_p1;
wire   [63:0] zext_ln587_65_fu_8197_p1;
wire   [63:0] zext_ln587_66_fu_8202_p1;
wire   [63:0] zext_ln587_67_fu_8207_p1;
wire   [63:0] zext_ln587_68_fu_8212_p1;
wire   [63:0] zext_ln587_69_fu_8217_p1;
wire   [63:0] zext_ln587_70_fu_8222_p1;
wire   [63:0] zext_ln587_71_fu_8227_p1;
wire   [63:0] zext_ln587_72_fu_8232_p1;
wire   [63:0] zext_ln587_73_fu_8237_p1;
wire   [63:0] zext_ln587_74_fu_8242_p1;
wire   [63:0] zext_ln587_75_fu_8247_p1;
wire   [63:0] zext_ln587_76_fu_8252_p1;
wire   [63:0] zext_ln587_77_fu_8257_p1;
wire   [63:0] zext_ln587_78_fu_8262_p1;
wire   [63:0] zext_ln587_79_fu_8267_p1;
wire   [63:0] zext_ln708_83_fu_8797_p1;
wire   [63:0] zext_ln708_84_fu_8812_p1;
wire   [63:0] zext_ln708_85_fu_8827_p1;
wire   [63:0] zext_ln708_86_fu_8842_p1;
wire   [63:0] zext_ln708_87_fu_8857_p1;
wire   [63:0] zext_ln708_88_fu_8872_p1;
wire   [63:0] zext_ln708_89_fu_8887_p1;
wire   [63:0] zext_ln708_90_fu_8902_p1;
wire   [63:0] zext_ln708_91_fu_8917_p1;
wire   [63:0] zext_ln708_92_fu_8932_p1;
wire   [63:0] zext_ln708_93_fu_8947_p1;
wire   [63:0] zext_ln708_94_fu_8962_p1;
wire   [63:0] zext_ln708_95_fu_8977_p1;
wire   [63:0] zext_ln708_96_fu_8992_p1;
wire   [63:0] zext_ln708_97_fu_9007_p1;
wire   [63:0] zext_ln708_98_fu_9022_p1;
wire   [63:0] zext_ln587_80_fu_9027_p1;
wire   [63:0] zext_ln587_81_fu_9032_p1;
wire   [63:0] zext_ln587_82_fu_9037_p1;
wire   [63:0] zext_ln587_83_fu_9042_p1;
wire   [63:0] zext_ln587_84_fu_9047_p1;
wire   [63:0] zext_ln587_85_fu_9052_p1;
wire   [63:0] zext_ln587_86_fu_9057_p1;
wire   [63:0] zext_ln587_87_fu_9062_p1;
wire   [63:0] zext_ln587_88_fu_9067_p1;
wire   [63:0] zext_ln587_89_fu_9072_p1;
wire   [63:0] zext_ln587_90_fu_9077_p1;
wire   [63:0] zext_ln587_91_fu_9082_p1;
wire   [63:0] zext_ln587_92_fu_9087_p1;
wire   [63:0] zext_ln587_93_fu_9092_p1;
wire   [63:0] zext_ln587_94_fu_9097_p1;
wire   [63:0] zext_ln587_95_fu_9102_p1;
wire   [63:0] zext_ln708_99_fu_9632_p1;
wire   [63:0] zext_ln708_100_fu_9647_p1;
wire   [63:0] zext_ln708_101_fu_9662_p1;
wire   [63:0] zext_ln708_102_fu_9677_p1;
wire   [63:0] zext_ln708_103_fu_9692_p1;
wire   [63:0] zext_ln708_104_fu_9707_p1;
wire   [63:0] zext_ln708_105_fu_9722_p1;
wire   [63:0] zext_ln708_106_fu_9737_p1;
wire   [63:0] zext_ln708_107_fu_9752_p1;
wire   [63:0] zext_ln708_108_fu_9767_p1;
wire   [63:0] zext_ln708_109_fu_9782_p1;
wire   [63:0] zext_ln708_110_fu_9797_p1;
wire   [63:0] zext_ln708_111_fu_9812_p1;
wire   [63:0] zext_ln708_112_fu_9827_p1;
wire   [63:0] zext_ln708_113_fu_9842_p1;
wire   [63:0] zext_ln708_114_fu_9857_p1;
wire   [63:0] zext_ln587_96_fu_9862_p1;
wire   [63:0] zext_ln587_97_fu_9867_p1;
wire   [63:0] zext_ln587_98_fu_9872_p1;
wire   [63:0] zext_ln587_99_fu_9877_p1;
wire   [63:0] zext_ln587_100_fu_9882_p1;
wire   [63:0] zext_ln587_101_fu_9887_p1;
wire   [63:0] zext_ln587_102_fu_9892_p1;
wire   [63:0] zext_ln587_103_fu_9897_p1;
wire   [63:0] zext_ln587_104_fu_9902_p1;
wire   [63:0] zext_ln587_105_fu_9907_p1;
wire   [63:0] zext_ln587_106_fu_9912_p1;
wire   [63:0] zext_ln587_107_fu_9917_p1;
wire   [63:0] zext_ln587_108_fu_9922_p1;
wire   [63:0] zext_ln587_109_fu_9927_p1;
wire   [63:0] zext_ln587_110_fu_9932_p1;
wire   [63:0] zext_ln587_111_fu_9937_p1;
wire   [63:0] zext_ln708_115_fu_10467_p1;
wire   [63:0] zext_ln708_116_fu_10482_p1;
wire   [63:0] zext_ln708_117_fu_10497_p1;
wire   [63:0] zext_ln708_118_fu_10512_p1;
wire   [63:0] zext_ln708_119_fu_10527_p1;
wire   [63:0] zext_ln708_120_fu_10542_p1;
wire   [63:0] zext_ln708_121_fu_10557_p1;
wire   [63:0] zext_ln708_122_fu_10572_p1;
wire   [63:0] zext_ln708_123_fu_10587_p1;
wire   [63:0] zext_ln708_124_fu_10602_p1;
wire   [63:0] zext_ln708_125_fu_10617_p1;
wire   [63:0] zext_ln708_126_fu_10632_p1;
wire   [63:0] zext_ln708_127_fu_10647_p1;
wire   [63:0] zext_ln708_128_fu_10662_p1;
wire   [63:0] zext_ln708_129_fu_10677_p1;
wire   [63:0] zext_ln708_130_fu_10692_p1;
wire   [63:0] zext_ln587_112_fu_10697_p1;
wire   [63:0] zext_ln587_113_fu_10702_p1;
wire   [63:0] zext_ln587_114_fu_10707_p1;
wire   [63:0] zext_ln587_115_fu_10712_p1;
wire   [63:0] zext_ln587_116_fu_10717_p1;
wire   [63:0] zext_ln587_117_fu_10722_p1;
wire   [63:0] zext_ln587_118_fu_10727_p1;
wire   [63:0] zext_ln587_119_fu_10732_p1;
wire   [63:0] zext_ln587_120_fu_10737_p1;
wire   [63:0] zext_ln587_121_fu_10742_p1;
wire   [63:0] zext_ln587_122_fu_10747_p1;
wire   [63:0] zext_ln587_123_fu_10752_p1;
wire   [63:0] zext_ln587_124_fu_10757_p1;
wire   [63:0] zext_ln587_125_fu_10762_p1;
wire   [63:0] zext_ln587_126_fu_10767_p1;
wire   [63:0] zext_ln587_127_fu_10772_p1;
wire   [63:0] zext_ln708_131_fu_11302_p1;
wire   [63:0] zext_ln708_132_fu_11317_p1;
wire   [63:0] zext_ln708_133_fu_11332_p1;
wire   [63:0] zext_ln708_134_fu_11347_p1;
wire   [63:0] zext_ln708_135_fu_11362_p1;
wire   [63:0] zext_ln708_136_fu_11377_p1;
wire   [63:0] zext_ln708_137_fu_11392_p1;
wire   [63:0] zext_ln708_138_fu_11407_p1;
wire   [63:0] zext_ln708_139_fu_11422_p1;
wire   [63:0] zext_ln708_140_fu_11437_p1;
wire   [63:0] zext_ln708_141_fu_11452_p1;
wire   [63:0] zext_ln708_142_fu_11467_p1;
wire   [63:0] zext_ln708_143_fu_11482_p1;
wire   [63:0] zext_ln708_144_fu_11497_p1;
wire   [63:0] zext_ln708_145_fu_11512_p1;
wire   [63:0] zext_ln708_146_fu_11527_p1;
wire   [63:0] zext_ln587_128_fu_11532_p1;
wire   [63:0] zext_ln587_129_fu_11537_p1;
wire   [63:0] zext_ln587_130_fu_11542_p1;
wire   [63:0] zext_ln587_131_fu_11547_p1;
wire   [63:0] zext_ln587_132_fu_11552_p1;
wire   [63:0] zext_ln587_133_fu_11557_p1;
wire   [63:0] zext_ln587_134_fu_11562_p1;
wire   [63:0] zext_ln587_135_fu_11567_p1;
wire   [63:0] zext_ln587_136_fu_11572_p1;
wire   [63:0] zext_ln587_137_fu_11577_p1;
wire   [63:0] zext_ln587_138_fu_11582_p1;
wire   [63:0] zext_ln587_139_fu_11587_p1;
wire   [63:0] zext_ln587_140_fu_11592_p1;
wire   [63:0] zext_ln587_141_fu_11597_p1;
wire   [63:0] zext_ln587_142_fu_11602_p1;
wire   [63:0] zext_ln587_143_fu_11607_p1;
wire   [63:0] zext_ln708_147_fu_12137_p1;
wire   [63:0] zext_ln708_148_fu_12152_p1;
wire   [63:0] zext_ln708_149_fu_12167_p1;
wire   [63:0] zext_ln708_150_fu_12182_p1;
wire   [63:0] zext_ln708_151_fu_12197_p1;
wire   [63:0] zext_ln708_152_fu_12212_p1;
wire   [63:0] zext_ln708_153_fu_12227_p1;
wire   [63:0] zext_ln708_154_fu_12242_p1;
wire   [63:0] zext_ln708_155_fu_12257_p1;
wire   [63:0] zext_ln708_156_fu_12272_p1;
wire   [63:0] zext_ln708_157_fu_12287_p1;
wire   [63:0] zext_ln708_158_fu_12302_p1;
wire   [63:0] zext_ln708_159_fu_12317_p1;
wire   [63:0] zext_ln708_160_fu_12332_p1;
wire   [63:0] zext_ln708_161_fu_12347_p1;
wire   [63:0] zext_ln708_162_fu_12362_p1;
wire   [63:0] zext_ln587_144_fu_12367_p1;
wire   [63:0] zext_ln587_145_fu_12372_p1;
wire   [63:0] zext_ln587_146_fu_12377_p1;
wire   [63:0] zext_ln587_147_fu_12382_p1;
wire   [63:0] zext_ln587_148_fu_12387_p1;
wire   [63:0] zext_ln587_149_fu_12392_p1;
wire   [63:0] zext_ln587_150_fu_12397_p1;
wire   [63:0] zext_ln587_151_fu_12402_p1;
wire   [63:0] zext_ln587_152_fu_12407_p1;
wire   [63:0] zext_ln587_153_fu_12412_p1;
wire   [63:0] zext_ln587_154_fu_12417_p1;
wire   [63:0] zext_ln587_155_fu_12422_p1;
wire   [63:0] zext_ln587_156_fu_12427_p1;
wire   [63:0] zext_ln587_157_fu_12432_p1;
wire   [63:0] zext_ln587_158_fu_12437_p1;
wire   [63:0] zext_ln587_159_fu_12442_p1;
wire   [63:0] zext_ln708_163_fu_12972_p1;
wire   [63:0] zext_ln708_164_fu_12987_p1;
wire   [63:0] zext_ln708_165_fu_13002_p1;
wire   [63:0] zext_ln708_166_fu_13017_p1;
wire   [63:0] zext_ln708_167_fu_13032_p1;
wire   [63:0] zext_ln708_168_fu_13047_p1;
wire   [63:0] zext_ln708_169_fu_13062_p1;
wire   [63:0] zext_ln708_170_fu_13077_p1;
wire   [63:0] zext_ln708_171_fu_13092_p1;
wire   [63:0] zext_ln708_172_fu_13107_p1;
wire   [63:0] zext_ln708_173_fu_13122_p1;
wire   [63:0] zext_ln708_174_fu_13137_p1;
wire   [63:0] zext_ln708_175_fu_13152_p1;
wire   [63:0] zext_ln708_176_fu_13167_p1;
wire   [63:0] zext_ln708_177_fu_13182_p1;
wire   [63:0] zext_ln708_178_fu_13197_p1;
wire   [63:0] zext_ln587_160_fu_13202_p1;
wire   [63:0] zext_ln587_161_fu_13207_p1;
wire   [63:0] zext_ln587_162_fu_13212_p1;
wire   [63:0] zext_ln587_163_fu_13217_p1;
wire   [63:0] zext_ln587_164_fu_13222_p1;
wire   [63:0] zext_ln587_165_fu_13227_p1;
wire   [63:0] zext_ln587_166_fu_13232_p1;
wire   [63:0] zext_ln587_167_fu_13237_p1;
wire   [63:0] zext_ln587_168_fu_13242_p1;
wire   [63:0] zext_ln587_169_fu_13247_p1;
wire   [63:0] zext_ln587_170_fu_13252_p1;
wire   [63:0] zext_ln587_171_fu_13257_p1;
wire   [63:0] zext_ln587_172_fu_13262_p1;
wire   [63:0] zext_ln587_173_fu_13267_p1;
wire   [63:0] zext_ln587_174_fu_13272_p1;
wire   [63:0] zext_ln587_175_fu_13277_p1;
wire   [63:0] zext_ln708_179_fu_13807_p1;
wire   [63:0] zext_ln708_180_fu_13822_p1;
wire   [63:0] zext_ln708_181_fu_13837_p1;
wire   [63:0] zext_ln708_182_fu_13852_p1;
wire   [63:0] zext_ln708_183_fu_13867_p1;
wire   [63:0] zext_ln708_184_fu_13882_p1;
wire   [63:0] zext_ln708_185_fu_13897_p1;
wire   [63:0] zext_ln708_186_fu_13912_p1;
wire   [63:0] zext_ln708_187_fu_13927_p1;
wire   [63:0] zext_ln708_188_fu_13942_p1;
wire   [63:0] zext_ln708_189_fu_13957_p1;
wire   [63:0] zext_ln708_190_fu_13972_p1;
wire   [63:0] zext_ln708_191_fu_13987_p1;
wire   [63:0] zext_ln708_192_fu_14002_p1;
wire   [63:0] zext_ln708_193_fu_14017_p1;
wire   [63:0] zext_ln708_194_fu_14032_p1;
wire   [127:0] ret_V_fu_4612_p2;
wire   [7:0] trunc_ln708_fu_4618_p1;
wire   [7:0] tmp_s_fu_4627_p4;
wire   [7:0] tmp_14_fu_4642_p4;
wire   [7:0] tmp_15_fu_4657_p4;
wire   [7:0] tmp_16_fu_4672_p4;
wire   [7:0] tmp_17_fu_4687_p4;
wire   [7:0] tmp_18_fu_4702_p4;
wire   [7:0] tmp_19_fu_4717_p4;
wire   [7:0] tmp_20_fu_4732_p4;
wire   [7:0] tmp_21_fu_4747_p4;
wire   [7:0] tmp_22_fu_4762_p4;
wire   [7:0] tmp_23_fu_4777_p4;
wire   [7:0] tmp_24_fu_4792_p4;
wire   [7:0] tmp_25_fu_4807_p4;
wire   [7:0] tmp_26_fu_4822_p4;
wire   [7:0] tmp_27_fu_4837_p4;
wire   [7:0] tmp_29_fu_4950_p4;
wire   [7:0] trunc_ln674_fu_4932_p1;
wire   [7:0] xor_ln1545_8_fu_5160_p2;
wire   [7:0] xor_ln1545_fu_5156_p2;
wire   [7:0] trunc_ln674_2_fu_4946_p1;
wire   [7:0] tmp_30_fu_4964_p4;
wire   [7:0] xor_ln1545_11_fu_5176_p2;
wire   [7:0] xor_ln1545_9_fu_5172_p2;
wire   [7:0] trunc_ln674_3_fu_4960_p1;
wire   [7:0] tmp_31_fu_4978_p4;
wire   [7:0] xor_ln1545_14_fu_5192_p2;
wire   [7:0] xor_ln1545_12_fu_5188_p2;
wire   [7:0] tmp_28_fu_4936_p4;
wire   [7:0] trunc_ln674_4_fu_4974_p1;
wire   [7:0] xor_ln1545_17_fu_5208_p2;
wire   [7:0] xor_ln1545_15_fu_5204_p2;
wire   [7:0] tmp_33_fu_5006_p4;
wire   [7:0] trunc_ln674_5_fu_4988_p1;
wire   [7:0] xor_ln1545_20_fu_5224_p2;
wire   [7:0] xor_ln1545_18_fu_5220_p2;
wire   [7:0] trunc_ln674_6_fu_5002_p1;
wire   [7:0] tmp_34_fu_5020_p4;
wire   [7:0] xor_ln1545_23_fu_5240_p2;
wire   [7:0] xor_ln1545_21_fu_5236_p2;
wire   [7:0] trunc_ln674_7_fu_5016_p1;
wire   [7:0] tmp_35_fu_5034_p4;
wire   [7:0] xor_ln1545_26_fu_5256_p2;
wire   [7:0] xor_ln1545_24_fu_5252_p2;
wire   [7:0] tmp_32_fu_4992_p4;
wire   [7:0] trunc_ln674_8_fu_5030_p1;
wire   [7:0] xor_ln1545_29_fu_5272_p2;
wire   [7:0] xor_ln1545_27_fu_5268_p2;
wire   [7:0] tmp_37_fu_5062_p4;
wire   [7:0] trunc_ln674_9_fu_5044_p1;
wire   [7:0] xor_ln1545_32_fu_5288_p2;
wire   [7:0] xor_ln1545_30_fu_5284_p2;
wire   [7:0] trunc_ln674_10_fu_5058_p1;
wire   [7:0] tmp_38_fu_5076_p4;
wire   [7:0] xor_ln1545_35_fu_5304_p2;
wire   [7:0] xor_ln1545_33_fu_5300_p2;
wire   [7:0] trunc_ln674_11_fu_5072_p1;
wire   [7:0] tmp_39_fu_5090_p4;
wire   [7:0] xor_ln1545_38_fu_5320_p2;
wire   [7:0] xor_ln1545_36_fu_5316_p2;
wire   [7:0] tmp_36_fu_5048_p4;
wire   [7:0] trunc_ln674_12_fu_5086_p1;
wire   [7:0] xor_ln1545_41_fu_5336_p2;
wire   [7:0] xor_ln1545_39_fu_5332_p2;
wire   [7:0] tmp_41_fu_5118_p4;
wire   [7:0] trunc_ln674_13_fu_5100_p1;
wire   [7:0] xor_ln1545_44_fu_5352_p2;
wire   [7:0] xor_ln1545_42_fu_5348_p2;
wire   [7:0] trunc_ln674_14_fu_5114_p1;
wire   [7:0] tmp_42_fu_5132_p4;
wire   [7:0] xor_ln1545_47_fu_5368_p2;
wire   [7:0] xor_ln1545_45_fu_5364_p2;
wire   [7:0] trunc_ln674_15_fu_5128_p1;
wire   [7:0] tmp_43_fu_5146_p4;
wire   [7:0] xor_ln1545_50_fu_5384_p2;
wire   [7:0] xor_ln1545_48_fu_5380_p2;
wire   [7:0] tmp_40_fu_5104_p4;
wire   [7:0] trunc_ln674_16_fu_5142_p1;
wire   [7:0] xor_ln1545_53_fu_5400_p2;
wire   [7:0] xor_ln1545_51_fu_5396_p2;
wire   [7:0] xor_ln1545_52_fu_5406_p2;
wire   [7:0] xor_ln1545_49_fu_5390_p2;
wire   [7:0] xor_ln1545_46_fu_5374_p2;
wire   [7:0] xor_ln1545_43_fu_5358_p2;
wire   [7:0] xor_ln1545_40_fu_5342_p2;
wire   [7:0] xor_ln1545_37_fu_5326_p2;
wire   [7:0] xor_ln1545_34_fu_5310_p2;
wire   [7:0] xor_ln1545_31_fu_5294_p2;
wire   [7:0] xor_ln1545_28_fu_5278_p2;
wire   [7:0] xor_ln1545_25_fu_5262_p2;
wire   [7:0] xor_ln1545_22_fu_5246_p2;
wire   [7:0] xor_ln1545_19_fu_5230_p2;
wire   [7:0] xor_ln1545_16_fu_5214_p2;
wire   [7:0] xor_ln1545_13_fu_5198_p2;
wire   [7:0] xor_ln1545_10_fu_5182_p2;
wire   [7:0] xor_ln1545_7_fu_5166_p2;
wire   [127:0] p_Result_s_fu_5412_p17;
wire   [127:0] state_V_24_fu_5448_p2;
wire   [7:0] trunc_ln708_1_fu_5453_p1;
wire   [7:0] tmp_44_fu_5462_p4;
wire   [7:0] tmp_45_fu_5477_p4;
wire   [7:0] tmp_46_fu_5492_p4;
wire   [7:0] tmp_47_fu_5507_p4;
wire   [7:0] tmp_48_fu_5522_p4;
wire   [7:0] tmp_49_fu_5537_p4;
wire   [7:0] tmp_50_fu_5552_p4;
wire   [7:0] tmp_51_fu_5567_p4;
wire   [7:0] tmp_52_fu_5582_p4;
wire   [7:0] tmp_53_fu_5597_p4;
wire   [7:0] tmp_54_fu_5612_p4;
wire   [7:0] tmp_55_fu_5627_p4;
wire   [7:0] tmp_56_fu_5642_p4;
wire   [7:0] tmp_57_fu_5657_p4;
wire   [7:0] tmp_58_fu_5672_p4;
wire   [7:0] tmp_60_fu_5785_p4;
wire   [7:0] trunc_ln674_17_fu_5767_p1;
wire   [7:0] xor_ln1545_56_fu_5995_p2;
wire   [7:0] xor_ln1545_54_fu_5991_p2;
wire   [7:0] trunc_ln674_18_fu_5781_p1;
wire   [7:0] tmp_61_fu_5799_p4;
wire   [7:0] xor_ln1545_59_fu_6011_p2;
wire   [7:0] xor_ln1545_57_fu_6007_p2;
wire   [7:0] trunc_ln674_19_fu_5795_p1;
wire   [7:0] tmp_62_fu_5813_p4;
wire   [7:0] xor_ln1545_62_fu_6027_p2;
wire   [7:0] xor_ln1545_60_fu_6023_p2;
wire   [7:0] tmp_59_fu_5771_p4;
wire   [7:0] trunc_ln674_20_fu_5809_p1;
wire   [7:0] xor_ln1545_65_fu_6043_p2;
wire   [7:0] xor_ln1545_63_fu_6039_p2;
wire   [7:0] tmp_64_fu_5841_p4;
wire   [7:0] trunc_ln674_21_fu_5823_p1;
wire   [7:0] xor_ln1545_68_fu_6059_p2;
wire   [7:0] xor_ln1545_66_fu_6055_p2;
wire   [7:0] trunc_ln674_22_fu_5837_p1;
wire   [7:0] tmp_65_fu_5855_p4;
wire   [7:0] xor_ln1545_71_fu_6075_p2;
wire   [7:0] xor_ln1545_69_fu_6071_p2;
wire   [7:0] trunc_ln674_23_fu_5851_p1;
wire   [7:0] tmp_66_fu_5869_p4;
wire   [7:0] xor_ln1545_74_fu_6091_p2;
wire   [7:0] xor_ln1545_72_fu_6087_p2;
wire   [7:0] tmp_63_fu_5827_p4;
wire   [7:0] trunc_ln674_24_fu_5865_p1;
wire   [7:0] xor_ln1545_77_fu_6107_p2;
wire   [7:0] xor_ln1545_75_fu_6103_p2;
wire   [7:0] tmp_68_fu_5897_p4;
wire   [7:0] trunc_ln674_25_fu_5879_p1;
wire   [7:0] xor_ln1545_80_fu_6123_p2;
wire   [7:0] xor_ln1545_78_fu_6119_p2;
wire   [7:0] trunc_ln674_26_fu_5893_p1;
wire   [7:0] tmp_69_fu_5911_p4;
wire   [7:0] xor_ln1545_83_fu_6139_p2;
wire   [7:0] xor_ln1545_81_fu_6135_p2;
wire   [7:0] trunc_ln674_27_fu_5907_p1;
wire   [7:0] tmp_70_fu_5925_p4;
wire   [7:0] xor_ln1545_86_fu_6155_p2;
wire   [7:0] xor_ln1545_84_fu_6151_p2;
wire   [7:0] tmp_67_fu_5883_p4;
wire   [7:0] trunc_ln674_28_fu_5921_p1;
wire   [7:0] xor_ln1545_89_fu_6171_p2;
wire   [7:0] xor_ln1545_87_fu_6167_p2;
wire   [7:0] tmp_72_fu_5953_p4;
wire   [7:0] trunc_ln674_29_fu_5935_p1;
wire   [7:0] xor_ln1545_92_fu_6187_p2;
wire   [7:0] xor_ln1545_90_fu_6183_p2;
wire   [7:0] trunc_ln674_30_fu_5949_p1;
wire   [7:0] tmp_73_fu_5967_p4;
wire   [7:0] xor_ln1545_95_fu_6203_p2;
wire   [7:0] xor_ln1545_93_fu_6199_p2;
wire   [7:0] trunc_ln674_31_fu_5963_p1;
wire   [7:0] tmp_74_fu_5981_p4;
wire   [7:0] xor_ln1545_98_fu_6219_p2;
wire   [7:0] xor_ln1545_96_fu_6215_p2;
wire   [7:0] tmp_71_fu_5939_p4;
wire   [7:0] trunc_ln674_32_fu_5977_p1;
wire   [7:0] xor_ln1545_101_fu_6235_p2;
wire   [7:0] xor_ln1545_99_fu_6231_p2;
wire   [7:0] xor_ln1545_100_fu_6241_p2;
wire   [7:0] xor_ln1545_97_fu_6225_p2;
wire   [7:0] xor_ln1545_94_fu_6209_p2;
wire   [7:0] xor_ln1545_91_fu_6193_p2;
wire   [7:0] xor_ln1545_88_fu_6177_p2;
wire   [7:0] xor_ln1545_85_fu_6161_p2;
wire   [7:0] xor_ln1545_82_fu_6145_p2;
wire   [7:0] xor_ln1545_79_fu_6129_p2;
wire   [7:0] xor_ln1545_76_fu_6113_p2;
wire   [7:0] xor_ln1545_73_fu_6097_p2;
wire   [7:0] xor_ln1545_70_fu_6081_p2;
wire   [7:0] xor_ln1545_67_fu_6065_p2;
wire   [7:0] xor_ln1545_64_fu_6049_p2;
wire   [7:0] xor_ln1545_61_fu_6033_p2;
wire   [7:0] xor_ln1545_58_fu_6017_p2;
wire   [7:0] xor_ln1545_55_fu_6001_p2;
wire   [127:0] p_Result_25_fu_6247_p17;
wire   [127:0] state_V_25_fu_6283_p2;
wire   [7:0] trunc_ln708_2_fu_6288_p1;
wire   [7:0] tmp_75_fu_6297_p4;
wire   [7:0] tmp_76_fu_6312_p4;
wire   [7:0] tmp_77_fu_6327_p4;
wire   [7:0] tmp_78_fu_6342_p4;
wire   [7:0] tmp_79_fu_6357_p4;
wire   [7:0] tmp_80_fu_6372_p4;
wire   [7:0] tmp_81_fu_6387_p4;
wire   [7:0] tmp_82_fu_6402_p4;
wire   [7:0] tmp_83_fu_6417_p4;
wire   [7:0] tmp_84_fu_6432_p4;
wire   [7:0] tmp_85_fu_6447_p4;
wire   [7:0] tmp_86_fu_6462_p4;
wire   [7:0] tmp_87_fu_6477_p4;
wire   [7:0] tmp_88_fu_6492_p4;
wire   [7:0] tmp_89_fu_6507_p4;
wire   [7:0] tmp_91_fu_6620_p4;
wire   [7:0] trunc_ln674_33_fu_6602_p1;
wire   [7:0] xor_ln1545_104_fu_6830_p2;
wire   [7:0] xor_ln1545_102_fu_6826_p2;
wire   [7:0] trunc_ln674_34_fu_6616_p1;
wire   [7:0] tmp_92_fu_6634_p4;
wire   [7:0] xor_ln1545_107_fu_6846_p2;
wire   [7:0] xor_ln1545_105_fu_6842_p2;
wire   [7:0] trunc_ln674_35_fu_6630_p1;
wire   [7:0] tmp_93_fu_6648_p4;
wire   [7:0] xor_ln1545_110_fu_6862_p2;
wire   [7:0] xor_ln1545_108_fu_6858_p2;
wire   [7:0] tmp_90_fu_6606_p4;
wire   [7:0] trunc_ln674_36_fu_6644_p1;
wire   [7:0] xor_ln1545_113_fu_6878_p2;
wire   [7:0] xor_ln1545_111_fu_6874_p2;
wire   [7:0] tmp_95_fu_6676_p4;
wire   [7:0] trunc_ln674_37_fu_6658_p1;
wire   [7:0] xor_ln1545_116_fu_6894_p2;
wire   [7:0] xor_ln1545_114_fu_6890_p2;
wire   [7:0] trunc_ln674_38_fu_6672_p1;
wire   [7:0] tmp_96_fu_6690_p4;
wire   [7:0] xor_ln1545_119_fu_6910_p2;
wire   [7:0] xor_ln1545_117_fu_6906_p2;
wire   [7:0] trunc_ln674_39_fu_6686_p1;
wire   [7:0] tmp_97_fu_6704_p4;
wire   [7:0] xor_ln1545_122_fu_6926_p2;
wire   [7:0] xor_ln1545_120_fu_6922_p2;
wire   [7:0] tmp_94_fu_6662_p4;
wire   [7:0] trunc_ln674_40_fu_6700_p1;
wire   [7:0] xor_ln1545_125_fu_6942_p2;
wire   [7:0] xor_ln1545_123_fu_6938_p2;
wire   [7:0] tmp_99_fu_6732_p4;
wire   [7:0] trunc_ln674_41_fu_6714_p1;
wire   [7:0] xor_ln1545_128_fu_6958_p2;
wire   [7:0] xor_ln1545_126_fu_6954_p2;
wire   [7:0] trunc_ln674_42_fu_6728_p1;
wire   [7:0] tmp_100_fu_6746_p4;
wire   [7:0] xor_ln1545_131_fu_6974_p2;
wire   [7:0] xor_ln1545_129_fu_6970_p2;
wire   [7:0] trunc_ln674_43_fu_6742_p1;
wire   [7:0] tmp_101_fu_6760_p4;
wire   [7:0] xor_ln1545_134_fu_6990_p2;
wire   [7:0] xor_ln1545_132_fu_6986_p2;
wire   [7:0] tmp_98_fu_6718_p4;
wire   [7:0] trunc_ln674_44_fu_6756_p1;
wire   [7:0] xor_ln1545_137_fu_7006_p2;
wire   [7:0] xor_ln1545_135_fu_7002_p2;
wire   [7:0] tmp_103_fu_6788_p4;
wire   [7:0] trunc_ln674_45_fu_6770_p1;
wire   [7:0] xor_ln1545_140_fu_7022_p2;
wire   [7:0] xor_ln1545_138_fu_7018_p2;
wire   [7:0] trunc_ln674_46_fu_6784_p1;
wire   [7:0] tmp_104_fu_6802_p4;
wire   [7:0] xor_ln1545_143_fu_7038_p2;
wire   [7:0] xor_ln1545_141_fu_7034_p2;
wire   [7:0] trunc_ln674_47_fu_6798_p1;
wire   [7:0] tmp_105_fu_6816_p4;
wire   [7:0] xor_ln1545_146_fu_7054_p2;
wire   [7:0] xor_ln1545_144_fu_7050_p2;
wire   [7:0] tmp_102_fu_6774_p4;
wire   [7:0] trunc_ln674_48_fu_6812_p1;
wire   [7:0] xor_ln1545_149_fu_7070_p2;
wire   [7:0] xor_ln1545_147_fu_7066_p2;
wire   [7:0] xor_ln1545_148_fu_7076_p2;
wire   [7:0] xor_ln1545_145_fu_7060_p2;
wire   [7:0] xor_ln1545_142_fu_7044_p2;
wire   [7:0] xor_ln1545_139_fu_7028_p2;
wire   [7:0] xor_ln1545_136_fu_7012_p2;
wire   [7:0] xor_ln1545_133_fu_6996_p2;
wire   [7:0] xor_ln1545_130_fu_6980_p2;
wire   [7:0] xor_ln1545_127_fu_6964_p2;
wire   [7:0] xor_ln1545_124_fu_6948_p2;
wire   [7:0] xor_ln1545_121_fu_6932_p2;
wire   [7:0] xor_ln1545_118_fu_6916_p2;
wire   [7:0] xor_ln1545_115_fu_6900_p2;
wire   [7:0] xor_ln1545_112_fu_6884_p2;
wire   [7:0] xor_ln1545_109_fu_6868_p2;
wire   [7:0] xor_ln1545_106_fu_6852_p2;
wire   [7:0] xor_ln1545_103_fu_6836_p2;
wire   [127:0] p_Result_26_fu_7082_p17;
wire   [127:0] state_V_26_fu_7118_p2;
wire   [7:0] trunc_ln708_3_fu_7123_p1;
wire   [7:0] tmp_106_fu_7132_p4;
wire   [7:0] tmp_107_fu_7147_p4;
wire   [7:0] tmp_108_fu_7162_p4;
wire   [7:0] tmp_109_fu_7177_p4;
wire   [7:0] tmp_110_fu_7192_p4;
wire   [7:0] tmp_111_fu_7207_p4;
wire   [7:0] tmp_112_fu_7222_p4;
wire   [7:0] tmp_113_fu_7237_p4;
wire   [7:0] tmp_114_fu_7252_p4;
wire   [7:0] tmp_115_fu_7267_p4;
wire   [7:0] tmp_116_fu_7282_p4;
wire   [7:0] tmp_117_fu_7297_p4;
wire   [7:0] tmp_118_fu_7312_p4;
wire   [7:0] tmp_119_fu_7327_p4;
wire   [7:0] tmp_120_fu_7342_p4;
wire   [7:0] tmp_122_fu_7455_p4;
wire   [7:0] trunc_ln674_49_fu_7437_p1;
wire   [7:0] xor_ln1545_152_fu_7665_p2;
wire   [7:0] xor_ln1545_150_fu_7661_p2;
wire   [7:0] trunc_ln674_50_fu_7451_p1;
wire   [7:0] tmp_123_fu_7469_p4;
wire   [7:0] xor_ln1545_155_fu_7681_p2;
wire   [7:0] xor_ln1545_153_fu_7677_p2;
wire   [7:0] trunc_ln674_51_fu_7465_p1;
wire   [7:0] tmp_124_fu_7483_p4;
wire   [7:0] xor_ln1545_158_fu_7697_p2;
wire   [7:0] xor_ln1545_156_fu_7693_p2;
wire   [7:0] tmp_121_fu_7441_p4;
wire   [7:0] trunc_ln674_52_fu_7479_p1;
wire   [7:0] xor_ln1545_161_fu_7713_p2;
wire   [7:0] xor_ln1545_159_fu_7709_p2;
wire   [7:0] tmp_126_fu_7511_p4;
wire   [7:0] trunc_ln674_53_fu_7493_p1;
wire   [7:0] xor_ln1545_164_fu_7729_p2;
wire   [7:0] xor_ln1545_162_fu_7725_p2;
wire   [7:0] trunc_ln674_54_fu_7507_p1;
wire   [7:0] tmp_127_fu_7525_p4;
wire   [7:0] xor_ln1545_167_fu_7745_p2;
wire   [7:0] xor_ln1545_165_fu_7741_p2;
wire   [7:0] trunc_ln674_55_fu_7521_p1;
wire   [7:0] tmp_128_fu_7539_p4;
wire   [7:0] xor_ln1545_170_fu_7761_p2;
wire   [7:0] xor_ln1545_168_fu_7757_p2;
wire   [7:0] tmp_125_fu_7497_p4;
wire   [7:0] trunc_ln674_56_fu_7535_p1;
wire   [7:0] xor_ln1545_173_fu_7777_p2;
wire   [7:0] xor_ln1545_171_fu_7773_p2;
wire   [7:0] tmp_130_fu_7567_p4;
wire   [7:0] trunc_ln674_57_fu_7549_p1;
wire   [7:0] xor_ln1545_176_fu_7793_p2;
wire   [7:0] xor_ln1545_174_fu_7789_p2;
wire   [7:0] trunc_ln674_58_fu_7563_p1;
wire   [7:0] tmp_131_fu_7581_p4;
wire   [7:0] xor_ln1545_179_fu_7809_p2;
wire   [7:0] xor_ln1545_177_fu_7805_p2;
wire   [7:0] trunc_ln674_59_fu_7577_p1;
wire   [7:0] tmp_132_fu_7595_p4;
wire   [7:0] xor_ln1545_182_fu_7825_p2;
wire   [7:0] xor_ln1545_180_fu_7821_p2;
wire   [7:0] tmp_129_fu_7553_p4;
wire   [7:0] trunc_ln674_60_fu_7591_p1;
wire   [7:0] xor_ln1545_185_fu_7841_p2;
wire   [7:0] xor_ln1545_183_fu_7837_p2;
wire   [7:0] tmp_134_fu_7623_p4;
wire   [7:0] trunc_ln674_61_fu_7605_p1;
wire   [7:0] xor_ln1545_188_fu_7857_p2;
wire   [7:0] xor_ln1545_186_fu_7853_p2;
wire   [7:0] trunc_ln674_62_fu_7619_p1;
wire   [7:0] tmp_135_fu_7637_p4;
wire   [7:0] xor_ln1545_191_fu_7873_p2;
wire   [7:0] xor_ln1545_189_fu_7869_p2;
wire   [7:0] trunc_ln674_63_fu_7633_p1;
wire   [7:0] tmp_136_fu_7651_p4;
wire   [7:0] xor_ln1545_194_fu_7889_p2;
wire   [7:0] xor_ln1545_192_fu_7885_p2;
wire   [7:0] tmp_133_fu_7609_p4;
wire   [7:0] trunc_ln674_64_fu_7647_p1;
wire   [7:0] xor_ln1545_197_fu_7905_p2;
wire   [7:0] xor_ln1545_195_fu_7901_p2;
wire   [7:0] xor_ln1545_196_fu_7911_p2;
wire   [7:0] xor_ln1545_193_fu_7895_p2;
wire   [7:0] xor_ln1545_190_fu_7879_p2;
wire   [7:0] xor_ln1545_187_fu_7863_p2;
wire   [7:0] xor_ln1545_184_fu_7847_p2;
wire   [7:0] xor_ln1545_181_fu_7831_p2;
wire   [7:0] xor_ln1545_178_fu_7815_p2;
wire   [7:0] xor_ln1545_175_fu_7799_p2;
wire   [7:0] xor_ln1545_172_fu_7783_p2;
wire   [7:0] xor_ln1545_169_fu_7767_p2;
wire   [7:0] xor_ln1545_166_fu_7751_p2;
wire   [7:0] xor_ln1545_163_fu_7735_p2;
wire   [7:0] xor_ln1545_160_fu_7719_p2;
wire   [7:0] xor_ln1545_157_fu_7703_p2;
wire   [7:0] xor_ln1545_154_fu_7687_p2;
wire   [7:0] xor_ln1545_151_fu_7671_p2;
wire   [127:0] p_Result_27_fu_7917_p17;
wire   [127:0] state_V_27_fu_7953_p2;
wire   [7:0] trunc_ln708_4_fu_7958_p1;
wire   [7:0] tmp_137_fu_7967_p4;
wire   [7:0] tmp_138_fu_7982_p4;
wire   [7:0] tmp_139_fu_7997_p4;
wire   [7:0] tmp_140_fu_8012_p4;
wire   [7:0] tmp_141_fu_8027_p4;
wire   [7:0] tmp_142_fu_8042_p4;
wire   [7:0] tmp_143_fu_8057_p4;
wire   [7:0] tmp_144_fu_8072_p4;
wire   [7:0] tmp_145_fu_8087_p4;
wire   [7:0] tmp_146_fu_8102_p4;
wire   [7:0] tmp_147_fu_8117_p4;
wire   [7:0] tmp_148_fu_8132_p4;
wire   [7:0] tmp_149_fu_8147_p4;
wire   [7:0] tmp_150_fu_8162_p4;
wire   [7:0] tmp_151_fu_8177_p4;
wire   [7:0] tmp_153_fu_8290_p4;
wire   [7:0] trunc_ln674_65_fu_8272_p1;
wire   [7:0] xor_ln1545_200_fu_8500_p2;
wire   [7:0] xor_ln1545_198_fu_8496_p2;
wire   [7:0] trunc_ln674_66_fu_8286_p1;
wire   [7:0] tmp_154_fu_8304_p4;
wire   [7:0] xor_ln1545_203_fu_8516_p2;
wire   [7:0] xor_ln1545_201_fu_8512_p2;
wire   [7:0] trunc_ln674_67_fu_8300_p1;
wire   [7:0] tmp_155_fu_8318_p4;
wire   [7:0] xor_ln1545_206_fu_8532_p2;
wire   [7:0] xor_ln1545_204_fu_8528_p2;
wire   [7:0] tmp_152_fu_8276_p4;
wire   [7:0] trunc_ln674_68_fu_8314_p1;
wire   [7:0] xor_ln1545_209_fu_8548_p2;
wire   [7:0] xor_ln1545_207_fu_8544_p2;
wire   [7:0] tmp_157_fu_8346_p4;
wire   [7:0] trunc_ln674_69_fu_8328_p1;
wire   [7:0] xor_ln1545_212_fu_8564_p2;
wire   [7:0] xor_ln1545_210_fu_8560_p2;
wire   [7:0] trunc_ln674_70_fu_8342_p1;
wire   [7:0] tmp_158_fu_8360_p4;
wire   [7:0] xor_ln1545_215_fu_8580_p2;
wire   [7:0] xor_ln1545_213_fu_8576_p2;
wire   [7:0] trunc_ln674_71_fu_8356_p1;
wire   [7:0] tmp_159_fu_8374_p4;
wire   [7:0] xor_ln1545_218_fu_8596_p2;
wire   [7:0] xor_ln1545_216_fu_8592_p2;
wire   [7:0] tmp_156_fu_8332_p4;
wire   [7:0] trunc_ln674_72_fu_8370_p1;
wire   [7:0] xor_ln1545_221_fu_8612_p2;
wire   [7:0] xor_ln1545_219_fu_8608_p2;
wire   [7:0] tmp_161_fu_8402_p4;
wire   [7:0] trunc_ln674_73_fu_8384_p1;
wire   [7:0] xor_ln1545_224_fu_8628_p2;
wire   [7:0] xor_ln1545_222_fu_8624_p2;
wire   [7:0] trunc_ln674_74_fu_8398_p1;
wire   [7:0] tmp_162_fu_8416_p4;
wire   [7:0] xor_ln1545_227_fu_8644_p2;
wire   [7:0] xor_ln1545_225_fu_8640_p2;
wire   [7:0] trunc_ln674_75_fu_8412_p1;
wire   [7:0] tmp_163_fu_8430_p4;
wire   [7:0] xor_ln1545_230_fu_8660_p2;
wire   [7:0] xor_ln1545_228_fu_8656_p2;
wire   [7:0] tmp_160_fu_8388_p4;
wire   [7:0] trunc_ln674_76_fu_8426_p1;
wire   [7:0] xor_ln1545_233_fu_8676_p2;
wire   [7:0] xor_ln1545_231_fu_8672_p2;
wire   [7:0] tmp_165_fu_8458_p4;
wire   [7:0] trunc_ln674_77_fu_8440_p1;
wire   [7:0] xor_ln1545_236_fu_8692_p2;
wire   [7:0] xor_ln1545_234_fu_8688_p2;
wire   [7:0] trunc_ln674_78_fu_8454_p1;
wire   [7:0] tmp_166_fu_8472_p4;
wire   [7:0] xor_ln1545_239_fu_8708_p2;
wire   [7:0] xor_ln1545_237_fu_8704_p2;
wire   [7:0] trunc_ln674_79_fu_8468_p1;
wire   [7:0] tmp_167_fu_8486_p4;
wire   [7:0] xor_ln1545_242_fu_8724_p2;
wire   [7:0] xor_ln1545_240_fu_8720_p2;
wire   [7:0] tmp_164_fu_8444_p4;
wire   [7:0] trunc_ln674_80_fu_8482_p1;
wire   [7:0] xor_ln1545_245_fu_8740_p2;
wire   [7:0] xor_ln1545_243_fu_8736_p2;
wire   [7:0] xor_ln1545_244_fu_8746_p2;
wire   [7:0] xor_ln1545_241_fu_8730_p2;
wire   [7:0] xor_ln1545_238_fu_8714_p2;
wire   [7:0] xor_ln1545_235_fu_8698_p2;
wire   [7:0] xor_ln1545_232_fu_8682_p2;
wire   [7:0] xor_ln1545_229_fu_8666_p2;
wire   [7:0] xor_ln1545_226_fu_8650_p2;
wire   [7:0] xor_ln1545_223_fu_8634_p2;
wire   [7:0] xor_ln1545_220_fu_8618_p2;
wire   [7:0] xor_ln1545_217_fu_8602_p2;
wire   [7:0] xor_ln1545_214_fu_8586_p2;
wire   [7:0] xor_ln1545_211_fu_8570_p2;
wire   [7:0] xor_ln1545_208_fu_8554_p2;
wire   [7:0] xor_ln1545_205_fu_8538_p2;
wire   [7:0] xor_ln1545_202_fu_8522_p2;
wire   [7:0] xor_ln1545_199_fu_8506_p2;
wire   [127:0] p_Result_28_fu_8752_p17;
wire   [127:0] state_V_28_fu_8788_p2;
wire   [7:0] trunc_ln708_5_fu_8793_p1;
wire   [7:0] tmp_168_fu_8802_p4;
wire   [7:0] tmp_169_fu_8817_p4;
wire   [7:0] tmp_170_fu_8832_p4;
wire   [7:0] tmp_171_fu_8847_p4;
wire   [7:0] tmp_172_fu_8862_p4;
wire   [7:0] tmp_173_fu_8877_p4;
wire   [7:0] tmp_174_fu_8892_p4;
wire   [7:0] tmp_175_fu_8907_p4;
wire   [7:0] tmp_176_fu_8922_p4;
wire   [7:0] tmp_177_fu_8937_p4;
wire   [7:0] tmp_178_fu_8952_p4;
wire   [7:0] tmp_179_fu_8967_p4;
wire   [7:0] tmp_180_fu_8982_p4;
wire   [7:0] tmp_181_fu_8997_p4;
wire   [7:0] tmp_182_fu_9012_p4;
wire   [7:0] tmp_184_fu_9125_p4;
wire   [7:0] trunc_ln674_81_fu_9107_p1;
wire   [7:0] xor_ln1545_248_fu_9335_p2;
wire   [7:0] xor_ln1545_246_fu_9331_p2;
wire   [7:0] trunc_ln674_82_fu_9121_p1;
wire   [7:0] tmp_185_fu_9139_p4;
wire   [7:0] xor_ln1545_251_fu_9351_p2;
wire   [7:0] xor_ln1545_249_fu_9347_p2;
wire   [7:0] trunc_ln674_83_fu_9135_p1;
wire   [7:0] tmp_186_fu_9153_p4;
wire   [7:0] xor_ln1545_254_fu_9367_p2;
wire   [7:0] xor_ln1545_252_fu_9363_p2;
wire   [7:0] tmp_183_fu_9111_p4;
wire   [7:0] trunc_ln674_84_fu_9149_p1;
wire   [7:0] xor_ln1545_257_fu_9383_p2;
wire   [7:0] xor_ln1545_255_fu_9379_p2;
wire   [7:0] tmp_188_fu_9181_p4;
wire   [7:0] trunc_ln674_85_fu_9163_p1;
wire   [7:0] xor_ln1545_260_fu_9399_p2;
wire   [7:0] xor_ln1545_258_fu_9395_p2;
wire   [7:0] trunc_ln674_86_fu_9177_p1;
wire   [7:0] tmp_189_fu_9195_p4;
wire   [7:0] xor_ln1545_263_fu_9415_p2;
wire   [7:0] xor_ln1545_261_fu_9411_p2;
wire   [7:0] trunc_ln674_87_fu_9191_p1;
wire   [7:0] tmp_190_fu_9209_p4;
wire   [7:0] xor_ln1545_266_fu_9431_p2;
wire   [7:0] xor_ln1545_264_fu_9427_p2;
wire   [7:0] tmp_187_fu_9167_p4;
wire   [7:0] trunc_ln674_88_fu_9205_p1;
wire   [7:0] xor_ln1545_269_fu_9447_p2;
wire   [7:0] xor_ln1545_267_fu_9443_p2;
wire   [7:0] tmp_192_fu_9237_p4;
wire   [7:0] trunc_ln674_89_fu_9219_p1;
wire   [7:0] xor_ln1545_272_fu_9463_p2;
wire   [7:0] xor_ln1545_270_fu_9459_p2;
wire   [7:0] trunc_ln674_90_fu_9233_p1;
wire   [7:0] tmp_193_fu_9251_p4;
wire   [7:0] xor_ln1545_275_fu_9479_p2;
wire   [7:0] xor_ln1545_273_fu_9475_p2;
wire   [7:0] trunc_ln674_91_fu_9247_p1;
wire   [7:0] tmp_194_fu_9265_p4;
wire   [7:0] xor_ln1545_278_fu_9495_p2;
wire   [7:0] xor_ln1545_276_fu_9491_p2;
wire   [7:0] tmp_191_fu_9223_p4;
wire   [7:0] trunc_ln674_92_fu_9261_p1;
wire   [7:0] xor_ln1545_281_fu_9511_p2;
wire   [7:0] xor_ln1545_279_fu_9507_p2;
wire   [7:0] tmp_196_fu_9293_p4;
wire   [7:0] trunc_ln674_93_fu_9275_p1;
wire   [7:0] xor_ln1545_284_fu_9527_p2;
wire   [7:0] xor_ln1545_282_fu_9523_p2;
wire   [7:0] trunc_ln674_94_fu_9289_p1;
wire   [7:0] tmp_197_fu_9307_p4;
wire   [7:0] xor_ln1545_287_fu_9543_p2;
wire   [7:0] xor_ln1545_285_fu_9539_p2;
wire   [7:0] trunc_ln674_95_fu_9303_p1;
wire   [7:0] tmp_198_fu_9321_p4;
wire   [7:0] xor_ln1545_290_fu_9559_p2;
wire   [7:0] xor_ln1545_288_fu_9555_p2;
wire   [7:0] tmp_195_fu_9279_p4;
wire   [7:0] trunc_ln674_96_fu_9317_p1;
wire   [7:0] xor_ln1545_293_fu_9575_p2;
wire   [7:0] xor_ln1545_291_fu_9571_p2;
wire   [7:0] xor_ln1545_292_fu_9581_p2;
wire   [7:0] xor_ln1545_289_fu_9565_p2;
wire   [7:0] xor_ln1545_286_fu_9549_p2;
wire   [7:0] xor_ln1545_283_fu_9533_p2;
wire   [7:0] xor_ln1545_280_fu_9517_p2;
wire   [7:0] xor_ln1545_277_fu_9501_p2;
wire   [7:0] xor_ln1545_274_fu_9485_p2;
wire   [7:0] xor_ln1545_271_fu_9469_p2;
wire   [7:0] xor_ln1545_268_fu_9453_p2;
wire   [7:0] xor_ln1545_265_fu_9437_p2;
wire   [7:0] xor_ln1545_262_fu_9421_p2;
wire   [7:0] xor_ln1545_259_fu_9405_p2;
wire   [7:0] xor_ln1545_256_fu_9389_p2;
wire   [7:0] xor_ln1545_253_fu_9373_p2;
wire   [7:0] xor_ln1545_250_fu_9357_p2;
wire   [7:0] xor_ln1545_247_fu_9341_p2;
wire   [127:0] p_Result_29_fu_9587_p17;
wire   [127:0] state_V_29_fu_9623_p2;
wire   [7:0] trunc_ln708_6_fu_9628_p1;
wire   [7:0] tmp_199_fu_9637_p4;
wire   [7:0] tmp_200_fu_9652_p4;
wire   [7:0] tmp_201_fu_9667_p4;
wire   [7:0] tmp_202_fu_9682_p4;
wire   [7:0] tmp_203_fu_9697_p4;
wire   [7:0] tmp_204_fu_9712_p4;
wire   [7:0] tmp_205_fu_9727_p4;
wire   [7:0] tmp_206_fu_9742_p4;
wire   [7:0] tmp_207_fu_9757_p4;
wire   [7:0] tmp_208_fu_9772_p4;
wire   [7:0] tmp_209_fu_9787_p4;
wire   [7:0] tmp_210_fu_9802_p4;
wire   [7:0] tmp_211_fu_9817_p4;
wire   [7:0] tmp_212_fu_9832_p4;
wire   [7:0] tmp_213_fu_9847_p4;
wire   [7:0] tmp_215_fu_9960_p4;
wire   [7:0] trunc_ln674_97_fu_9942_p1;
wire   [7:0] xor_ln1545_296_fu_10170_p2;
wire   [7:0] xor_ln1545_294_fu_10166_p2;
wire   [7:0] trunc_ln674_98_fu_9956_p1;
wire   [7:0] tmp_216_fu_9974_p4;
wire   [7:0] xor_ln1545_299_fu_10186_p2;
wire   [7:0] xor_ln1545_297_fu_10182_p2;
wire   [7:0] trunc_ln674_99_fu_9970_p1;
wire   [7:0] tmp_217_fu_9988_p4;
wire   [7:0] xor_ln1545_302_fu_10202_p2;
wire   [7:0] xor_ln1545_300_fu_10198_p2;
wire   [7:0] tmp_214_fu_9946_p4;
wire   [7:0] trunc_ln674_100_fu_9984_p1;
wire   [7:0] xor_ln1545_305_fu_10218_p2;
wire   [7:0] xor_ln1545_303_fu_10214_p2;
wire   [7:0] tmp_219_fu_10016_p4;
wire   [7:0] trunc_ln674_101_fu_9998_p1;
wire   [7:0] xor_ln1545_308_fu_10234_p2;
wire   [7:0] xor_ln1545_306_fu_10230_p2;
wire   [7:0] trunc_ln674_102_fu_10012_p1;
wire   [7:0] tmp_220_fu_10030_p4;
wire   [7:0] xor_ln1545_311_fu_10250_p2;
wire   [7:0] xor_ln1545_309_fu_10246_p2;
wire   [7:0] trunc_ln674_103_fu_10026_p1;
wire   [7:0] tmp_221_fu_10044_p4;
wire   [7:0] xor_ln1545_314_fu_10266_p2;
wire   [7:0] xor_ln1545_312_fu_10262_p2;
wire   [7:0] tmp_218_fu_10002_p4;
wire   [7:0] trunc_ln674_104_fu_10040_p1;
wire   [7:0] xor_ln1545_317_fu_10282_p2;
wire   [7:0] xor_ln1545_315_fu_10278_p2;
wire   [7:0] tmp_223_fu_10072_p4;
wire   [7:0] trunc_ln674_105_fu_10054_p1;
wire   [7:0] xor_ln1545_320_fu_10298_p2;
wire   [7:0] xor_ln1545_318_fu_10294_p2;
wire   [7:0] trunc_ln674_106_fu_10068_p1;
wire   [7:0] tmp_224_fu_10086_p4;
wire   [7:0] xor_ln1545_323_fu_10314_p2;
wire   [7:0] xor_ln1545_321_fu_10310_p2;
wire   [7:0] trunc_ln674_107_fu_10082_p1;
wire   [7:0] tmp_225_fu_10100_p4;
wire   [7:0] xor_ln1545_326_fu_10330_p2;
wire   [7:0] xor_ln1545_324_fu_10326_p2;
wire   [7:0] tmp_222_fu_10058_p4;
wire   [7:0] trunc_ln674_108_fu_10096_p1;
wire   [7:0] xor_ln1545_329_fu_10346_p2;
wire   [7:0] xor_ln1545_327_fu_10342_p2;
wire   [7:0] tmp_227_fu_10128_p4;
wire   [7:0] trunc_ln674_109_fu_10110_p1;
wire   [7:0] xor_ln1545_332_fu_10362_p2;
wire   [7:0] xor_ln1545_330_fu_10358_p2;
wire   [7:0] trunc_ln674_110_fu_10124_p1;
wire   [7:0] tmp_228_fu_10142_p4;
wire   [7:0] xor_ln1545_335_fu_10378_p2;
wire   [7:0] xor_ln1545_333_fu_10374_p2;
wire   [7:0] trunc_ln674_111_fu_10138_p1;
wire   [7:0] tmp_229_fu_10156_p4;
wire   [7:0] xor_ln1545_338_fu_10394_p2;
wire   [7:0] xor_ln1545_336_fu_10390_p2;
wire   [7:0] tmp_226_fu_10114_p4;
wire   [7:0] trunc_ln674_112_fu_10152_p1;
wire   [7:0] xor_ln1545_341_fu_10410_p2;
wire   [7:0] xor_ln1545_339_fu_10406_p2;
wire   [7:0] xor_ln1545_340_fu_10416_p2;
wire   [7:0] xor_ln1545_337_fu_10400_p2;
wire   [7:0] xor_ln1545_334_fu_10384_p2;
wire   [7:0] xor_ln1545_331_fu_10368_p2;
wire   [7:0] xor_ln1545_328_fu_10352_p2;
wire   [7:0] xor_ln1545_325_fu_10336_p2;
wire   [7:0] xor_ln1545_322_fu_10320_p2;
wire   [7:0] xor_ln1545_319_fu_10304_p2;
wire   [7:0] xor_ln1545_316_fu_10288_p2;
wire   [7:0] xor_ln1545_313_fu_10272_p2;
wire   [7:0] xor_ln1545_310_fu_10256_p2;
wire   [7:0] xor_ln1545_307_fu_10240_p2;
wire   [7:0] xor_ln1545_304_fu_10224_p2;
wire   [7:0] xor_ln1545_301_fu_10208_p2;
wire   [7:0] xor_ln1545_298_fu_10192_p2;
wire   [7:0] xor_ln1545_295_fu_10176_p2;
wire   [127:0] p_Result_30_fu_10422_p17;
wire   [127:0] state_V_fu_10458_p2;
wire   [7:0] trunc_ln708_7_fu_10463_p1;
wire   [7:0] tmp_230_fu_10472_p4;
wire   [7:0] tmp_231_fu_10487_p4;
wire   [7:0] tmp_232_fu_10502_p4;
wire   [7:0] tmp_233_fu_10517_p4;
wire   [7:0] tmp_234_fu_10532_p4;
wire   [7:0] tmp_235_fu_10547_p4;
wire   [7:0] tmp_236_fu_10562_p4;
wire   [7:0] tmp_237_fu_10577_p4;
wire   [7:0] tmp_238_fu_10592_p4;
wire   [7:0] tmp_239_fu_10607_p4;
wire   [7:0] tmp_240_fu_10622_p4;
wire   [7:0] tmp_241_fu_10637_p4;
wire   [7:0] tmp_242_fu_10652_p4;
wire   [7:0] tmp_243_fu_10667_p4;
wire   [7:0] tmp_244_fu_10682_p4;
wire   [7:0] tmp_246_fu_10795_p4;
wire   [7:0] trunc_ln674_113_fu_10777_p1;
wire   [7:0] xor_ln1545_344_fu_11005_p2;
wire   [7:0] xor_ln1545_342_fu_11001_p2;
wire   [7:0] trunc_ln674_114_fu_10791_p1;
wire   [7:0] tmp_247_fu_10809_p4;
wire   [7:0] xor_ln1545_347_fu_11021_p2;
wire   [7:0] xor_ln1545_345_fu_11017_p2;
wire   [7:0] trunc_ln674_115_fu_10805_p1;
wire   [7:0] tmp_248_fu_10823_p4;
wire   [7:0] xor_ln1545_350_fu_11037_p2;
wire   [7:0] xor_ln1545_348_fu_11033_p2;
wire   [7:0] tmp_245_fu_10781_p4;
wire   [7:0] trunc_ln674_116_fu_10819_p1;
wire   [7:0] xor_ln1545_353_fu_11053_p2;
wire   [7:0] xor_ln1545_351_fu_11049_p2;
wire   [7:0] tmp_250_fu_10851_p4;
wire   [7:0] trunc_ln674_117_fu_10833_p1;
wire   [7:0] xor_ln1545_356_fu_11069_p2;
wire   [7:0] xor_ln1545_354_fu_11065_p2;
wire   [7:0] trunc_ln674_118_fu_10847_p1;
wire   [7:0] tmp_251_fu_10865_p4;
wire   [7:0] xor_ln1545_359_fu_11085_p2;
wire   [7:0] xor_ln1545_357_fu_11081_p2;
wire   [7:0] trunc_ln674_119_fu_10861_p1;
wire   [7:0] tmp_252_fu_10879_p4;
wire   [7:0] xor_ln1545_362_fu_11101_p2;
wire   [7:0] xor_ln1545_360_fu_11097_p2;
wire   [7:0] tmp_249_fu_10837_p4;
wire   [7:0] trunc_ln674_120_fu_10875_p1;
wire   [7:0] xor_ln1545_365_fu_11117_p2;
wire   [7:0] xor_ln1545_363_fu_11113_p2;
wire   [7:0] tmp_254_fu_10907_p4;
wire   [7:0] trunc_ln674_121_fu_10889_p1;
wire   [7:0] xor_ln1545_368_fu_11133_p2;
wire   [7:0] xor_ln1545_366_fu_11129_p2;
wire   [7:0] trunc_ln674_122_fu_10903_p1;
wire   [7:0] tmp_255_fu_10921_p4;
wire   [7:0] xor_ln1545_371_fu_11149_p2;
wire   [7:0] xor_ln1545_369_fu_11145_p2;
wire   [7:0] trunc_ln674_123_fu_10917_p1;
wire   [7:0] tmp_256_fu_10935_p4;
wire   [7:0] xor_ln1545_374_fu_11165_p2;
wire   [7:0] xor_ln1545_372_fu_11161_p2;
wire   [7:0] tmp_253_fu_10893_p4;
wire   [7:0] trunc_ln674_124_fu_10931_p1;
wire   [7:0] xor_ln1545_377_fu_11181_p2;
wire   [7:0] xor_ln1545_375_fu_11177_p2;
wire   [7:0] tmp_258_fu_10963_p4;
wire   [7:0] trunc_ln674_125_fu_10945_p1;
wire   [7:0] xor_ln1545_380_fu_11197_p2;
wire   [7:0] xor_ln1545_378_fu_11193_p2;
wire   [7:0] trunc_ln674_126_fu_10959_p1;
wire   [7:0] tmp_259_fu_10977_p4;
wire   [7:0] xor_ln1545_383_fu_11213_p2;
wire   [7:0] xor_ln1545_381_fu_11209_p2;
wire   [7:0] trunc_ln674_127_fu_10973_p1;
wire   [7:0] tmp_260_fu_10991_p4;
wire   [7:0] xor_ln1545_386_fu_11229_p2;
wire   [7:0] xor_ln1545_384_fu_11225_p2;
wire   [7:0] tmp_257_fu_10949_p4;
wire   [7:0] trunc_ln674_128_fu_10987_p1;
wire   [7:0] xor_ln1545_389_fu_11245_p2;
wire   [7:0] xor_ln1545_387_fu_11241_p2;
wire   [7:0] xor_ln1545_388_fu_11251_p2;
wire   [7:0] xor_ln1545_385_fu_11235_p2;
wire   [7:0] xor_ln1545_382_fu_11219_p2;
wire   [7:0] xor_ln1545_379_fu_11203_p2;
wire   [7:0] xor_ln1545_376_fu_11187_p2;
wire   [7:0] xor_ln1545_373_fu_11171_p2;
wire   [7:0] xor_ln1545_370_fu_11155_p2;
wire   [7:0] xor_ln1545_367_fu_11139_p2;
wire   [7:0] xor_ln1545_364_fu_11123_p2;
wire   [7:0] xor_ln1545_361_fu_11107_p2;
wire   [7:0] xor_ln1545_358_fu_11091_p2;
wire   [7:0] xor_ln1545_355_fu_11075_p2;
wire   [7:0] xor_ln1545_352_fu_11059_p2;
wire   [7:0] xor_ln1545_349_fu_11043_p2;
wire   [7:0] xor_ln1545_346_fu_11027_p2;
wire   [7:0] xor_ln1545_343_fu_11011_p2;
wire   [127:0] p_Result_31_fu_11257_p17;
wire   [127:0] state_V_30_fu_11293_p2;
wire   [7:0] trunc_ln708_8_fu_11298_p1;
wire   [7:0] tmp_261_fu_11307_p4;
wire   [7:0] tmp_262_fu_11322_p4;
wire   [7:0] tmp_263_fu_11337_p4;
wire   [7:0] tmp_264_fu_11352_p4;
wire   [7:0] tmp_265_fu_11367_p4;
wire   [7:0] tmp_266_fu_11382_p4;
wire   [7:0] tmp_267_fu_11397_p4;
wire   [7:0] tmp_268_fu_11412_p4;
wire   [7:0] tmp_269_fu_11427_p4;
wire   [7:0] tmp_270_fu_11442_p4;
wire   [7:0] tmp_271_fu_11457_p4;
wire   [7:0] tmp_272_fu_11472_p4;
wire   [7:0] tmp_273_fu_11487_p4;
wire   [7:0] tmp_274_fu_11502_p4;
wire   [7:0] tmp_275_fu_11517_p4;
wire   [7:0] tmp_277_fu_11630_p4;
wire   [7:0] trunc_ln674_129_fu_11612_p1;
wire   [7:0] xor_ln1545_392_fu_11840_p2;
wire   [7:0] xor_ln1545_390_fu_11836_p2;
wire   [7:0] trunc_ln674_130_fu_11626_p1;
wire   [7:0] tmp_278_fu_11644_p4;
wire   [7:0] xor_ln1545_395_fu_11856_p2;
wire   [7:0] xor_ln1545_393_fu_11852_p2;
wire   [7:0] trunc_ln674_131_fu_11640_p1;
wire   [7:0] tmp_279_fu_11658_p4;
wire   [7:0] xor_ln1545_398_fu_11872_p2;
wire   [7:0] xor_ln1545_396_fu_11868_p2;
wire   [7:0] tmp_276_fu_11616_p4;
wire   [7:0] trunc_ln674_132_fu_11654_p1;
wire   [7:0] xor_ln1545_401_fu_11888_p2;
wire   [7:0] xor_ln1545_399_fu_11884_p2;
wire   [7:0] tmp_281_fu_11686_p4;
wire   [7:0] trunc_ln674_133_fu_11668_p1;
wire   [7:0] xor_ln1545_404_fu_11904_p2;
wire   [7:0] xor_ln1545_402_fu_11900_p2;
wire   [7:0] trunc_ln674_134_fu_11682_p1;
wire   [7:0] tmp_282_fu_11700_p4;
wire   [7:0] xor_ln1545_407_fu_11920_p2;
wire   [7:0] xor_ln1545_405_fu_11916_p2;
wire   [7:0] trunc_ln674_135_fu_11696_p1;
wire   [7:0] tmp_283_fu_11714_p4;
wire   [7:0] xor_ln1545_410_fu_11936_p2;
wire   [7:0] xor_ln1545_408_fu_11932_p2;
wire   [7:0] tmp_280_fu_11672_p4;
wire   [7:0] trunc_ln674_136_fu_11710_p1;
wire   [7:0] xor_ln1545_413_fu_11952_p2;
wire   [7:0] xor_ln1545_411_fu_11948_p2;
wire   [7:0] tmp_285_fu_11742_p4;
wire   [7:0] trunc_ln674_137_fu_11724_p1;
wire   [7:0] xor_ln1545_416_fu_11968_p2;
wire   [7:0] xor_ln1545_414_fu_11964_p2;
wire   [7:0] trunc_ln674_138_fu_11738_p1;
wire   [7:0] tmp_286_fu_11756_p4;
wire   [7:0] xor_ln1545_419_fu_11984_p2;
wire   [7:0] xor_ln1545_417_fu_11980_p2;
wire   [7:0] trunc_ln674_139_fu_11752_p1;
wire   [7:0] tmp_287_fu_11770_p4;
wire   [7:0] xor_ln1545_422_fu_12000_p2;
wire   [7:0] xor_ln1545_420_fu_11996_p2;
wire   [7:0] tmp_284_fu_11728_p4;
wire   [7:0] trunc_ln674_140_fu_11766_p1;
wire   [7:0] xor_ln1545_425_fu_12016_p2;
wire   [7:0] xor_ln1545_423_fu_12012_p2;
wire   [7:0] tmp_289_fu_11798_p4;
wire   [7:0] trunc_ln674_141_fu_11780_p1;
wire   [7:0] xor_ln1545_428_fu_12032_p2;
wire   [7:0] xor_ln1545_426_fu_12028_p2;
wire   [7:0] trunc_ln674_142_fu_11794_p1;
wire   [7:0] tmp_290_fu_11812_p4;
wire   [7:0] xor_ln1545_431_fu_12048_p2;
wire   [7:0] xor_ln1545_429_fu_12044_p2;
wire   [7:0] trunc_ln674_143_fu_11808_p1;
wire   [7:0] tmp_291_fu_11826_p4;
wire   [7:0] xor_ln1545_434_fu_12064_p2;
wire   [7:0] xor_ln1545_432_fu_12060_p2;
wire   [7:0] tmp_288_fu_11784_p4;
wire   [7:0] trunc_ln674_144_fu_11822_p1;
wire   [7:0] xor_ln1545_437_fu_12080_p2;
wire   [7:0] xor_ln1545_435_fu_12076_p2;
wire   [7:0] xor_ln1545_436_fu_12086_p2;
wire   [7:0] xor_ln1545_433_fu_12070_p2;
wire   [7:0] xor_ln1545_430_fu_12054_p2;
wire   [7:0] xor_ln1545_427_fu_12038_p2;
wire   [7:0] xor_ln1545_424_fu_12022_p2;
wire   [7:0] xor_ln1545_421_fu_12006_p2;
wire   [7:0] xor_ln1545_418_fu_11990_p2;
wire   [7:0] xor_ln1545_415_fu_11974_p2;
wire   [7:0] xor_ln1545_412_fu_11958_p2;
wire   [7:0] xor_ln1545_409_fu_11942_p2;
wire   [7:0] xor_ln1545_406_fu_11926_p2;
wire   [7:0] xor_ln1545_403_fu_11910_p2;
wire   [7:0] xor_ln1545_400_fu_11894_p2;
wire   [7:0] xor_ln1545_397_fu_11878_p2;
wire   [7:0] xor_ln1545_394_fu_11862_p2;
wire   [7:0] xor_ln1545_391_fu_11846_p2;
wire   [127:0] p_Result_32_fu_12092_p17;
wire   [127:0] state_V_31_fu_12128_p2;
wire   [7:0] trunc_ln708_9_fu_12133_p1;
wire   [7:0] tmp_292_fu_12142_p4;
wire   [7:0] tmp_293_fu_12157_p4;
wire   [7:0] tmp_294_fu_12172_p4;
wire   [7:0] tmp_295_fu_12187_p4;
wire   [7:0] tmp_296_fu_12202_p4;
wire   [7:0] tmp_297_fu_12217_p4;
wire   [7:0] tmp_298_fu_12232_p4;
wire   [7:0] tmp_299_fu_12247_p4;
wire   [7:0] tmp_300_fu_12262_p4;
wire   [7:0] tmp_301_fu_12277_p4;
wire   [7:0] tmp_302_fu_12292_p4;
wire   [7:0] tmp_303_fu_12307_p4;
wire   [7:0] tmp_304_fu_12322_p4;
wire   [7:0] tmp_305_fu_12337_p4;
wire   [7:0] tmp_306_fu_12352_p4;
wire   [7:0] tmp_308_fu_12465_p4;
wire   [7:0] trunc_ln674_145_fu_12447_p1;
wire   [7:0] xor_ln1545_440_fu_12675_p2;
wire   [7:0] xor_ln1545_438_fu_12671_p2;
wire   [7:0] trunc_ln674_146_fu_12461_p1;
wire   [7:0] tmp_309_fu_12479_p4;
wire   [7:0] xor_ln1545_443_fu_12691_p2;
wire   [7:0] xor_ln1545_441_fu_12687_p2;
wire   [7:0] trunc_ln674_147_fu_12475_p1;
wire   [7:0] tmp_310_fu_12493_p4;
wire   [7:0] xor_ln1545_446_fu_12707_p2;
wire   [7:0] xor_ln1545_444_fu_12703_p2;
wire   [7:0] tmp_307_fu_12451_p4;
wire   [7:0] trunc_ln674_148_fu_12489_p1;
wire   [7:0] xor_ln1545_449_fu_12723_p2;
wire   [7:0] xor_ln1545_447_fu_12719_p2;
wire   [7:0] tmp_312_fu_12521_p4;
wire   [7:0] trunc_ln674_149_fu_12503_p1;
wire   [7:0] xor_ln1545_452_fu_12739_p2;
wire   [7:0] xor_ln1545_450_fu_12735_p2;
wire   [7:0] trunc_ln674_150_fu_12517_p1;
wire   [7:0] tmp_313_fu_12535_p4;
wire   [7:0] xor_ln1545_455_fu_12755_p2;
wire   [7:0] xor_ln1545_453_fu_12751_p2;
wire   [7:0] trunc_ln674_151_fu_12531_p1;
wire   [7:0] tmp_314_fu_12549_p4;
wire   [7:0] xor_ln1545_458_fu_12771_p2;
wire   [7:0] xor_ln1545_456_fu_12767_p2;
wire   [7:0] tmp_311_fu_12507_p4;
wire   [7:0] trunc_ln674_152_fu_12545_p1;
wire   [7:0] xor_ln1545_461_fu_12787_p2;
wire   [7:0] xor_ln1545_459_fu_12783_p2;
wire   [7:0] tmp_316_fu_12577_p4;
wire   [7:0] trunc_ln674_153_fu_12559_p1;
wire   [7:0] xor_ln1545_464_fu_12803_p2;
wire   [7:0] xor_ln1545_462_fu_12799_p2;
wire   [7:0] trunc_ln674_154_fu_12573_p1;
wire   [7:0] tmp_317_fu_12591_p4;
wire   [7:0] xor_ln1545_467_fu_12819_p2;
wire   [7:0] xor_ln1545_465_fu_12815_p2;
wire   [7:0] trunc_ln674_155_fu_12587_p1;
wire   [7:0] tmp_318_fu_12605_p4;
wire   [7:0] xor_ln1545_470_fu_12835_p2;
wire   [7:0] xor_ln1545_468_fu_12831_p2;
wire   [7:0] tmp_315_fu_12563_p4;
wire   [7:0] trunc_ln674_156_fu_12601_p1;
wire   [7:0] xor_ln1545_473_fu_12851_p2;
wire   [7:0] xor_ln1545_471_fu_12847_p2;
wire   [7:0] tmp_320_fu_12633_p4;
wire   [7:0] trunc_ln674_157_fu_12615_p1;
wire   [7:0] xor_ln1545_476_fu_12867_p2;
wire   [7:0] xor_ln1545_474_fu_12863_p2;
wire   [7:0] trunc_ln674_158_fu_12629_p1;
wire   [7:0] tmp_321_fu_12647_p4;
wire   [7:0] xor_ln1545_479_fu_12883_p2;
wire   [7:0] xor_ln1545_477_fu_12879_p2;
wire   [7:0] trunc_ln674_159_fu_12643_p1;
wire   [7:0] tmp_322_fu_12661_p4;
wire   [7:0] xor_ln1545_482_fu_12899_p2;
wire   [7:0] xor_ln1545_480_fu_12895_p2;
wire   [7:0] tmp_319_fu_12619_p4;
wire   [7:0] trunc_ln674_160_fu_12657_p1;
wire   [7:0] xor_ln1545_485_fu_12915_p2;
wire   [7:0] xor_ln1545_483_fu_12911_p2;
wire   [7:0] xor_ln1545_484_fu_12921_p2;
wire   [7:0] xor_ln1545_481_fu_12905_p2;
wire   [7:0] xor_ln1545_478_fu_12889_p2;
wire   [7:0] xor_ln1545_475_fu_12873_p2;
wire   [7:0] xor_ln1545_472_fu_12857_p2;
wire   [7:0] xor_ln1545_469_fu_12841_p2;
wire   [7:0] xor_ln1545_466_fu_12825_p2;
wire   [7:0] xor_ln1545_463_fu_12809_p2;
wire   [7:0] xor_ln1545_460_fu_12793_p2;
wire   [7:0] xor_ln1545_457_fu_12777_p2;
wire   [7:0] xor_ln1545_454_fu_12761_p2;
wire   [7:0] xor_ln1545_451_fu_12745_p2;
wire   [7:0] xor_ln1545_448_fu_12729_p2;
wire   [7:0] xor_ln1545_445_fu_12713_p2;
wire   [7:0] xor_ln1545_442_fu_12697_p2;
wire   [7:0] xor_ln1545_439_fu_12681_p2;
wire   [127:0] p_Result_33_fu_12927_p17;
wire   [127:0] state_V_32_fu_12963_p2;
wire   [7:0] trunc_ln708_10_fu_12968_p1;
wire   [7:0] tmp_323_fu_12977_p4;
wire   [7:0] tmp_324_fu_12992_p4;
wire   [7:0] tmp_325_fu_13007_p4;
wire   [7:0] tmp_326_fu_13022_p4;
wire   [7:0] tmp_327_fu_13037_p4;
wire   [7:0] tmp_328_fu_13052_p4;
wire   [7:0] tmp_329_fu_13067_p4;
wire   [7:0] tmp_330_fu_13082_p4;
wire   [7:0] tmp_331_fu_13097_p4;
wire   [7:0] tmp_332_fu_13112_p4;
wire   [7:0] tmp_333_fu_13127_p4;
wire   [7:0] tmp_334_fu_13142_p4;
wire   [7:0] tmp_335_fu_13157_p4;
wire   [7:0] tmp_336_fu_13172_p4;
wire   [7:0] tmp_337_fu_13187_p4;
wire   [7:0] tmp_339_fu_13300_p4;
wire   [7:0] trunc_ln674_161_fu_13282_p1;
wire   [7:0] xor_ln1545_488_fu_13510_p2;
wire   [7:0] xor_ln1545_486_fu_13506_p2;
wire   [7:0] trunc_ln674_162_fu_13296_p1;
wire   [7:0] tmp_340_fu_13314_p4;
wire   [7:0] xor_ln1545_491_fu_13526_p2;
wire   [7:0] xor_ln1545_489_fu_13522_p2;
wire   [7:0] trunc_ln674_163_fu_13310_p1;
wire   [7:0] tmp_341_fu_13328_p4;
wire   [7:0] xor_ln1545_494_fu_13542_p2;
wire   [7:0] xor_ln1545_492_fu_13538_p2;
wire   [7:0] tmp_338_fu_13286_p4;
wire   [7:0] trunc_ln674_164_fu_13324_p1;
wire   [7:0] xor_ln1545_497_fu_13558_p2;
wire   [7:0] xor_ln1545_495_fu_13554_p2;
wire   [7:0] tmp_343_fu_13356_p4;
wire   [7:0] trunc_ln674_165_fu_13338_p1;
wire   [7:0] xor_ln1545_500_fu_13574_p2;
wire   [7:0] xor_ln1545_498_fu_13570_p2;
wire   [7:0] trunc_ln674_166_fu_13352_p1;
wire   [7:0] tmp_344_fu_13370_p4;
wire   [7:0] xor_ln1545_503_fu_13590_p2;
wire   [7:0] xor_ln1545_501_fu_13586_p2;
wire   [7:0] trunc_ln674_167_fu_13366_p1;
wire   [7:0] tmp_345_fu_13384_p4;
wire   [7:0] xor_ln1545_506_fu_13606_p2;
wire   [7:0] xor_ln1545_504_fu_13602_p2;
wire   [7:0] tmp_342_fu_13342_p4;
wire   [7:0] trunc_ln674_168_fu_13380_p1;
wire   [7:0] xor_ln1545_509_fu_13622_p2;
wire   [7:0] xor_ln1545_507_fu_13618_p2;
wire   [7:0] tmp_347_fu_13412_p4;
wire   [7:0] trunc_ln674_169_fu_13394_p1;
wire   [7:0] xor_ln1545_512_fu_13638_p2;
wire   [7:0] xor_ln1545_510_fu_13634_p2;
wire   [7:0] trunc_ln674_170_fu_13408_p1;
wire   [7:0] tmp_348_fu_13426_p4;
wire   [7:0] xor_ln1545_515_fu_13654_p2;
wire   [7:0] xor_ln1545_513_fu_13650_p2;
wire   [7:0] trunc_ln674_171_fu_13422_p1;
wire   [7:0] tmp_349_fu_13440_p4;
wire   [7:0] xor_ln1545_518_fu_13670_p2;
wire   [7:0] xor_ln1545_516_fu_13666_p2;
wire   [7:0] tmp_346_fu_13398_p4;
wire   [7:0] trunc_ln674_172_fu_13436_p1;
wire   [7:0] xor_ln1545_521_fu_13686_p2;
wire   [7:0] xor_ln1545_519_fu_13682_p2;
wire   [7:0] tmp_351_fu_13468_p4;
wire   [7:0] trunc_ln674_173_fu_13450_p1;
wire   [7:0] xor_ln1545_524_fu_13702_p2;
wire   [7:0] xor_ln1545_522_fu_13698_p2;
wire   [7:0] trunc_ln674_174_fu_13464_p1;
wire   [7:0] tmp_352_fu_13482_p4;
wire   [7:0] xor_ln1545_527_fu_13718_p2;
wire   [7:0] xor_ln1545_525_fu_13714_p2;
wire   [7:0] trunc_ln674_175_fu_13478_p1;
wire   [7:0] tmp_353_fu_13496_p4;
wire   [7:0] xor_ln1545_530_fu_13734_p2;
wire   [7:0] xor_ln1545_528_fu_13730_p2;
wire   [7:0] tmp_350_fu_13454_p4;
wire   [7:0] trunc_ln674_176_fu_13492_p1;
wire   [7:0] xor_ln1545_533_fu_13750_p2;
wire   [7:0] xor_ln1545_531_fu_13746_p2;
wire   [7:0] xor_ln1545_532_fu_13756_p2;
wire   [7:0] xor_ln1545_529_fu_13740_p2;
wire   [7:0] xor_ln1545_526_fu_13724_p2;
wire   [7:0] xor_ln1545_523_fu_13708_p2;
wire   [7:0] xor_ln1545_520_fu_13692_p2;
wire   [7:0] xor_ln1545_517_fu_13676_p2;
wire   [7:0] xor_ln1545_514_fu_13660_p2;
wire   [7:0] xor_ln1545_511_fu_13644_p2;
wire   [7:0] xor_ln1545_508_fu_13628_p2;
wire   [7:0] xor_ln1545_505_fu_13612_p2;
wire   [7:0] xor_ln1545_502_fu_13596_p2;
wire   [7:0] xor_ln1545_499_fu_13580_p2;
wire   [7:0] xor_ln1545_496_fu_13564_p2;
wire   [7:0] xor_ln1545_493_fu_13548_p2;
wire   [7:0] xor_ln1545_490_fu_13532_p2;
wire   [7:0] xor_ln1545_487_fu_13516_p2;
wire   [127:0] p_Result_34_fu_13762_p17;
wire   [127:0] state_V_33_fu_13798_p2;
wire   [7:0] trunc_ln708_11_fu_13803_p1;
wire   [7:0] tmp_354_fu_13812_p4;
wire   [7:0] tmp_355_fu_13827_p4;
wire   [7:0] tmp_356_fu_13842_p4;
wire   [7:0] tmp_357_fu_13857_p4;
wire   [7:0] tmp_358_fu_13872_p4;
wire   [7:0] tmp_359_fu_13887_p4;
wire   [7:0] tmp_360_fu_13902_p4;
wire   [7:0] tmp_361_fu_13917_p4;
wire   [7:0] tmp_362_fu_13932_p4;
wire   [7:0] tmp_363_fu_13947_p4;
wire   [7:0] tmp_364_fu_13962_p4;
wire   [7:0] tmp_365_fu_13977_p4;
wire   [7:0] tmp_366_fu_13992_p4;
wire   [7:0] tmp_367_fu_14007_p4;
wire   [7:0] tmp_368_fu_14022_p4;
wire   [127:0] p_Result_35_fu_14037_p17;
reg   [0:0] ap_NS_fsm;
reg    ap_idle_pp0_0to22;
reg    ap_reset_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 1'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter5 = 1'b0;
#0 ap_enable_reg_pp0_iter6 = 1'b0;
#0 ap_enable_reg_pp0_iter7 = 1'b0;
#0 ap_enable_reg_pp0_iter8 = 1'b0;
#0 ap_enable_reg_pp0_iter9 = 1'b0;
#0 ap_enable_reg_pp0_iter10 = 1'b0;
#0 ap_enable_reg_pp0_iter11 = 1'b0;
#0 ap_enable_reg_pp0_iter12 = 1'b0;
#0 ap_enable_reg_pp0_iter13 = 1'b0;
#0 ap_enable_reg_pp0_iter14 = 1'b0;
#0 ap_enable_reg_pp0_iter15 = 1'b0;
#0 ap_enable_reg_pp0_iter16 = 1'b0;
#0 ap_enable_reg_pp0_iter17 = 1'b0;
#0 ap_enable_reg_pp0_iter18 = 1'b0;
#0 ap_enable_reg_pp0_iter19 = 1'b0;
#0 ap_enable_reg_pp0_iter20 = 1'b0;
#0 ap_enable_reg_pp0_iter21 = 1'b0;
#0 ap_enable_reg_pp0_iter22 = 1'b0;
#0 ap_enable_reg_pp0_iter23 = 1'b0;
end

testEnc_process_r_cipher_0_ssbox_ROM_NP_LUTRAM_1R #(
    .DataWidth( 8 ),
    .AddressRange( 256 ),
    .AddressWidth( 8 ))
cipher_0_ssbox_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(cipher_0_ssbox_address0),
    .ce0(cipher_0_ssbox_ce0),
    .q0(cipher_0_ssbox_q0),
    .address1(cipher_0_ssbox_address1),
    .ce1(cipher_0_ssbox_ce1),
    .q1(cipher_0_ssbox_q1),
    .address2(cipher_0_ssbox_address2),
    .ce2(cipher_0_ssbox_ce2),
    .q2(cipher_0_ssbox_q2),
    .address3(cipher_0_ssbox_address3),
    .ce3(cipher_0_ssbox_ce3),
    .q3(cipher_0_ssbox_q3),
    .address4(cipher_0_ssbox_address4),
    .ce4(cipher_0_ssbox_ce4),
    .q4(cipher_0_ssbox_q4),
    .address5(cipher_0_ssbox_address5),
    .ce5(cipher_0_ssbox_ce5),
    .q5(cipher_0_ssbox_q5),
    .address6(cipher_0_ssbox_address6),
    .ce6(cipher_0_ssbox_ce6),
    .q6(cipher_0_ssbox_q6),
    .address7(cipher_0_ssbox_address7),
    .ce7(cipher_0_ssbox_ce7),
    .q7(cipher_0_ssbox_q7),
    .address8(cipher_0_ssbox_address8),
    .ce8(cipher_0_ssbox_ce8),
    .q8(cipher_0_ssbox_q8),
    .address9(cipher_0_ssbox_address9),
    .ce9(cipher_0_ssbox_ce9),
    .q9(cipher_0_ssbox_q9),
    .address10(cipher_0_ssbox_address10),
    .ce10(cipher_0_ssbox_ce10),
    .q10(cipher_0_ssbox_q10),
    .address11(cipher_0_ssbox_address11),
    .ce11(cipher_0_ssbox_ce11),
    .q11(cipher_0_ssbox_q11),
    .address12(cipher_0_ssbox_address12),
    .ce12(cipher_0_ssbox_ce12),
    .q12(cipher_0_ssbox_q12),
    .address13(cipher_0_ssbox_address13),
    .ce13(cipher_0_ssbox_ce13),
    .q13(cipher_0_ssbox_q13),
    .address14(cipher_0_ssbox_address14),
    .ce14(cipher_0_ssbox_ce14),
    .q14(cipher_0_ssbox_q14),
    .address15(cipher_0_ssbox_address15),
    .ce15(cipher_0_ssbox_ce15),
    .q15(cipher_0_ssbox_q15),
    .address16(cipher_0_ssbox_address16),
    .ce16(cipher_0_ssbox_ce16),
    .q16(cipher_0_ssbox_q16),
    .address17(cipher_0_ssbox_address17),
    .ce17(cipher_0_ssbox_ce17),
    .q17(cipher_0_ssbox_q17),
    .address18(cipher_0_ssbox_address18),
    .ce18(cipher_0_ssbox_ce18),
    .q18(cipher_0_ssbox_q18),
    .address19(cipher_0_ssbox_address19),
    .ce19(cipher_0_ssbox_ce19),
    .q19(cipher_0_ssbox_q19),
    .address20(cipher_0_ssbox_address20),
    .ce20(cipher_0_ssbox_ce20),
    .q20(cipher_0_ssbox_q20),
    .address21(cipher_0_ssbox_address21),
    .ce21(cipher_0_ssbox_ce21),
    .q21(cipher_0_ssbox_q21),
    .address22(cipher_0_ssbox_address22),
    .ce22(cipher_0_ssbox_ce22),
    .q22(cipher_0_ssbox_q22),
    .address23(cipher_0_ssbox_address23),
    .ce23(cipher_0_ssbox_ce23),
    .q23(cipher_0_ssbox_q23),
    .address24(cipher_0_ssbox_address24),
    .ce24(cipher_0_ssbox_ce24),
    .q24(cipher_0_ssbox_q24),
    .address25(cipher_0_ssbox_address25),
    .ce25(cipher_0_ssbox_ce25),
    .q25(cipher_0_ssbox_q25),
    .address26(cipher_0_ssbox_address26),
    .ce26(cipher_0_ssbox_ce26),
    .q26(cipher_0_ssbox_q26),
    .address27(cipher_0_ssbox_address27),
    .ce27(cipher_0_ssbox_ce27),
    .q27(cipher_0_ssbox_q27),
    .address28(cipher_0_ssbox_address28),
    .ce28(cipher_0_ssbox_ce28),
    .q28(cipher_0_ssbox_q28),
    .address29(cipher_0_ssbox_address29),
    .ce29(cipher_0_ssbox_ce29),
    .q29(cipher_0_ssbox_q29),
    .address30(cipher_0_ssbox_address30),
    .ce30(cipher_0_ssbox_ce30),
    .q30(cipher_0_ssbox_q30),
    .address31(cipher_0_ssbox_address31),
    .ce31(cipher_0_ssbox_ce31),
    .q31(cipher_0_ssbox_q31),
    .address32(cipher_0_ssbox_address32),
    .ce32(cipher_0_ssbox_ce32),
    .q32(cipher_0_ssbox_q32),
    .address33(cipher_0_ssbox_address33),
    .ce33(cipher_0_ssbox_ce33),
    .q33(cipher_0_ssbox_q33),
    .address34(cipher_0_ssbox_address34),
    .ce34(cipher_0_ssbox_ce34),
    .q34(cipher_0_ssbox_q34),
    .address35(cipher_0_ssbox_address35),
    .ce35(cipher_0_ssbox_ce35),
    .q35(cipher_0_ssbox_q35),
    .address36(cipher_0_ssbox_address36),
    .ce36(cipher_0_ssbox_ce36),
    .q36(cipher_0_ssbox_q36),
    .address37(cipher_0_ssbox_address37),
    .ce37(cipher_0_ssbox_ce37),
    .q37(cipher_0_ssbox_q37),
    .address38(cipher_0_ssbox_address38),
    .ce38(cipher_0_ssbox_ce38),
    .q38(cipher_0_ssbox_q38),
    .address39(cipher_0_ssbox_address39),
    .ce39(cipher_0_ssbox_ce39),
    .q39(cipher_0_ssbox_q39),
    .address40(cipher_0_ssbox_address40),
    .ce40(cipher_0_ssbox_ce40),
    .q40(cipher_0_ssbox_q40),
    .address41(cipher_0_ssbox_address41),
    .ce41(cipher_0_ssbox_ce41),
    .q41(cipher_0_ssbox_q41),
    .address42(cipher_0_ssbox_address42),
    .ce42(cipher_0_ssbox_ce42),
    .q42(cipher_0_ssbox_q42),
    .address43(cipher_0_ssbox_address43),
    .ce43(cipher_0_ssbox_ce43),
    .q43(cipher_0_ssbox_q43),
    .address44(cipher_0_ssbox_address44),
    .ce44(cipher_0_ssbox_ce44),
    .q44(cipher_0_ssbox_q44),
    .address45(cipher_0_ssbox_address45),
    .ce45(cipher_0_ssbox_ce45),
    .q45(cipher_0_ssbox_q45),
    .address46(cipher_0_ssbox_address46),
    .ce46(cipher_0_ssbox_ce46),
    .q46(cipher_0_ssbox_q46),
    .address47(cipher_0_ssbox_address47),
    .ce47(cipher_0_ssbox_ce47),
    .q47(cipher_0_ssbox_q47),
    .address48(cipher_0_ssbox_address48),
    .ce48(cipher_0_ssbox_ce48),
    .q48(cipher_0_ssbox_q48),
    .address49(cipher_0_ssbox_address49),
    .ce49(cipher_0_ssbox_ce49),
    .q49(cipher_0_ssbox_q49),
    .address50(cipher_0_ssbox_address50),
    .ce50(cipher_0_ssbox_ce50),
    .q50(cipher_0_ssbox_q50),
    .address51(cipher_0_ssbox_address51),
    .ce51(cipher_0_ssbox_ce51),
    .q51(cipher_0_ssbox_q51),
    .address52(cipher_0_ssbox_address52),
    .ce52(cipher_0_ssbox_ce52),
    .q52(cipher_0_ssbox_q52),
    .address53(cipher_0_ssbox_address53),
    .ce53(cipher_0_ssbox_ce53),
    .q53(cipher_0_ssbox_q53),
    .address54(cipher_0_ssbox_address54),
    .ce54(cipher_0_ssbox_ce54),
    .q54(cipher_0_ssbox_q54),
    .address55(cipher_0_ssbox_address55),
    .ce55(cipher_0_ssbox_ce55),
    .q55(cipher_0_ssbox_q55),
    .address56(cipher_0_ssbox_address56),
    .ce56(cipher_0_ssbox_ce56),
    .q56(cipher_0_ssbox_q56),
    .address57(cipher_0_ssbox_address57),
    .ce57(cipher_0_ssbox_ce57),
    .q57(cipher_0_ssbox_q57),
    .address58(cipher_0_ssbox_address58),
    .ce58(cipher_0_ssbox_ce58),
    .q58(cipher_0_ssbox_q58),
    .address59(cipher_0_ssbox_address59),
    .ce59(cipher_0_ssbox_ce59),
    .q59(cipher_0_ssbox_q59),
    .address60(cipher_0_ssbox_address60),
    .ce60(cipher_0_ssbox_ce60),
    .q60(cipher_0_ssbox_q60),
    .address61(cipher_0_ssbox_address61),
    .ce61(cipher_0_ssbox_ce61),
    .q61(cipher_0_ssbox_q61),
    .address62(cipher_0_ssbox_address62),
    .ce62(cipher_0_ssbox_ce62),
    .q62(cipher_0_ssbox_q62),
    .address63(cipher_0_ssbox_address63),
    .ce63(cipher_0_ssbox_ce63),
    .q63(cipher_0_ssbox_q63),
    .address64(cipher_0_ssbox_address64),
    .ce64(cipher_0_ssbox_ce64),
    .q64(cipher_0_ssbox_q64),
    .address65(cipher_0_ssbox_address65),
    .ce65(cipher_0_ssbox_ce65),
    .q65(cipher_0_ssbox_q65),
    .address66(cipher_0_ssbox_address66),
    .ce66(cipher_0_ssbox_ce66),
    .q66(cipher_0_ssbox_q66),
    .address67(cipher_0_ssbox_address67),
    .ce67(cipher_0_ssbox_ce67),
    .q67(cipher_0_ssbox_q67),
    .address68(cipher_0_ssbox_address68),
    .ce68(cipher_0_ssbox_ce68),
    .q68(cipher_0_ssbox_q68),
    .address69(cipher_0_ssbox_address69),
    .ce69(cipher_0_ssbox_ce69),
    .q69(cipher_0_ssbox_q69),
    .address70(cipher_0_ssbox_address70),
    .ce70(cipher_0_ssbox_ce70),
    .q70(cipher_0_ssbox_q70),
    .address71(cipher_0_ssbox_address71),
    .ce71(cipher_0_ssbox_ce71),
    .q71(cipher_0_ssbox_q71),
    .address72(cipher_0_ssbox_address72),
    .ce72(cipher_0_ssbox_ce72),
    .q72(cipher_0_ssbox_q72),
    .address73(cipher_0_ssbox_address73),
    .ce73(cipher_0_ssbox_ce73),
    .q73(cipher_0_ssbox_q73),
    .address74(cipher_0_ssbox_address74),
    .ce74(cipher_0_ssbox_ce74),
    .q74(cipher_0_ssbox_q74),
    .address75(cipher_0_ssbox_address75),
    .ce75(cipher_0_ssbox_ce75),
    .q75(cipher_0_ssbox_q75),
    .address76(cipher_0_ssbox_address76),
    .ce76(cipher_0_ssbox_ce76),
    .q76(cipher_0_ssbox_q76),
    .address77(cipher_0_ssbox_address77),
    .ce77(cipher_0_ssbox_ce77),
    .q77(cipher_0_ssbox_q77),
    .address78(cipher_0_ssbox_address78),
    .ce78(cipher_0_ssbox_ce78),
    .q78(cipher_0_ssbox_q78),
    .address79(cipher_0_ssbox_address79),
    .ce79(cipher_0_ssbox_ce79),
    .q79(cipher_0_ssbox_q79),
    .address80(cipher_0_ssbox_address80),
    .ce80(cipher_0_ssbox_ce80),
    .q80(cipher_0_ssbox_q80),
    .address81(cipher_0_ssbox_address81),
    .ce81(cipher_0_ssbox_ce81),
    .q81(cipher_0_ssbox_q81),
    .address82(cipher_0_ssbox_address82),
    .ce82(cipher_0_ssbox_ce82),
    .q82(cipher_0_ssbox_q82),
    .address83(cipher_0_ssbox_address83),
    .ce83(cipher_0_ssbox_ce83),
    .q83(cipher_0_ssbox_q83),
    .address84(cipher_0_ssbox_address84),
    .ce84(cipher_0_ssbox_ce84),
    .q84(cipher_0_ssbox_q84),
    .address85(cipher_0_ssbox_address85),
    .ce85(cipher_0_ssbox_ce85),
    .q85(cipher_0_ssbox_q85),
    .address86(cipher_0_ssbox_address86),
    .ce86(cipher_0_ssbox_ce86),
    .q86(cipher_0_ssbox_q86),
    .address87(cipher_0_ssbox_address87),
    .ce87(cipher_0_ssbox_ce87),
    .q87(cipher_0_ssbox_q87),
    .address88(cipher_0_ssbox_address88),
    .ce88(cipher_0_ssbox_ce88),
    .q88(cipher_0_ssbox_q88),
    .address89(cipher_0_ssbox_address89),
    .ce89(cipher_0_ssbox_ce89),
    .q89(cipher_0_ssbox_q89),
    .address90(cipher_0_ssbox_address90),
    .ce90(cipher_0_ssbox_ce90),
    .q90(cipher_0_ssbox_q90),
    .address91(cipher_0_ssbox_address91),
    .ce91(cipher_0_ssbox_ce91),
    .q91(cipher_0_ssbox_q91),
    .address92(cipher_0_ssbox_address92),
    .ce92(cipher_0_ssbox_ce92),
    .q92(cipher_0_ssbox_q92),
    .address93(cipher_0_ssbox_address93),
    .ce93(cipher_0_ssbox_ce93),
    .q93(cipher_0_ssbox_q93),
    .address94(cipher_0_ssbox_address94),
    .ce94(cipher_0_ssbox_ce94),
    .q94(cipher_0_ssbox_q94),
    .address95(cipher_0_ssbox_address95),
    .ce95(cipher_0_ssbox_ce95),
    .q95(cipher_0_ssbox_q95),
    .address96(cipher_0_ssbox_address96),
    .ce96(cipher_0_ssbox_ce96),
    .q96(cipher_0_ssbox_q96),
    .address97(cipher_0_ssbox_address97),
    .ce97(cipher_0_ssbox_ce97),
    .q97(cipher_0_ssbox_q97),
    .address98(cipher_0_ssbox_address98),
    .ce98(cipher_0_ssbox_ce98),
    .q98(cipher_0_ssbox_q98),
    .address99(cipher_0_ssbox_address99),
    .ce99(cipher_0_ssbox_ce99),
    .q99(cipher_0_ssbox_q99),
    .address100(cipher_0_ssbox_address100),
    .ce100(cipher_0_ssbox_ce100),
    .q100(cipher_0_ssbox_q100),
    .address101(cipher_0_ssbox_address101),
    .ce101(cipher_0_ssbox_ce101),
    .q101(cipher_0_ssbox_q101),
    .address102(cipher_0_ssbox_address102),
    .ce102(cipher_0_ssbox_ce102),
    .q102(cipher_0_ssbox_q102),
    .address103(cipher_0_ssbox_address103),
    .ce103(cipher_0_ssbox_ce103),
    .q103(cipher_0_ssbox_q103),
    .address104(cipher_0_ssbox_address104),
    .ce104(cipher_0_ssbox_ce104),
    .q104(cipher_0_ssbox_q104),
    .address105(cipher_0_ssbox_address105),
    .ce105(cipher_0_ssbox_ce105),
    .q105(cipher_0_ssbox_q105),
    .address106(cipher_0_ssbox_address106),
    .ce106(cipher_0_ssbox_ce106),
    .q106(cipher_0_ssbox_q106),
    .address107(cipher_0_ssbox_address107),
    .ce107(cipher_0_ssbox_ce107),
    .q107(cipher_0_ssbox_q107),
    .address108(cipher_0_ssbox_address108),
    .ce108(cipher_0_ssbox_ce108),
    .q108(cipher_0_ssbox_q108),
    .address109(cipher_0_ssbox_address109),
    .ce109(cipher_0_ssbox_ce109),
    .q109(cipher_0_ssbox_q109),
    .address110(cipher_0_ssbox_address110),
    .ce110(cipher_0_ssbox_ce110),
    .q110(cipher_0_ssbox_q110),
    .address111(cipher_0_ssbox_address111),
    .ce111(cipher_0_ssbox_ce111),
    .q111(cipher_0_ssbox_q111),
    .address112(cipher_0_ssbox_address112),
    .ce112(cipher_0_ssbox_ce112),
    .q112(cipher_0_ssbox_q112),
    .address113(cipher_0_ssbox_address113),
    .ce113(cipher_0_ssbox_ce113),
    .q113(cipher_0_ssbox_q113),
    .address114(cipher_0_ssbox_address114),
    .ce114(cipher_0_ssbox_ce114),
    .q114(cipher_0_ssbox_q114),
    .address115(cipher_0_ssbox_address115),
    .ce115(cipher_0_ssbox_ce115),
    .q115(cipher_0_ssbox_q115),
    .address116(cipher_0_ssbox_address116),
    .ce116(cipher_0_ssbox_ce116),
    .q116(cipher_0_ssbox_q116),
    .address117(cipher_0_ssbox_address117),
    .ce117(cipher_0_ssbox_ce117),
    .q117(cipher_0_ssbox_q117),
    .address118(cipher_0_ssbox_address118),
    .ce118(cipher_0_ssbox_ce118),
    .q118(cipher_0_ssbox_q118),
    .address119(cipher_0_ssbox_address119),
    .ce119(cipher_0_ssbox_ce119),
    .q119(cipher_0_ssbox_q119),
    .address120(cipher_0_ssbox_address120),
    .ce120(cipher_0_ssbox_ce120),
    .q120(cipher_0_ssbox_q120),
    .address121(cipher_0_ssbox_address121),
    .ce121(cipher_0_ssbox_ce121),
    .q121(cipher_0_ssbox_q121),
    .address122(cipher_0_ssbox_address122),
    .ce122(cipher_0_ssbox_ce122),
    .q122(cipher_0_ssbox_q122),
    .address123(cipher_0_ssbox_address123),
    .ce123(cipher_0_ssbox_ce123),
    .q123(cipher_0_ssbox_q123),
    .address124(cipher_0_ssbox_address124),
    .ce124(cipher_0_ssbox_ce124),
    .q124(cipher_0_ssbox_q124),
    .address125(cipher_0_ssbox_address125),
    .ce125(cipher_0_ssbox_ce125),
    .q125(cipher_0_ssbox_q125),
    .address126(cipher_0_ssbox_address126),
    .ce126(cipher_0_ssbox_ce126),
    .q126(cipher_0_ssbox_q126),
    .address127(cipher_0_ssbox_address127),
    .ce127(cipher_0_ssbox_ce127),
    .q127(cipher_0_ssbox_q127),
    .address128(cipher_0_ssbox_address128),
    .ce128(cipher_0_ssbox_ce128),
    .q128(cipher_0_ssbox_q128),
    .address129(cipher_0_ssbox_address129),
    .ce129(cipher_0_ssbox_ce129),
    .q129(cipher_0_ssbox_q129),
    .address130(cipher_0_ssbox_address130),
    .ce130(cipher_0_ssbox_ce130),
    .q130(cipher_0_ssbox_q130),
    .address131(cipher_0_ssbox_address131),
    .ce131(cipher_0_ssbox_ce131),
    .q131(cipher_0_ssbox_q131),
    .address132(cipher_0_ssbox_address132),
    .ce132(cipher_0_ssbox_ce132),
    .q132(cipher_0_ssbox_q132),
    .address133(cipher_0_ssbox_address133),
    .ce133(cipher_0_ssbox_ce133),
    .q133(cipher_0_ssbox_q133),
    .address134(cipher_0_ssbox_address134),
    .ce134(cipher_0_ssbox_ce134),
    .q134(cipher_0_ssbox_q134),
    .address135(cipher_0_ssbox_address135),
    .ce135(cipher_0_ssbox_ce135),
    .q135(cipher_0_ssbox_q135),
    .address136(cipher_0_ssbox_address136),
    .ce136(cipher_0_ssbox_ce136),
    .q136(cipher_0_ssbox_q136),
    .address137(cipher_0_ssbox_address137),
    .ce137(cipher_0_ssbox_ce137),
    .q137(cipher_0_ssbox_q137),
    .address138(cipher_0_ssbox_address138),
    .ce138(cipher_0_ssbox_ce138),
    .q138(cipher_0_ssbox_q138),
    .address139(cipher_0_ssbox_address139),
    .ce139(cipher_0_ssbox_ce139),
    .q139(cipher_0_ssbox_q139),
    .address140(cipher_0_ssbox_address140),
    .ce140(cipher_0_ssbox_ce140),
    .q140(cipher_0_ssbox_q140),
    .address141(cipher_0_ssbox_address141),
    .ce141(cipher_0_ssbox_ce141),
    .q141(cipher_0_ssbox_q141),
    .address142(cipher_0_ssbox_address142),
    .ce142(cipher_0_ssbox_ce142),
    .q142(cipher_0_ssbox_q142),
    .address143(cipher_0_ssbox_address143),
    .ce143(cipher_0_ssbox_ce143),
    .q143(cipher_0_ssbox_q143),
    .address144(cipher_0_ssbox_address144),
    .ce144(cipher_0_ssbox_ce144),
    .q144(cipher_0_ssbox_q144),
    .address145(cipher_0_ssbox_address145),
    .ce145(cipher_0_ssbox_ce145),
    .q145(cipher_0_ssbox_q145),
    .address146(cipher_0_ssbox_address146),
    .ce146(cipher_0_ssbox_ce146),
    .q146(cipher_0_ssbox_q146),
    .address147(cipher_0_ssbox_address147),
    .ce147(cipher_0_ssbox_ce147),
    .q147(cipher_0_ssbox_q147),
    .address148(cipher_0_ssbox_address148),
    .ce148(cipher_0_ssbox_ce148),
    .q148(cipher_0_ssbox_q148),
    .address149(cipher_0_ssbox_address149),
    .ce149(cipher_0_ssbox_ce149),
    .q149(cipher_0_ssbox_q149),
    .address150(cipher_0_ssbox_address150),
    .ce150(cipher_0_ssbox_ce150),
    .q150(cipher_0_ssbox_q150),
    .address151(cipher_0_ssbox_address151),
    .ce151(cipher_0_ssbox_ce151),
    .q151(cipher_0_ssbox_q151),
    .address152(cipher_0_ssbox_address152),
    .ce152(cipher_0_ssbox_ce152),
    .q152(cipher_0_ssbox_q152),
    .address153(cipher_0_ssbox_address153),
    .ce153(cipher_0_ssbox_ce153),
    .q153(cipher_0_ssbox_q153),
    .address154(cipher_0_ssbox_address154),
    .ce154(cipher_0_ssbox_ce154),
    .q154(cipher_0_ssbox_q154),
    .address155(cipher_0_ssbox_address155),
    .ce155(cipher_0_ssbox_ce155),
    .q155(cipher_0_ssbox_q155),
    .address156(cipher_0_ssbox_address156),
    .ce156(cipher_0_ssbox_ce156),
    .q156(cipher_0_ssbox_q156),
    .address157(cipher_0_ssbox_address157),
    .ce157(cipher_0_ssbox_ce157),
    .q157(cipher_0_ssbox_q157),
    .address158(cipher_0_ssbox_address158),
    .ce158(cipher_0_ssbox_ce158),
    .q158(cipher_0_ssbox_q158),
    .address159(cipher_0_ssbox_address159),
    .ce159(cipher_0_ssbox_ce159),
    .q159(cipher_0_ssbox_q159),
    .address160(cipher_0_ssbox_address160),
    .ce160(cipher_0_ssbox_ce160),
    .q160(cipher_0_ssbox_q160),
    .address161(cipher_0_ssbox_address161),
    .ce161(cipher_0_ssbox_ce161),
    .q161(cipher_0_ssbox_q161),
    .address162(cipher_0_ssbox_address162),
    .ce162(cipher_0_ssbox_ce162),
    .q162(cipher_0_ssbox_q162),
    .address163(cipher_0_ssbox_address163),
    .ce163(cipher_0_ssbox_ce163),
    .q163(cipher_0_ssbox_q163),
    .address164(cipher_0_ssbox_address164),
    .ce164(cipher_0_ssbox_ce164),
    .q164(cipher_0_ssbox_q164),
    .address165(cipher_0_ssbox_address165),
    .ce165(cipher_0_ssbox_ce165),
    .q165(cipher_0_ssbox_q165),
    .address166(cipher_0_ssbox_address166),
    .ce166(cipher_0_ssbox_ce166),
    .q166(cipher_0_ssbox_q166),
    .address167(cipher_0_ssbox_address167),
    .ce167(cipher_0_ssbox_ce167),
    .q167(cipher_0_ssbox_q167),
    .address168(cipher_0_ssbox_address168),
    .ce168(cipher_0_ssbox_ce168),
    .q168(cipher_0_ssbox_q168),
    .address169(cipher_0_ssbox_address169),
    .ce169(cipher_0_ssbox_ce169),
    .q169(cipher_0_ssbox_q169),
    .address170(cipher_0_ssbox_address170),
    .ce170(cipher_0_ssbox_ce170),
    .q170(cipher_0_ssbox_q170),
    .address171(cipher_0_ssbox_address171),
    .ce171(cipher_0_ssbox_ce171),
    .q171(cipher_0_ssbox_q171),
    .address172(cipher_0_ssbox_address172),
    .ce172(cipher_0_ssbox_ce172),
    .q172(cipher_0_ssbox_q172),
    .address173(cipher_0_ssbox_address173),
    .ce173(cipher_0_ssbox_ce173),
    .q173(cipher_0_ssbox_q173),
    .address174(cipher_0_ssbox_address174),
    .ce174(cipher_0_ssbox_ce174),
    .q174(cipher_0_ssbox_q174),
    .address175(cipher_0_ssbox_address175),
    .ce175(cipher_0_ssbox_ce175),
    .q175(cipher_0_ssbox_q175),
    .address176(cipher_0_ssbox_address176),
    .ce176(cipher_0_ssbox_ce176),
    .q176(cipher_0_ssbox_q176),
    .address177(cipher_0_ssbox_address177),
    .ce177(cipher_0_ssbox_ce177),
    .q177(cipher_0_ssbox_q177),
    .address178(cipher_0_ssbox_address178),
    .ce178(cipher_0_ssbox_ce178),
    .q178(cipher_0_ssbox_q178),
    .address179(cipher_0_ssbox_address179),
    .ce179(cipher_0_ssbox_ce179),
    .q179(cipher_0_ssbox_q179),
    .address180(cipher_0_ssbox_address180),
    .ce180(cipher_0_ssbox_ce180),
    .q180(cipher_0_ssbox_q180),
    .address181(cipher_0_ssbox_address181),
    .ce181(cipher_0_ssbox_ce181),
    .q181(cipher_0_ssbox_q181),
    .address182(cipher_0_ssbox_address182),
    .ce182(cipher_0_ssbox_ce182),
    .q182(cipher_0_ssbox_q182),
    .address183(cipher_0_ssbox_address183),
    .ce183(cipher_0_ssbox_ce183),
    .q183(cipher_0_ssbox_q183),
    .address184(cipher_0_ssbox_address184),
    .ce184(cipher_0_ssbox_ce184),
    .q184(cipher_0_ssbox_q184),
    .address185(cipher_0_ssbox_address185),
    .ce185(cipher_0_ssbox_ce185),
    .q185(cipher_0_ssbox_q185),
    .address186(cipher_0_ssbox_address186),
    .ce186(cipher_0_ssbox_ce186),
    .q186(cipher_0_ssbox_q186),
    .address187(cipher_0_ssbox_address187),
    .ce187(cipher_0_ssbox_ce187),
    .q187(cipher_0_ssbox_q187),
    .address188(cipher_0_ssbox_address188),
    .ce188(cipher_0_ssbox_ce188),
    .q188(cipher_0_ssbox_q188),
    .address189(cipher_0_ssbox_address189),
    .ce189(cipher_0_ssbox_ce189),
    .q189(cipher_0_ssbox_q189),
    .address190(cipher_0_ssbox_address190),
    .ce190(cipher_0_ssbox_ce190),
    .q190(cipher_0_ssbox_q190),
    .address191(cipher_0_ssbox_address191),
    .ce191(cipher_0_ssbox_ce191),
    .q191(cipher_0_ssbox_q191)
);

testEnc_process_r_cipher_0_p16box_ROM_NP_LUTRAM_1R #(
    .DataWidth( 16 ),
    .AddressRange( 256 ),
    .AddressWidth( 8 ))
cipher_0_p16box_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(cipher_0_p16box_address0),
    .ce0(cipher_0_p16box_ce0),
    .q0(cipher_0_p16box_q0),
    .address1(cipher_0_p16box_address1),
    .ce1(cipher_0_p16box_ce1),
    .q1(cipher_0_p16box_q1),
    .address2(cipher_0_p16box_address2),
    .ce2(cipher_0_p16box_ce2),
    .q2(cipher_0_p16box_q2),
    .address3(cipher_0_p16box_address3),
    .ce3(cipher_0_p16box_ce3),
    .q3(cipher_0_p16box_q3),
    .address4(cipher_0_p16box_address4),
    .ce4(cipher_0_p16box_ce4),
    .q4(cipher_0_p16box_q4),
    .address5(cipher_0_p16box_address5),
    .ce5(cipher_0_p16box_ce5),
    .q5(cipher_0_p16box_q5),
    .address6(cipher_0_p16box_address6),
    .ce6(cipher_0_p16box_ce6),
    .q6(cipher_0_p16box_q6),
    .address7(cipher_0_p16box_address7),
    .ce7(cipher_0_p16box_ce7),
    .q7(cipher_0_p16box_q7),
    .address8(cipher_0_p16box_address8),
    .ce8(cipher_0_p16box_ce8),
    .q8(cipher_0_p16box_q8),
    .address9(cipher_0_p16box_address9),
    .ce9(cipher_0_p16box_ce9),
    .q9(cipher_0_p16box_q9),
    .address10(cipher_0_p16box_address10),
    .ce10(cipher_0_p16box_ce10),
    .q10(cipher_0_p16box_q10),
    .address11(cipher_0_p16box_address11),
    .ce11(cipher_0_p16box_ce11),
    .q11(cipher_0_p16box_q11),
    .address12(cipher_0_p16box_address12),
    .ce12(cipher_0_p16box_ce12),
    .q12(cipher_0_p16box_q12),
    .address13(cipher_0_p16box_address13),
    .ce13(cipher_0_p16box_ce13),
    .q13(cipher_0_p16box_q13),
    .address14(cipher_0_p16box_address14),
    .ce14(cipher_0_p16box_ce14),
    .q14(cipher_0_p16box_q14),
    .address15(cipher_0_p16box_address15),
    .ce15(cipher_0_p16box_ce15),
    .q15(cipher_0_p16box_q15),
    .address16(cipher_0_p16box_address16),
    .ce16(cipher_0_p16box_ce16),
    .q16(cipher_0_p16box_q16),
    .address17(cipher_0_p16box_address17),
    .ce17(cipher_0_p16box_ce17),
    .q17(cipher_0_p16box_q17),
    .address18(cipher_0_p16box_address18),
    .ce18(cipher_0_p16box_ce18),
    .q18(cipher_0_p16box_q18),
    .address19(cipher_0_p16box_address19),
    .ce19(cipher_0_p16box_ce19),
    .q19(cipher_0_p16box_q19),
    .address20(cipher_0_p16box_address20),
    .ce20(cipher_0_p16box_ce20),
    .q20(cipher_0_p16box_q20),
    .address21(cipher_0_p16box_address21),
    .ce21(cipher_0_p16box_ce21),
    .q21(cipher_0_p16box_q21),
    .address22(cipher_0_p16box_address22),
    .ce22(cipher_0_p16box_ce22),
    .q22(cipher_0_p16box_q22),
    .address23(cipher_0_p16box_address23),
    .ce23(cipher_0_p16box_ce23),
    .q23(cipher_0_p16box_q23),
    .address24(cipher_0_p16box_address24),
    .ce24(cipher_0_p16box_ce24),
    .q24(cipher_0_p16box_q24),
    .address25(cipher_0_p16box_address25),
    .ce25(cipher_0_p16box_ce25),
    .q25(cipher_0_p16box_q25),
    .address26(cipher_0_p16box_address26),
    .ce26(cipher_0_p16box_ce26),
    .q26(cipher_0_p16box_q26),
    .address27(cipher_0_p16box_address27),
    .ce27(cipher_0_p16box_ce27),
    .q27(cipher_0_p16box_q27),
    .address28(cipher_0_p16box_address28),
    .ce28(cipher_0_p16box_ce28),
    .q28(cipher_0_p16box_q28),
    .address29(cipher_0_p16box_address29),
    .ce29(cipher_0_p16box_ce29),
    .q29(cipher_0_p16box_q29),
    .address30(cipher_0_p16box_address30),
    .ce30(cipher_0_p16box_ce30),
    .q30(cipher_0_p16box_q30),
    .address31(cipher_0_p16box_address31),
    .ce31(cipher_0_p16box_ce31),
    .q31(cipher_0_p16box_q31),
    .address32(cipher_0_p16box_address32),
    .ce32(cipher_0_p16box_ce32),
    .q32(cipher_0_p16box_q32),
    .address33(cipher_0_p16box_address33),
    .ce33(cipher_0_p16box_ce33),
    .q33(cipher_0_p16box_q33),
    .address34(cipher_0_p16box_address34),
    .ce34(cipher_0_p16box_ce34),
    .q34(cipher_0_p16box_q34),
    .address35(cipher_0_p16box_address35),
    .ce35(cipher_0_p16box_ce35),
    .q35(cipher_0_p16box_q35),
    .address36(cipher_0_p16box_address36),
    .ce36(cipher_0_p16box_ce36),
    .q36(cipher_0_p16box_q36),
    .address37(cipher_0_p16box_address37),
    .ce37(cipher_0_p16box_ce37),
    .q37(cipher_0_p16box_q37),
    .address38(cipher_0_p16box_address38),
    .ce38(cipher_0_p16box_ce38),
    .q38(cipher_0_p16box_q38),
    .address39(cipher_0_p16box_address39),
    .ce39(cipher_0_p16box_ce39),
    .q39(cipher_0_p16box_q39),
    .address40(cipher_0_p16box_address40),
    .ce40(cipher_0_p16box_ce40),
    .q40(cipher_0_p16box_q40),
    .address41(cipher_0_p16box_address41),
    .ce41(cipher_0_p16box_ce41),
    .q41(cipher_0_p16box_q41),
    .address42(cipher_0_p16box_address42),
    .ce42(cipher_0_p16box_ce42),
    .q42(cipher_0_p16box_q42),
    .address43(cipher_0_p16box_address43),
    .ce43(cipher_0_p16box_ce43),
    .q43(cipher_0_p16box_q43),
    .address44(cipher_0_p16box_address44),
    .ce44(cipher_0_p16box_ce44),
    .q44(cipher_0_p16box_q44),
    .address45(cipher_0_p16box_address45),
    .ce45(cipher_0_p16box_ce45),
    .q45(cipher_0_p16box_q45),
    .address46(cipher_0_p16box_address46),
    .ce46(cipher_0_p16box_ce46),
    .q46(cipher_0_p16box_q46),
    .address47(cipher_0_p16box_address47),
    .ce47(cipher_0_p16box_ce47),
    .q47(cipher_0_p16box_q47),
    .address48(cipher_0_p16box_address48),
    .ce48(cipher_0_p16box_ce48),
    .q48(cipher_0_p16box_q48),
    .address49(cipher_0_p16box_address49),
    .ce49(cipher_0_p16box_ce49),
    .q49(cipher_0_p16box_q49),
    .address50(cipher_0_p16box_address50),
    .ce50(cipher_0_p16box_ce50),
    .q50(cipher_0_p16box_q50),
    .address51(cipher_0_p16box_address51),
    .ce51(cipher_0_p16box_ce51),
    .q51(cipher_0_p16box_q51),
    .address52(cipher_0_p16box_address52),
    .ce52(cipher_0_p16box_ce52),
    .q52(cipher_0_p16box_q52),
    .address53(cipher_0_p16box_address53),
    .ce53(cipher_0_p16box_ce53),
    .q53(cipher_0_p16box_q53),
    .address54(cipher_0_p16box_address54),
    .ce54(cipher_0_p16box_ce54),
    .q54(cipher_0_p16box_q54),
    .address55(cipher_0_p16box_address55),
    .ce55(cipher_0_p16box_ce55),
    .q55(cipher_0_p16box_q55),
    .address56(cipher_0_p16box_address56),
    .ce56(cipher_0_p16box_ce56),
    .q56(cipher_0_p16box_q56),
    .address57(cipher_0_p16box_address57),
    .ce57(cipher_0_p16box_ce57),
    .q57(cipher_0_p16box_q57),
    .address58(cipher_0_p16box_address58),
    .ce58(cipher_0_p16box_ce58),
    .q58(cipher_0_p16box_q58),
    .address59(cipher_0_p16box_address59),
    .ce59(cipher_0_p16box_ce59),
    .q59(cipher_0_p16box_q59),
    .address60(cipher_0_p16box_address60),
    .ce60(cipher_0_p16box_ce60),
    .q60(cipher_0_p16box_q60),
    .address61(cipher_0_p16box_address61),
    .ce61(cipher_0_p16box_ce61),
    .q61(cipher_0_p16box_q61),
    .address62(cipher_0_p16box_address62),
    .ce62(cipher_0_p16box_ce62),
    .q62(cipher_0_p16box_q62),
    .address63(cipher_0_p16box_address63),
    .ce63(cipher_0_p16box_ce63),
    .q63(cipher_0_p16box_q63),
    .address64(cipher_0_p16box_address64),
    .ce64(cipher_0_p16box_ce64),
    .q64(cipher_0_p16box_q64),
    .address65(cipher_0_p16box_address65),
    .ce65(cipher_0_p16box_ce65),
    .q65(cipher_0_p16box_q65),
    .address66(cipher_0_p16box_address66),
    .ce66(cipher_0_p16box_ce66),
    .q66(cipher_0_p16box_q66),
    .address67(cipher_0_p16box_address67),
    .ce67(cipher_0_p16box_ce67),
    .q67(cipher_0_p16box_q67),
    .address68(cipher_0_p16box_address68),
    .ce68(cipher_0_p16box_ce68),
    .q68(cipher_0_p16box_q68),
    .address69(cipher_0_p16box_address69),
    .ce69(cipher_0_p16box_ce69),
    .q69(cipher_0_p16box_q69),
    .address70(cipher_0_p16box_address70),
    .ce70(cipher_0_p16box_ce70),
    .q70(cipher_0_p16box_q70),
    .address71(cipher_0_p16box_address71),
    .ce71(cipher_0_p16box_ce71),
    .q71(cipher_0_p16box_q71),
    .address72(cipher_0_p16box_address72),
    .ce72(cipher_0_p16box_ce72),
    .q72(cipher_0_p16box_q72),
    .address73(cipher_0_p16box_address73),
    .ce73(cipher_0_p16box_ce73),
    .q73(cipher_0_p16box_q73),
    .address74(cipher_0_p16box_address74),
    .ce74(cipher_0_p16box_ce74),
    .q74(cipher_0_p16box_q74),
    .address75(cipher_0_p16box_address75),
    .ce75(cipher_0_p16box_ce75),
    .q75(cipher_0_p16box_q75),
    .address76(cipher_0_p16box_address76),
    .ce76(cipher_0_p16box_ce76),
    .q76(cipher_0_p16box_q76),
    .address77(cipher_0_p16box_address77),
    .ce77(cipher_0_p16box_ce77),
    .q77(cipher_0_p16box_q77),
    .address78(cipher_0_p16box_address78),
    .ce78(cipher_0_p16box_ce78),
    .q78(cipher_0_p16box_q78),
    .address79(cipher_0_p16box_address79),
    .ce79(cipher_0_p16box_ce79),
    .q79(cipher_0_p16box_q79),
    .address80(cipher_0_p16box_address80),
    .ce80(cipher_0_p16box_ce80),
    .q80(cipher_0_p16box_q80),
    .address81(cipher_0_p16box_address81),
    .ce81(cipher_0_p16box_ce81),
    .q81(cipher_0_p16box_q81),
    .address82(cipher_0_p16box_address82),
    .ce82(cipher_0_p16box_ce82),
    .q82(cipher_0_p16box_q82),
    .address83(cipher_0_p16box_address83),
    .ce83(cipher_0_p16box_ce83),
    .q83(cipher_0_p16box_q83),
    .address84(cipher_0_p16box_address84),
    .ce84(cipher_0_p16box_ce84),
    .q84(cipher_0_p16box_q84),
    .address85(cipher_0_p16box_address85),
    .ce85(cipher_0_p16box_ce85),
    .q85(cipher_0_p16box_q85),
    .address86(cipher_0_p16box_address86),
    .ce86(cipher_0_p16box_ce86),
    .q86(cipher_0_p16box_q86),
    .address87(cipher_0_p16box_address87),
    .ce87(cipher_0_p16box_ce87),
    .q87(cipher_0_p16box_q87),
    .address88(cipher_0_p16box_address88),
    .ce88(cipher_0_p16box_ce88),
    .q88(cipher_0_p16box_q88),
    .address89(cipher_0_p16box_address89),
    .ce89(cipher_0_p16box_ce89),
    .q89(cipher_0_p16box_q89),
    .address90(cipher_0_p16box_address90),
    .ce90(cipher_0_p16box_ce90),
    .q90(cipher_0_p16box_q90),
    .address91(cipher_0_p16box_address91),
    .ce91(cipher_0_p16box_ce91),
    .q91(cipher_0_p16box_q91),
    .address92(cipher_0_p16box_address92),
    .ce92(cipher_0_p16box_ce92),
    .q92(cipher_0_p16box_q92),
    .address93(cipher_0_p16box_address93),
    .ce93(cipher_0_p16box_ce93),
    .q93(cipher_0_p16box_q93),
    .address94(cipher_0_p16box_address94),
    .ce94(cipher_0_p16box_ce94),
    .q94(cipher_0_p16box_q94),
    .address95(cipher_0_p16box_address95),
    .ce95(cipher_0_p16box_ce95),
    .q95(cipher_0_p16box_q95),
    .address96(cipher_0_p16box_address96),
    .ce96(cipher_0_p16box_ce96),
    .q96(cipher_0_p16box_q96),
    .address97(cipher_0_p16box_address97),
    .ce97(cipher_0_p16box_ce97),
    .q97(cipher_0_p16box_q97),
    .address98(cipher_0_p16box_address98),
    .ce98(cipher_0_p16box_ce98),
    .q98(cipher_0_p16box_q98),
    .address99(cipher_0_p16box_address99),
    .ce99(cipher_0_p16box_ce99),
    .q99(cipher_0_p16box_q99),
    .address100(cipher_0_p16box_address100),
    .ce100(cipher_0_p16box_ce100),
    .q100(cipher_0_p16box_q100),
    .address101(cipher_0_p16box_address101),
    .ce101(cipher_0_p16box_ce101),
    .q101(cipher_0_p16box_q101),
    .address102(cipher_0_p16box_address102),
    .ce102(cipher_0_p16box_ce102),
    .q102(cipher_0_p16box_q102),
    .address103(cipher_0_p16box_address103),
    .ce103(cipher_0_p16box_ce103),
    .q103(cipher_0_p16box_q103),
    .address104(cipher_0_p16box_address104),
    .ce104(cipher_0_p16box_ce104),
    .q104(cipher_0_p16box_q104),
    .address105(cipher_0_p16box_address105),
    .ce105(cipher_0_p16box_ce105),
    .q105(cipher_0_p16box_q105),
    .address106(cipher_0_p16box_address106),
    .ce106(cipher_0_p16box_ce106),
    .q106(cipher_0_p16box_q106),
    .address107(cipher_0_p16box_address107),
    .ce107(cipher_0_p16box_ce107),
    .q107(cipher_0_p16box_q107),
    .address108(cipher_0_p16box_address108),
    .ce108(cipher_0_p16box_ce108),
    .q108(cipher_0_p16box_q108),
    .address109(cipher_0_p16box_address109),
    .ce109(cipher_0_p16box_ce109),
    .q109(cipher_0_p16box_q109),
    .address110(cipher_0_p16box_address110),
    .ce110(cipher_0_p16box_ce110),
    .q110(cipher_0_p16box_q110),
    .address111(cipher_0_p16box_address111),
    .ce111(cipher_0_p16box_ce111),
    .q111(cipher_0_p16box_q111),
    .address112(cipher_0_p16box_address112),
    .ce112(cipher_0_p16box_ce112),
    .q112(cipher_0_p16box_q112),
    .address113(cipher_0_p16box_address113),
    .ce113(cipher_0_p16box_ce113),
    .q113(cipher_0_p16box_q113),
    .address114(cipher_0_p16box_address114),
    .ce114(cipher_0_p16box_ce114),
    .q114(cipher_0_p16box_q114),
    .address115(cipher_0_p16box_address115),
    .ce115(cipher_0_p16box_ce115),
    .q115(cipher_0_p16box_q115),
    .address116(cipher_0_p16box_address116),
    .ce116(cipher_0_p16box_ce116),
    .q116(cipher_0_p16box_q116),
    .address117(cipher_0_p16box_address117),
    .ce117(cipher_0_p16box_ce117),
    .q117(cipher_0_p16box_q117),
    .address118(cipher_0_p16box_address118),
    .ce118(cipher_0_p16box_ce118),
    .q118(cipher_0_p16box_q118),
    .address119(cipher_0_p16box_address119),
    .ce119(cipher_0_p16box_ce119),
    .q119(cipher_0_p16box_q119),
    .address120(cipher_0_p16box_address120),
    .ce120(cipher_0_p16box_ce120),
    .q120(cipher_0_p16box_q120),
    .address121(cipher_0_p16box_address121),
    .ce121(cipher_0_p16box_ce121),
    .q121(cipher_0_p16box_q121),
    .address122(cipher_0_p16box_address122),
    .ce122(cipher_0_p16box_ce122),
    .q122(cipher_0_p16box_q122),
    .address123(cipher_0_p16box_address123),
    .ce123(cipher_0_p16box_ce123),
    .q123(cipher_0_p16box_q123),
    .address124(cipher_0_p16box_address124),
    .ce124(cipher_0_p16box_ce124),
    .q124(cipher_0_p16box_q124),
    .address125(cipher_0_p16box_address125),
    .ce125(cipher_0_p16box_ce125),
    .q125(cipher_0_p16box_q125),
    .address126(cipher_0_p16box_address126),
    .ce126(cipher_0_p16box_ce126),
    .q126(cipher_0_p16box_q126),
    .address127(cipher_0_p16box_address127),
    .ce127(cipher_0_p16box_ce127),
    .q127(cipher_0_p16box_q127),
    .address128(cipher_0_p16box_address128),
    .ce128(cipher_0_p16box_ce128),
    .q128(cipher_0_p16box_q128),
    .address129(cipher_0_p16box_address129),
    .ce129(cipher_0_p16box_ce129),
    .q129(cipher_0_p16box_q129),
    .address130(cipher_0_p16box_address130),
    .ce130(cipher_0_p16box_ce130),
    .q130(cipher_0_p16box_q130),
    .address131(cipher_0_p16box_address131),
    .ce131(cipher_0_p16box_ce131),
    .q131(cipher_0_p16box_q131),
    .address132(cipher_0_p16box_address132),
    .ce132(cipher_0_p16box_ce132),
    .q132(cipher_0_p16box_q132),
    .address133(cipher_0_p16box_address133),
    .ce133(cipher_0_p16box_ce133),
    .q133(cipher_0_p16box_q133),
    .address134(cipher_0_p16box_address134),
    .ce134(cipher_0_p16box_ce134),
    .q134(cipher_0_p16box_q134),
    .address135(cipher_0_p16box_address135),
    .ce135(cipher_0_p16box_ce135),
    .q135(cipher_0_p16box_q135),
    .address136(cipher_0_p16box_address136),
    .ce136(cipher_0_p16box_ce136),
    .q136(cipher_0_p16box_q136),
    .address137(cipher_0_p16box_address137),
    .ce137(cipher_0_p16box_ce137),
    .q137(cipher_0_p16box_q137),
    .address138(cipher_0_p16box_address138),
    .ce138(cipher_0_p16box_ce138),
    .q138(cipher_0_p16box_q138),
    .address139(cipher_0_p16box_address139),
    .ce139(cipher_0_p16box_ce139),
    .q139(cipher_0_p16box_q139),
    .address140(cipher_0_p16box_address140),
    .ce140(cipher_0_p16box_ce140),
    .q140(cipher_0_p16box_q140),
    .address141(cipher_0_p16box_address141),
    .ce141(cipher_0_p16box_ce141),
    .q141(cipher_0_p16box_q141),
    .address142(cipher_0_p16box_address142),
    .ce142(cipher_0_p16box_ce142),
    .q142(cipher_0_p16box_q142),
    .address143(cipher_0_p16box_address143),
    .ce143(cipher_0_p16box_ce143),
    .q143(cipher_0_p16box_q143),
    .address144(cipher_0_p16box_address144),
    .ce144(cipher_0_p16box_ce144),
    .q144(cipher_0_p16box_q144),
    .address145(cipher_0_p16box_address145),
    .ce145(cipher_0_p16box_ce145),
    .q145(cipher_0_p16box_q145),
    .address146(cipher_0_p16box_address146),
    .ce146(cipher_0_p16box_ce146),
    .q146(cipher_0_p16box_q146),
    .address147(cipher_0_p16box_address147),
    .ce147(cipher_0_p16box_ce147),
    .q147(cipher_0_p16box_q147),
    .address148(cipher_0_p16box_address148),
    .ce148(cipher_0_p16box_ce148),
    .q148(cipher_0_p16box_q148),
    .address149(cipher_0_p16box_address149),
    .ce149(cipher_0_p16box_ce149),
    .q149(cipher_0_p16box_q149),
    .address150(cipher_0_p16box_address150),
    .ce150(cipher_0_p16box_ce150),
    .q150(cipher_0_p16box_q150),
    .address151(cipher_0_p16box_address151),
    .ce151(cipher_0_p16box_ce151),
    .q151(cipher_0_p16box_q151),
    .address152(cipher_0_p16box_address152),
    .ce152(cipher_0_p16box_ce152),
    .q152(cipher_0_p16box_q152),
    .address153(cipher_0_p16box_address153),
    .ce153(cipher_0_p16box_ce153),
    .q153(cipher_0_p16box_q153),
    .address154(cipher_0_p16box_address154),
    .ce154(cipher_0_p16box_ce154),
    .q154(cipher_0_p16box_q154),
    .address155(cipher_0_p16box_address155),
    .ce155(cipher_0_p16box_ce155),
    .q155(cipher_0_p16box_q155),
    .address156(cipher_0_p16box_address156),
    .ce156(cipher_0_p16box_ce156),
    .q156(cipher_0_p16box_q156),
    .address157(cipher_0_p16box_address157),
    .ce157(cipher_0_p16box_ce157),
    .q157(cipher_0_p16box_q157),
    .address158(cipher_0_p16box_address158),
    .ce158(cipher_0_p16box_ce158),
    .q158(cipher_0_p16box_q158),
    .address159(cipher_0_p16box_address159),
    .ce159(cipher_0_p16box_ce159),
    .q159(cipher_0_p16box_q159),
    .address160(cipher_0_p16box_address160),
    .ce160(cipher_0_p16box_ce160),
    .q160(cipher_0_p16box_q160),
    .address161(cipher_0_p16box_address161),
    .ce161(cipher_0_p16box_ce161),
    .q161(cipher_0_p16box_q161),
    .address162(cipher_0_p16box_address162),
    .ce162(cipher_0_p16box_ce162),
    .q162(cipher_0_p16box_q162),
    .address163(cipher_0_p16box_address163),
    .ce163(cipher_0_p16box_ce163),
    .q163(cipher_0_p16box_q163),
    .address164(cipher_0_p16box_address164),
    .ce164(cipher_0_p16box_ce164),
    .q164(cipher_0_p16box_q164),
    .address165(cipher_0_p16box_address165),
    .ce165(cipher_0_p16box_ce165),
    .q165(cipher_0_p16box_q165),
    .address166(cipher_0_p16box_address166),
    .ce166(cipher_0_p16box_ce166),
    .q166(cipher_0_p16box_q166),
    .address167(cipher_0_p16box_address167),
    .ce167(cipher_0_p16box_ce167),
    .q167(cipher_0_p16box_q167),
    .address168(cipher_0_p16box_address168),
    .ce168(cipher_0_p16box_ce168),
    .q168(cipher_0_p16box_q168),
    .address169(cipher_0_p16box_address169),
    .ce169(cipher_0_p16box_ce169),
    .q169(cipher_0_p16box_q169),
    .address170(cipher_0_p16box_address170),
    .ce170(cipher_0_p16box_ce170),
    .q170(cipher_0_p16box_q170),
    .address171(cipher_0_p16box_address171),
    .ce171(cipher_0_p16box_ce171),
    .q171(cipher_0_p16box_q171),
    .address172(cipher_0_p16box_address172),
    .ce172(cipher_0_p16box_ce172),
    .q172(cipher_0_p16box_q172),
    .address173(cipher_0_p16box_address173),
    .ce173(cipher_0_p16box_ce173),
    .q173(cipher_0_p16box_q173),
    .address174(cipher_0_p16box_address174),
    .ce174(cipher_0_p16box_ce174),
    .q174(cipher_0_p16box_q174),
    .address175(cipher_0_p16box_address175),
    .ce175(cipher_0_p16box_ce175),
    .q175(cipher_0_p16box_q175)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_enable_reg_pp0_iter1 <= ap_start;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter10 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter10 <= ap_enable_reg_pp0_iter9;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter11 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter11 <= ap_enable_reg_pp0_iter10;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter12 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter12 <= ap_enable_reg_pp0_iter11;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter13 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter13 <= ap_enable_reg_pp0_iter12;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter14 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter14 <= ap_enable_reg_pp0_iter13;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter15 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter15 <= ap_enable_reg_pp0_iter14;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter16 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter16 <= ap_enable_reg_pp0_iter15;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter17 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter17 <= ap_enable_reg_pp0_iter16;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter18 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter18 <= ap_enable_reg_pp0_iter17;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter19 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter19 <= ap_enable_reg_pp0_iter18;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter20 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter20 <= ap_enable_reg_pp0_iter19;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter21 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter21 <= ap_enable_reg_pp0_iter20;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter22 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter22 <= ap_enable_reg_pp0_iter21;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter23 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter23 <= ap_enable_reg_pp0_iter22;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter5 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter6 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter7 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter8 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter8 <= ap_enable_reg_pp0_iter7;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter9 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter9 <= ap_enable_reg_pp0_iter8;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        p_read_10_reg_14123 <= p_read3;
        p_read_10_reg_14123_pp0_iter1_reg <= p_read_10_reg_14123;
        p_read_11_reg_14128 <= p_read2;
        p_read_11_reg_14128_pp0_iter1_reg <= p_read_11_reg_14128;
        p_read_12_reg_14133 <= p_read1;
        p_read_12_reg_14133_pp0_iter1_reg <= p_read_12_reg_14133;
        p_read_1_reg_14078 <= p_read12;
        p_read_1_reg_14078_pp0_iter1_reg <= p_read_1_reg_14078;
        p_read_2_reg_14083 <= p_read11;
        p_read_2_reg_14083_pp0_iter1_reg <= p_read_2_reg_14083;
        p_read_3_reg_14088 <= p_read10;
        p_read_3_reg_14088_pp0_iter1_reg <= p_read_3_reg_14088;
        p_read_4_reg_14093 <= p_read9;
        p_read_4_reg_14093_pp0_iter1_reg <= p_read_4_reg_14093;
        p_read_5_reg_14098 <= p_read8;
        p_read_5_reg_14098_pp0_iter1_reg <= p_read_5_reg_14098;
        p_read_6_reg_14103 <= p_read7;
        p_read_6_reg_14103_pp0_iter1_reg <= p_read_6_reg_14103;
        p_read_7_reg_14108 <= p_read6;
        p_read_7_reg_14108_pp0_iter1_reg <= p_read_7_reg_14108;
        p_read_8_reg_14113 <= p_read5;
        p_read_8_reg_14113_pp0_iter1_reg <= p_read_8_reg_14113;
        p_read_9_reg_14118 <= p_read4;
        p_read_9_reg_14118_pp0_iter1_reg <= p_read_9_reg_14118;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        p_read_10_reg_14123_pp0_iter2_reg <= p_read_10_reg_14123_pp0_iter1_reg;
        p_read_10_reg_14123_pp0_iter3_reg <= p_read_10_reg_14123_pp0_iter2_reg;
        p_read_10_reg_14123_pp0_iter4_reg <= p_read_10_reg_14123_pp0_iter3_reg;
        p_read_10_reg_14123_pp0_iter5_reg <= p_read_10_reg_14123_pp0_iter4_reg;
        p_read_11_reg_14128_pp0_iter2_reg <= p_read_11_reg_14128_pp0_iter1_reg;
        p_read_11_reg_14128_pp0_iter3_reg <= p_read_11_reg_14128_pp0_iter2_reg;
        p_read_1_reg_14078_pp0_iter10_reg <= p_read_1_reg_14078_pp0_iter9_reg;
        p_read_1_reg_14078_pp0_iter11_reg <= p_read_1_reg_14078_pp0_iter10_reg;
        p_read_1_reg_14078_pp0_iter12_reg <= p_read_1_reg_14078_pp0_iter11_reg;
        p_read_1_reg_14078_pp0_iter13_reg <= p_read_1_reg_14078_pp0_iter12_reg;
        p_read_1_reg_14078_pp0_iter14_reg <= p_read_1_reg_14078_pp0_iter13_reg;
        p_read_1_reg_14078_pp0_iter15_reg <= p_read_1_reg_14078_pp0_iter14_reg;
        p_read_1_reg_14078_pp0_iter16_reg <= p_read_1_reg_14078_pp0_iter15_reg;
        p_read_1_reg_14078_pp0_iter17_reg <= p_read_1_reg_14078_pp0_iter16_reg;
        p_read_1_reg_14078_pp0_iter18_reg <= p_read_1_reg_14078_pp0_iter17_reg;
        p_read_1_reg_14078_pp0_iter19_reg <= p_read_1_reg_14078_pp0_iter18_reg;
        p_read_1_reg_14078_pp0_iter20_reg <= p_read_1_reg_14078_pp0_iter19_reg;
        p_read_1_reg_14078_pp0_iter21_reg <= p_read_1_reg_14078_pp0_iter20_reg;
        p_read_1_reg_14078_pp0_iter22_reg <= p_read_1_reg_14078_pp0_iter21_reg;
        p_read_1_reg_14078_pp0_iter2_reg <= p_read_1_reg_14078_pp0_iter1_reg;
        p_read_1_reg_14078_pp0_iter3_reg <= p_read_1_reg_14078_pp0_iter2_reg;
        p_read_1_reg_14078_pp0_iter4_reg <= p_read_1_reg_14078_pp0_iter3_reg;
        p_read_1_reg_14078_pp0_iter5_reg <= p_read_1_reg_14078_pp0_iter4_reg;
        p_read_1_reg_14078_pp0_iter6_reg <= p_read_1_reg_14078_pp0_iter5_reg;
        p_read_1_reg_14078_pp0_iter7_reg <= p_read_1_reg_14078_pp0_iter6_reg;
        p_read_1_reg_14078_pp0_iter8_reg <= p_read_1_reg_14078_pp0_iter7_reg;
        p_read_1_reg_14078_pp0_iter9_reg <= p_read_1_reg_14078_pp0_iter8_reg;
        p_read_2_reg_14083_pp0_iter10_reg <= p_read_2_reg_14083_pp0_iter9_reg;
        p_read_2_reg_14083_pp0_iter11_reg <= p_read_2_reg_14083_pp0_iter10_reg;
        p_read_2_reg_14083_pp0_iter12_reg <= p_read_2_reg_14083_pp0_iter11_reg;
        p_read_2_reg_14083_pp0_iter13_reg <= p_read_2_reg_14083_pp0_iter12_reg;
        p_read_2_reg_14083_pp0_iter14_reg <= p_read_2_reg_14083_pp0_iter13_reg;
        p_read_2_reg_14083_pp0_iter15_reg <= p_read_2_reg_14083_pp0_iter14_reg;
        p_read_2_reg_14083_pp0_iter16_reg <= p_read_2_reg_14083_pp0_iter15_reg;
        p_read_2_reg_14083_pp0_iter17_reg <= p_read_2_reg_14083_pp0_iter16_reg;
        p_read_2_reg_14083_pp0_iter18_reg <= p_read_2_reg_14083_pp0_iter17_reg;
        p_read_2_reg_14083_pp0_iter19_reg <= p_read_2_reg_14083_pp0_iter18_reg;
        p_read_2_reg_14083_pp0_iter20_reg <= p_read_2_reg_14083_pp0_iter19_reg;
        p_read_2_reg_14083_pp0_iter21_reg <= p_read_2_reg_14083_pp0_iter20_reg;
        p_read_2_reg_14083_pp0_iter2_reg <= p_read_2_reg_14083_pp0_iter1_reg;
        p_read_2_reg_14083_pp0_iter3_reg <= p_read_2_reg_14083_pp0_iter2_reg;
        p_read_2_reg_14083_pp0_iter4_reg <= p_read_2_reg_14083_pp0_iter3_reg;
        p_read_2_reg_14083_pp0_iter5_reg <= p_read_2_reg_14083_pp0_iter4_reg;
        p_read_2_reg_14083_pp0_iter6_reg <= p_read_2_reg_14083_pp0_iter5_reg;
        p_read_2_reg_14083_pp0_iter7_reg <= p_read_2_reg_14083_pp0_iter6_reg;
        p_read_2_reg_14083_pp0_iter8_reg <= p_read_2_reg_14083_pp0_iter7_reg;
        p_read_2_reg_14083_pp0_iter9_reg <= p_read_2_reg_14083_pp0_iter8_reg;
        p_read_3_reg_14088_pp0_iter10_reg <= p_read_3_reg_14088_pp0_iter9_reg;
        p_read_3_reg_14088_pp0_iter11_reg <= p_read_3_reg_14088_pp0_iter10_reg;
        p_read_3_reg_14088_pp0_iter12_reg <= p_read_3_reg_14088_pp0_iter11_reg;
        p_read_3_reg_14088_pp0_iter13_reg <= p_read_3_reg_14088_pp0_iter12_reg;
        p_read_3_reg_14088_pp0_iter14_reg <= p_read_3_reg_14088_pp0_iter13_reg;
        p_read_3_reg_14088_pp0_iter15_reg <= p_read_3_reg_14088_pp0_iter14_reg;
        p_read_3_reg_14088_pp0_iter16_reg <= p_read_3_reg_14088_pp0_iter15_reg;
        p_read_3_reg_14088_pp0_iter17_reg <= p_read_3_reg_14088_pp0_iter16_reg;
        p_read_3_reg_14088_pp0_iter18_reg <= p_read_3_reg_14088_pp0_iter17_reg;
        p_read_3_reg_14088_pp0_iter19_reg <= p_read_3_reg_14088_pp0_iter18_reg;
        p_read_3_reg_14088_pp0_iter2_reg <= p_read_3_reg_14088_pp0_iter1_reg;
        p_read_3_reg_14088_pp0_iter3_reg <= p_read_3_reg_14088_pp0_iter2_reg;
        p_read_3_reg_14088_pp0_iter4_reg <= p_read_3_reg_14088_pp0_iter3_reg;
        p_read_3_reg_14088_pp0_iter5_reg <= p_read_3_reg_14088_pp0_iter4_reg;
        p_read_3_reg_14088_pp0_iter6_reg <= p_read_3_reg_14088_pp0_iter5_reg;
        p_read_3_reg_14088_pp0_iter7_reg <= p_read_3_reg_14088_pp0_iter6_reg;
        p_read_3_reg_14088_pp0_iter8_reg <= p_read_3_reg_14088_pp0_iter7_reg;
        p_read_3_reg_14088_pp0_iter9_reg <= p_read_3_reg_14088_pp0_iter8_reg;
        p_read_4_reg_14093_pp0_iter10_reg <= p_read_4_reg_14093_pp0_iter9_reg;
        p_read_4_reg_14093_pp0_iter11_reg <= p_read_4_reg_14093_pp0_iter10_reg;
        p_read_4_reg_14093_pp0_iter12_reg <= p_read_4_reg_14093_pp0_iter11_reg;
        p_read_4_reg_14093_pp0_iter13_reg <= p_read_4_reg_14093_pp0_iter12_reg;
        p_read_4_reg_14093_pp0_iter14_reg <= p_read_4_reg_14093_pp0_iter13_reg;
        p_read_4_reg_14093_pp0_iter15_reg <= p_read_4_reg_14093_pp0_iter14_reg;
        p_read_4_reg_14093_pp0_iter16_reg <= p_read_4_reg_14093_pp0_iter15_reg;
        p_read_4_reg_14093_pp0_iter17_reg <= p_read_4_reg_14093_pp0_iter16_reg;
        p_read_4_reg_14093_pp0_iter2_reg <= p_read_4_reg_14093_pp0_iter1_reg;
        p_read_4_reg_14093_pp0_iter3_reg <= p_read_4_reg_14093_pp0_iter2_reg;
        p_read_4_reg_14093_pp0_iter4_reg <= p_read_4_reg_14093_pp0_iter3_reg;
        p_read_4_reg_14093_pp0_iter5_reg <= p_read_4_reg_14093_pp0_iter4_reg;
        p_read_4_reg_14093_pp0_iter6_reg <= p_read_4_reg_14093_pp0_iter5_reg;
        p_read_4_reg_14093_pp0_iter7_reg <= p_read_4_reg_14093_pp0_iter6_reg;
        p_read_4_reg_14093_pp0_iter8_reg <= p_read_4_reg_14093_pp0_iter7_reg;
        p_read_4_reg_14093_pp0_iter9_reg <= p_read_4_reg_14093_pp0_iter8_reg;
        p_read_5_reg_14098_pp0_iter10_reg <= p_read_5_reg_14098_pp0_iter9_reg;
        p_read_5_reg_14098_pp0_iter11_reg <= p_read_5_reg_14098_pp0_iter10_reg;
        p_read_5_reg_14098_pp0_iter12_reg <= p_read_5_reg_14098_pp0_iter11_reg;
        p_read_5_reg_14098_pp0_iter13_reg <= p_read_5_reg_14098_pp0_iter12_reg;
        p_read_5_reg_14098_pp0_iter14_reg <= p_read_5_reg_14098_pp0_iter13_reg;
        p_read_5_reg_14098_pp0_iter15_reg <= p_read_5_reg_14098_pp0_iter14_reg;
        p_read_5_reg_14098_pp0_iter2_reg <= p_read_5_reg_14098_pp0_iter1_reg;
        p_read_5_reg_14098_pp0_iter3_reg <= p_read_5_reg_14098_pp0_iter2_reg;
        p_read_5_reg_14098_pp0_iter4_reg <= p_read_5_reg_14098_pp0_iter3_reg;
        p_read_5_reg_14098_pp0_iter5_reg <= p_read_5_reg_14098_pp0_iter4_reg;
        p_read_5_reg_14098_pp0_iter6_reg <= p_read_5_reg_14098_pp0_iter5_reg;
        p_read_5_reg_14098_pp0_iter7_reg <= p_read_5_reg_14098_pp0_iter6_reg;
        p_read_5_reg_14098_pp0_iter8_reg <= p_read_5_reg_14098_pp0_iter7_reg;
        p_read_5_reg_14098_pp0_iter9_reg <= p_read_5_reg_14098_pp0_iter8_reg;
        p_read_6_reg_14103_pp0_iter10_reg <= p_read_6_reg_14103_pp0_iter9_reg;
        p_read_6_reg_14103_pp0_iter11_reg <= p_read_6_reg_14103_pp0_iter10_reg;
        p_read_6_reg_14103_pp0_iter12_reg <= p_read_6_reg_14103_pp0_iter11_reg;
        p_read_6_reg_14103_pp0_iter13_reg <= p_read_6_reg_14103_pp0_iter12_reg;
        p_read_6_reg_14103_pp0_iter2_reg <= p_read_6_reg_14103_pp0_iter1_reg;
        p_read_6_reg_14103_pp0_iter3_reg <= p_read_6_reg_14103_pp0_iter2_reg;
        p_read_6_reg_14103_pp0_iter4_reg <= p_read_6_reg_14103_pp0_iter3_reg;
        p_read_6_reg_14103_pp0_iter5_reg <= p_read_6_reg_14103_pp0_iter4_reg;
        p_read_6_reg_14103_pp0_iter6_reg <= p_read_6_reg_14103_pp0_iter5_reg;
        p_read_6_reg_14103_pp0_iter7_reg <= p_read_6_reg_14103_pp0_iter6_reg;
        p_read_6_reg_14103_pp0_iter8_reg <= p_read_6_reg_14103_pp0_iter7_reg;
        p_read_6_reg_14103_pp0_iter9_reg <= p_read_6_reg_14103_pp0_iter8_reg;
        p_read_7_reg_14108_pp0_iter10_reg <= p_read_7_reg_14108_pp0_iter9_reg;
        p_read_7_reg_14108_pp0_iter11_reg <= p_read_7_reg_14108_pp0_iter10_reg;
        p_read_7_reg_14108_pp0_iter2_reg <= p_read_7_reg_14108_pp0_iter1_reg;
        p_read_7_reg_14108_pp0_iter3_reg <= p_read_7_reg_14108_pp0_iter2_reg;
        p_read_7_reg_14108_pp0_iter4_reg <= p_read_7_reg_14108_pp0_iter3_reg;
        p_read_7_reg_14108_pp0_iter5_reg <= p_read_7_reg_14108_pp0_iter4_reg;
        p_read_7_reg_14108_pp0_iter6_reg <= p_read_7_reg_14108_pp0_iter5_reg;
        p_read_7_reg_14108_pp0_iter7_reg <= p_read_7_reg_14108_pp0_iter6_reg;
        p_read_7_reg_14108_pp0_iter8_reg <= p_read_7_reg_14108_pp0_iter7_reg;
        p_read_7_reg_14108_pp0_iter9_reg <= p_read_7_reg_14108_pp0_iter8_reg;
        p_read_8_reg_14113_pp0_iter2_reg <= p_read_8_reg_14113_pp0_iter1_reg;
        p_read_8_reg_14113_pp0_iter3_reg <= p_read_8_reg_14113_pp0_iter2_reg;
        p_read_8_reg_14113_pp0_iter4_reg <= p_read_8_reg_14113_pp0_iter3_reg;
        p_read_8_reg_14113_pp0_iter5_reg <= p_read_8_reg_14113_pp0_iter4_reg;
        p_read_8_reg_14113_pp0_iter6_reg <= p_read_8_reg_14113_pp0_iter5_reg;
        p_read_8_reg_14113_pp0_iter7_reg <= p_read_8_reg_14113_pp0_iter6_reg;
        p_read_8_reg_14113_pp0_iter8_reg <= p_read_8_reg_14113_pp0_iter7_reg;
        p_read_8_reg_14113_pp0_iter9_reg <= p_read_8_reg_14113_pp0_iter8_reg;
        p_read_9_reg_14118_pp0_iter2_reg <= p_read_9_reg_14118_pp0_iter1_reg;
        p_read_9_reg_14118_pp0_iter3_reg <= p_read_9_reg_14118_pp0_iter2_reg;
        p_read_9_reg_14118_pp0_iter4_reg <= p_read_9_reg_14118_pp0_iter3_reg;
        p_read_9_reg_14118_pp0_iter5_reg <= p_read_9_reg_14118_pp0_iter4_reg;
        p_read_9_reg_14118_pp0_iter6_reg <= p_read_9_reg_14118_pp0_iter5_reg;
        p_read_9_reg_14118_pp0_iter7_reg <= p_read_9_reg_14118_pp0_iter6_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        tmp_1_V_12_reg_14224 <= cipher_0_ssbox_q190;
        tmp_2_1_V_12_reg_14230 <= cipher_0_ssbox_q189;
        tmp_2_2_V_12_reg_14254 <= cipher_0_ssbox_q185;
        tmp_3_V_12_reg_14308 <= cipher_0_ssbox_q176;
        tmp_V_11_reg_14260 <= cipher_0_ssbox_q184;
        tmp_V_12_reg_14290 <= cipher_0_ssbox_q179;
        tmp_V_15_reg_14284 <= cipher_0_ssbox_q180;
        tmp_V_1_reg_14248 <= cipher_0_ssbox_q186;
        tmp_V_2_reg_14278 <= cipher_0_ssbox_q181;
        tmp_V_4_reg_14242 <= cipher_0_ssbox_q187;
        tmp_V_5_reg_14272 <= cipher_0_ssbox_q182;
        tmp_V_6_reg_14302 <= cipher_0_ssbox_q177;
        tmp_V_7_reg_14236 <= cipher_0_ssbox_q188;
        tmp_V_8_reg_14266 <= cipher_0_ssbox_q183;
        tmp_V_9_reg_14296 <= cipher_0_ssbox_q178;
        tmp_V_reg_14218 <= cipher_0_ssbox_q191;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        tmp_1_V_13_reg_14480 <= cipher_0_ssbox_q174;
        tmp_2_1_V_13_reg_14486 <= cipher_0_ssbox_q173;
        tmp_2_2_V_13_reg_14510 <= cipher_0_ssbox_q169;
        tmp_3_V_13_reg_14564 <= cipher_0_ssbox_q160;
        tmp_V_16_reg_14474 <= cipher_0_ssbox_q175;
        tmp_V_17_reg_14504 <= cipher_0_ssbox_q170;
        tmp_V_18_reg_14534 <= cipher_0_ssbox_q165;
        tmp_V_20_reg_14498 <= cipher_0_ssbox_q171;
        tmp_V_21_reg_14528 <= cipher_0_ssbox_q166;
        tmp_V_22_reg_14558 <= cipher_0_ssbox_q161;
        tmp_V_23_reg_14492 <= cipher_0_ssbox_q172;
        tmp_V_24_reg_14522 <= cipher_0_ssbox_q167;
        tmp_V_25_reg_14552 <= cipher_0_ssbox_q162;
        tmp_V_27_reg_14516 <= cipher_0_ssbox_q168;
        tmp_V_28_reg_14546 <= cipher_0_ssbox_q163;
        tmp_V_31_reg_14540 <= cipher_0_ssbox_q164;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        tmp_1_V_14_reg_14736 <= cipher_0_ssbox_q158;
        tmp_2_1_V_14_reg_14742 <= cipher_0_ssbox_q157;
        tmp_2_2_V_14_reg_14766 <= cipher_0_ssbox_q153;
        tmp_3_V_14_reg_14820 <= cipher_0_ssbox_q144;
        tmp_V_32_reg_14730 <= cipher_0_ssbox_q159;
        tmp_V_33_reg_14760 <= cipher_0_ssbox_q154;
        tmp_V_34_reg_14790 <= cipher_0_ssbox_q149;
        tmp_V_36_reg_14754 <= cipher_0_ssbox_q155;
        tmp_V_37_reg_14784 <= cipher_0_ssbox_q150;
        tmp_V_38_reg_14814 <= cipher_0_ssbox_q145;
        tmp_V_39_reg_14748 <= cipher_0_ssbox_q156;
        tmp_V_40_reg_14778 <= cipher_0_ssbox_q151;
        tmp_V_41_reg_14808 <= cipher_0_ssbox_q146;
        tmp_V_43_reg_14772 <= cipher_0_ssbox_q152;
        tmp_V_44_reg_14802 <= cipher_0_ssbox_q147;
        tmp_V_47_reg_14796 <= cipher_0_ssbox_q148;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        tmp_1_V_15_reg_14992 <= cipher_0_ssbox_q142;
        tmp_2_1_V_15_reg_14998 <= cipher_0_ssbox_q141;
        tmp_2_2_V_15_reg_15022 <= cipher_0_ssbox_q137;
        tmp_3_V_15_reg_15076 <= cipher_0_ssbox_q128;
        tmp_V_48_reg_14986 <= cipher_0_ssbox_q143;
        tmp_V_49_reg_15016 <= cipher_0_ssbox_q138;
        tmp_V_50_reg_15046 <= cipher_0_ssbox_q133;
        tmp_V_52_reg_15010 <= cipher_0_ssbox_q139;
        tmp_V_53_reg_15040 <= cipher_0_ssbox_q134;
        tmp_V_54_reg_15070 <= cipher_0_ssbox_q129;
        tmp_V_55_reg_15004 <= cipher_0_ssbox_q140;
        tmp_V_56_reg_15034 <= cipher_0_ssbox_q135;
        tmp_V_57_reg_15064 <= cipher_0_ssbox_q130;
        tmp_V_59_reg_15028 <= cipher_0_ssbox_q136;
        tmp_V_60_reg_15058 <= cipher_0_ssbox_q131;
        tmp_V_63_reg_15052 <= cipher_0_ssbox_q132;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        tmp_1_V_16_reg_15248 <= cipher_0_ssbox_q126;
        tmp_2_1_V_16_reg_15254 <= cipher_0_ssbox_q125;
        tmp_2_2_V_16_reg_15278 <= cipher_0_ssbox_q121;
        tmp_3_V_16_reg_15332 <= cipher_0_ssbox_q112;
        tmp_V_64_reg_15242 <= cipher_0_ssbox_q127;
        tmp_V_65_reg_15272 <= cipher_0_ssbox_q122;
        tmp_V_66_reg_15302 <= cipher_0_ssbox_q117;
        tmp_V_68_reg_15266 <= cipher_0_ssbox_q123;
        tmp_V_69_reg_15296 <= cipher_0_ssbox_q118;
        tmp_V_70_reg_15326 <= cipher_0_ssbox_q113;
        tmp_V_71_reg_15260 <= cipher_0_ssbox_q124;
        tmp_V_72_reg_15290 <= cipher_0_ssbox_q119;
        tmp_V_73_reg_15320 <= cipher_0_ssbox_q114;
        tmp_V_75_reg_15284 <= cipher_0_ssbox_q120;
        tmp_V_76_reg_15314 <= cipher_0_ssbox_q115;
        tmp_V_79_reg_15308 <= cipher_0_ssbox_q116;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        tmp_1_V_17_reg_15504 <= cipher_0_ssbox_q110;
        tmp_2_1_V_17_reg_15510 <= cipher_0_ssbox_q109;
        tmp_2_2_V_17_reg_15534 <= cipher_0_ssbox_q105;
        tmp_3_V_17_reg_15588 <= cipher_0_ssbox_q96;
        tmp_V_80_reg_15498 <= cipher_0_ssbox_q111;
        tmp_V_81_reg_15528 <= cipher_0_ssbox_q106;
        tmp_V_82_reg_15558 <= cipher_0_ssbox_q101;
        tmp_V_84_reg_15522 <= cipher_0_ssbox_q107;
        tmp_V_85_reg_15552 <= cipher_0_ssbox_q102;
        tmp_V_86_reg_15582 <= cipher_0_ssbox_q97;
        tmp_V_87_reg_15516 <= cipher_0_ssbox_q108;
        tmp_V_88_reg_15546 <= cipher_0_ssbox_q103;
        tmp_V_89_reg_15576 <= cipher_0_ssbox_q98;
        tmp_V_91_reg_15540 <= cipher_0_ssbox_q104;
        tmp_V_92_reg_15570 <= cipher_0_ssbox_q99;
        tmp_V_95_reg_15564 <= cipher_0_ssbox_q100;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        tmp_1_V_18_reg_15760 <= cipher_0_ssbox_q94;
        tmp_2_1_V_18_reg_15766 <= cipher_0_ssbox_q93;
        tmp_2_2_V_18_reg_15790 <= cipher_0_ssbox_q89;
        tmp_3_V_18_reg_15844 <= cipher_0_ssbox_q80;
        tmp_V_100_reg_15778 <= cipher_0_ssbox_q91;
        tmp_V_101_reg_15808 <= cipher_0_ssbox_q86;
        tmp_V_102_reg_15838 <= cipher_0_ssbox_q81;
        tmp_V_103_reg_15772 <= cipher_0_ssbox_q92;
        tmp_V_104_reg_15802 <= cipher_0_ssbox_q87;
        tmp_V_105_reg_15832 <= cipher_0_ssbox_q82;
        tmp_V_107_reg_15796 <= cipher_0_ssbox_q88;
        tmp_V_108_reg_15826 <= cipher_0_ssbox_q83;
        tmp_V_111_reg_15820 <= cipher_0_ssbox_q84;
        tmp_V_96_reg_15754 <= cipher_0_ssbox_q95;
        tmp_V_97_reg_15784 <= cipher_0_ssbox_q90;
        tmp_V_98_reg_15814 <= cipher_0_ssbox_q85;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        tmp_1_V_19_reg_16016 <= cipher_0_ssbox_q78;
        tmp_2_1_V_19_reg_16022 <= cipher_0_ssbox_q77;
        tmp_2_2_V_19_reg_16046 <= cipher_0_ssbox_q73;
        tmp_3_V_19_reg_16100 <= cipher_0_ssbox_q64;
        tmp_V_112_reg_16010 <= cipher_0_ssbox_q79;
        tmp_V_113_reg_16040 <= cipher_0_ssbox_q74;
        tmp_V_114_reg_16070 <= cipher_0_ssbox_q69;
        tmp_V_116_reg_16034 <= cipher_0_ssbox_q75;
        tmp_V_117_reg_16064 <= cipher_0_ssbox_q70;
        tmp_V_118_reg_16094 <= cipher_0_ssbox_q65;
        tmp_V_119_reg_16028 <= cipher_0_ssbox_q76;
        tmp_V_120_reg_16058 <= cipher_0_ssbox_q71;
        tmp_V_121_reg_16088 <= cipher_0_ssbox_q66;
        tmp_V_123_reg_16052 <= cipher_0_ssbox_q72;
        tmp_V_124_reg_16082 <= cipher_0_ssbox_q67;
        tmp_V_127_reg_16076 <= cipher_0_ssbox_q68;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        tmp_1_V_20_reg_16272 <= cipher_0_ssbox_q62;
        tmp_2_1_V_20_reg_16278 <= cipher_0_ssbox_q61;
        tmp_2_2_V_20_reg_16302 <= cipher_0_ssbox_q57;
        tmp_3_V_20_reg_16356 <= cipher_0_ssbox_q48;
        tmp_V_128_reg_16266 <= cipher_0_ssbox_q63;
        tmp_V_129_reg_16296 <= cipher_0_ssbox_q58;
        tmp_V_130_reg_16326 <= cipher_0_ssbox_q53;
        tmp_V_132_reg_16290 <= cipher_0_ssbox_q59;
        tmp_V_133_reg_16320 <= cipher_0_ssbox_q54;
        tmp_V_134_reg_16350 <= cipher_0_ssbox_q49;
        tmp_V_135_reg_16284 <= cipher_0_ssbox_q60;
        tmp_V_136_reg_16314 <= cipher_0_ssbox_q55;
        tmp_V_137_reg_16344 <= cipher_0_ssbox_q50;
        tmp_V_139_reg_16308 <= cipher_0_ssbox_q56;
        tmp_V_140_reg_16338 <= cipher_0_ssbox_q51;
        tmp_V_143_reg_16332 <= cipher_0_ssbox_q52;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        tmp_1_V_21_reg_16528 <= cipher_0_ssbox_q46;
        tmp_2_1_V_21_reg_16534 <= cipher_0_ssbox_q45;
        tmp_2_2_V_21_reg_16558 <= cipher_0_ssbox_q41;
        tmp_3_V_21_reg_16612 <= cipher_0_ssbox_q32;
        tmp_V_144_reg_16522 <= cipher_0_ssbox_q47;
        tmp_V_145_reg_16552 <= cipher_0_ssbox_q42;
        tmp_V_146_reg_16582 <= cipher_0_ssbox_q37;
        tmp_V_148_reg_16546 <= cipher_0_ssbox_q43;
        tmp_V_149_reg_16576 <= cipher_0_ssbox_q38;
        tmp_V_150_reg_16606 <= cipher_0_ssbox_q33;
        tmp_V_151_reg_16540 <= cipher_0_ssbox_q44;
        tmp_V_152_reg_16570 <= cipher_0_ssbox_q39;
        tmp_V_153_reg_16600 <= cipher_0_ssbox_q34;
        tmp_V_155_reg_16564 <= cipher_0_ssbox_q40;
        tmp_V_156_reg_16594 <= cipher_0_ssbox_q35;
        tmp_V_159_reg_16588 <= cipher_0_ssbox_q36;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        tmp_1_V_22_reg_16784 <= cipher_0_ssbox_q30;
        tmp_2_1_V_22_reg_16790 <= cipher_0_ssbox_q29;
        tmp_2_2_V_22_reg_16814 <= cipher_0_ssbox_q25;
        tmp_3_V_22_reg_16868 <= cipher_0_ssbox_q16;
        tmp_V_160_reg_16778 <= cipher_0_ssbox_q31;
        tmp_V_161_reg_16808 <= cipher_0_ssbox_q26;
        tmp_V_162_reg_16838 <= cipher_0_ssbox_q21;
        tmp_V_164_reg_16802 <= cipher_0_ssbox_q27;
        tmp_V_165_reg_16832 <= cipher_0_ssbox_q22;
        tmp_V_166_reg_16862 <= cipher_0_ssbox_q17;
        tmp_V_167_reg_16796 <= cipher_0_ssbox_q28;
        tmp_V_168_reg_16826 <= cipher_0_ssbox_q23;
        tmp_V_169_reg_16856 <= cipher_0_ssbox_q18;
        tmp_V_171_reg_16820 <= cipher_0_ssbox_q24;
        tmp_V_172_reg_16850 <= cipher_0_ssbox_q19;
        tmp_V_175_reg_16844 <= cipher_0_ssbox_q20;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter23 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_idle_pp0 == 1'b1) & (ap_start == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter23 == 1'b0) & (ap_enable_reg_pp0_iter22 == 1'b0) & (ap_enable_reg_pp0_iter21 == 1'b0) & (ap_enable_reg_pp0_iter20 == 1'b0) & (ap_enable_reg_pp0_iter19 == 1'b0) & (ap_enable_reg_pp0_iter18 == 1'b0) & (ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b0) & (ap_enable_reg_pp0_iter21 == 1'b0) & (ap_enable_reg_pp0_iter20 == 1'b0) & (ap_enable_reg_pp0_iter19 == 1'b0) & (ap_enable_reg_pp0_iter18 == 1'b0) & (ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0_0to22 = 1'b1;
    end else begin
        ap_idle_pp0_0to22 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((ap_idle_pp0_0to22 == 1'b1) & (ap_start == 1'b0))) begin
        ap_reset_idle_pp0 = 1'b1;
    end else begin
        ap_reset_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce0 = 1'b1;
    end else begin
        cipher_0_p16box_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce1 = 1'b1;
    end else begin
        cipher_0_p16box_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce10 = 1'b1;
    end else begin
        cipher_0_p16box_ce10 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce100 = 1'b1;
    end else begin
        cipher_0_p16box_ce100 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce101 = 1'b1;
    end else begin
        cipher_0_p16box_ce101 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce102 = 1'b1;
    end else begin
        cipher_0_p16box_ce102 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce103 = 1'b1;
    end else begin
        cipher_0_p16box_ce103 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce104 = 1'b1;
    end else begin
        cipher_0_p16box_ce104 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce105 = 1'b1;
    end else begin
        cipher_0_p16box_ce105 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce106 = 1'b1;
    end else begin
        cipher_0_p16box_ce106 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce107 = 1'b1;
    end else begin
        cipher_0_p16box_ce107 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce108 = 1'b1;
    end else begin
        cipher_0_p16box_ce108 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce109 = 1'b1;
    end else begin
        cipher_0_p16box_ce109 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce11 = 1'b1;
    end else begin
        cipher_0_p16box_ce11 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce110 = 1'b1;
    end else begin
        cipher_0_p16box_ce110 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce111 = 1'b1;
    end else begin
        cipher_0_p16box_ce111 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce112 = 1'b1;
    end else begin
        cipher_0_p16box_ce112 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce113 = 1'b1;
    end else begin
        cipher_0_p16box_ce113 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce114 = 1'b1;
    end else begin
        cipher_0_p16box_ce114 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce115 = 1'b1;
    end else begin
        cipher_0_p16box_ce115 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce116 = 1'b1;
    end else begin
        cipher_0_p16box_ce116 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce117 = 1'b1;
    end else begin
        cipher_0_p16box_ce117 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce118 = 1'b1;
    end else begin
        cipher_0_p16box_ce118 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce119 = 1'b1;
    end else begin
        cipher_0_p16box_ce119 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce12 = 1'b1;
    end else begin
        cipher_0_p16box_ce12 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce120 = 1'b1;
    end else begin
        cipher_0_p16box_ce120 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce121 = 1'b1;
    end else begin
        cipher_0_p16box_ce121 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce122 = 1'b1;
    end else begin
        cipher_0_p16box_ce122 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce123 = 1'b1;
    end else begin
        cipher_0_p16box_ce123 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce124 = 1'b1;
    end else begin
        cipher_0_p16box_ce124 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce125 = 1'b1;
    end else begin
        cipher_0_p16box_ce125 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce126 = 1'b1;
    end else begin
        cipher_0_p16box_ce126 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce127 = 1'b1;
    end else begin
        cipher_0_p16box_ce127 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce128 = 1'b1;
    end else begin
        cipher_0_p16box_ce128 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce129 = 1'b1;
    end else begin
        cipher_0_p16box_ce129 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce13 = 1'b1;
    end else begin
        cipher_0_p16box_ce13 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce130 = 1'b1;
    end else begin
        cipher_0_p16box_ce130 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce131 = 1'b1;
    end else begin
        cipher_0_p16box_ce131 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce132 = 1'b1;
    end else begin
        cipher_0_p16box_ce132 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce133 = 1'b1;
    end else begin
        cipher_0_p16box_ce133 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce134 = 1'b1;
    end else begin
        cipher_0_p16box_ce134 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce135 = 1'b1;
    end else begin
        cipher_0_p16box_ce135 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce136 = 1'b1;
    end else begin
        cipher_0_p16box_ce136 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce137 = 1'b1;
    end else begin
        cipher_0_p16box_ce137 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce138 = 1'b1;
    end else begin
        cipher_0_p16box_ce138 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce139 = 1'b1;
    end else begin
        cipher_0_p16box_ce139 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce14 = 1'b1;
    end else begin
        cipher_0_p16box_ce14 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce140 = 1'b1;
    end else begin
        cipher_0_p16box_ce140 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce141 = 1'b1;
    end else begin
        cipher_0_p16box_ce141 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce142 = 1'b1;
    end else begin
        cipher_0_p16box_ce142 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce143 = 1'b1;
    end else begin
        cipher_0_p16box_ce143 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce144 = 1'b1;
    end else begin
        cipher_0_p16box_ce144 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce145 = 1'b1;
    end else begin
        cipher_0_p16box_ce145 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce146 = 1'b1;
    end else begin
        cipher_0_p16box_ce146 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce147 = 1'b1;
    end else begin
        cipher_0_p16box_ce147 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce148 = 1'b1;
    end else begin
        cipher_0_p16box_ce148 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce149 = 1'b1;
    end else begin
        cipher_0_p16box_ce149 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce15 = 1'b1;
    end else begin
        cipher_0_p16box_ce15 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce150 = 1'b1;
    end else begin
        cipher_0_p16box_ce150 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce151 = 1'b1;
    end else begin
        cipher_0_p16box_ce151 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce152 = 1'b1;
    end else begin
        cipher_0_p16box_ce152 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce153 = 1'b1;
    end else begin
        cipher_0_p16box_ce153 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce154 = 1'b1;
    end else begin
        cipher_0_p16box_ce154 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce155 = 1'b1;
    end else begin
        cipher_0_p16box_ce155 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce156 = 1'b1;
    end else begin
        cipher_0_p16box_ce156 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce157 = 1'b1;
    end else begin
        cipher_0_p16box_ce157 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce158 = 1'b1;
    end else begin
        cipher_0_p16box_ce158 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce159 = 1'b1;
    end else begin
        cipher_0_p16box_ce159 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce16 = 1'b1;
    end else begin
        cipher_0_p16box_ce16 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce160 = 1'b1;
    end else begin
        cipher_0_p16box_ce160 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce161 = 1'b1;
    end else begin
        cipher_0_p16box_ce161 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce162 = 1'b1;
    end else begin
        cipher_0_p16box_ce162 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce163 = 1'b1;
    end else begin
        cipher_0_p16box_ce163 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce164 = 1'b1;
    end else begin
        cipher_0_p16box_ce164 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce165 = 1'b1;
    end else begin
        cipher_0_p16box_ce165 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce166 = 1'b1;
    end else begin
        cipher_0_p16box_ce166 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce167 = 1'b1;
    end else begin
        cipher_0_p16box_ce167 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce168 = 1'b1;
    end else begin
        cipher_0_p16box_ce168 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce169 = 1'b1;
    end else begin
        cipher_0_p16box_ce169 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce17 = 1'b1;
    end else begin
        cipher_0_p16box_ce17 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce170 = 1'b1;
    end else begin
        cipher_0_p16box_ce170 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce171 = 1'b1;
    end else begin
        cipher_0_p16box_ce171 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce172 = 1'b1;
    end else begin
        cipher_0_p16box_ce172 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce173 = 1'b1;
    end else begin
        cipher_0_p16box_ce173 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce174 = 1'b1;
    end else begin
        cipher_0_p16box_ce174 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce175 = 1'b1;
    end else begin
        cipher_0_p16box_ce175 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce18 = 1'b1;
    end else begin
        cipher_0_p16box_ce18 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce19 = 1'b1;
    end else begin
        cipher_0_p16box_ce19 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce2 = 1'b1;
    end else begin
        cipher_0_p16box_ce2 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce20 = 1'b1;
    end else begin
        cipher_0_p16box_ce20 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce21 = 1'b1;
    end else begin
        cipher_0_p16box_ce21 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce22 = 1'b1;
    end else begin
        cipher_0_p16box_ce22 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce23 = 1'b1;
    end else begin
        cipher_0_p16box_ce23 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce24 = 1'b1;
    end else begin
        cipher_0_p16box_ce24 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce25 = 1'b1;
    end else begin
        cipher_0_p16box_ce25 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce26 = 1'b1;
    end else begin
        cipher_0_p16box_ce26 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce27 = 1'b1;
    end else begin
        cipher_0_p16box_ce27 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce28 = 1'b1;
    end else begin
        cipher_0_p16box_ce28 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce29 = 1'b1;
    end else begin
        cipher_0_p16box_ce29 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce3 = 1'b1;
    end else begin
        cipher_0_p16box_ce3 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce30 = 1'b1;
    end else begin
        cipher_0_p16box_ce30 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce31 = 1'b1;
    end else begin
        cipher_0_p16box_ce31 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce32 = 1'b1;
    end else begin
        cipher_0_p16box_ce32 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce33 = 1'b1;
    end else begin
        cipher_0_p16box_ce33 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce34 = 1'b1;
    end else begin
        cipher_0_p16box_ce34 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce35 = 1'b1;
    end else begin
        cipher_0_p16box_ce35 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce36 = 1'b1;
    end else begin
        cipher_0_p16box_ce36 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce37 = 1'b1;
    end else begin
        cipher_0_p16box_ce37 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce38 = 1'b1;
    end else begin
        cipher_0_p16box_ce38 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce39 = 1'b1;
    end else begin
        cipher_0_p16box_ce39 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce4 = 1'b1;
    end else begin
        cipher_0_p16box_ce4 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce40 = 1'b1;
    end else begin
        cipher_0_p16box_ce40 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce41 = 1'b1;
    end else begin
        cipher_0_p16box_ce41 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce42 = 1'b1;
    end else begin
        cipher_0_p16box_ce42 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce43 = 1'b1;
    end else begin
        cipher_0_p16box_ce43 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce44 = 1'b1;
    end else begin
        cipher_0_p16box_ce44 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce45 = 1'b1;
    end else begin
        cipher_0_p16box_ce45 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce46 = 1'b1;
    end else begin
        cipher_0_p16box_ce46 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce47 = 1'b1;
    end else begin
        cipher_0_p16box_ce47 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce48 = 1'b1;
    end else begin
        cipher_0_p16box_ce48 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce49 = 1'b1;
    end else begin
        cipher_0_p16box_ce49 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce5 = 1'b1;
    end else begin
        cipher_0_p16box_ce5 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce50 = 1'b1;
    end else begin
        cipher_0_p16box_ce50 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce51 = 1'b1;
    end else begin
        cipher_0_p16box_ce51 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce52 = 1'b1;
    end else begin
        cipher_0_p16box_ce52 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce53 = 1'b1;
    end else begin
        cipher_0_p16box_ce53 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce54 = 1'b1;
    end else begin
        cipher_0_p16box_ce54 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce55 = 1'b1;
    end else begin
        cipher_0_p16box_ce55 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce56 = 1'b1;
    end else begin
        cipher_0_p16box_ce56 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce57 = 1'b1;
    end else begin
        cipher_0_p16box_ce57 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce58 = 1'b1;
    end else begin
        cipher_0_p16box_ce58 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce59 = 1'b1;
    end else begin
        cipher_0_p16box_ce59 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce6 = 1'b1;
    end else begin
        cipher_0_p16box_ce6 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce60 = 1'b1;
    end else begin
        cipher_0_p16box_ce60 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce61 = 1'b1;
    end else begin
        cipher_0_p16box_ce61 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce62 = 1'b1;
    end else begin
        cipher_0_p16box_ce62 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce63 = 1'b1;
    end else begin
        cipher_0_p16box_ce63 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce64 = 1'b1;
    end else begin
        cipher_0_p16box_ce64 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce65 = 1'b1;
    end else begin
        cipher_0_p16box_ce65 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce66 = 1'b1;
    end else begin
        cipher_0_p16box_ce66 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce67 = 1'b1;
    end else begin
        cipher_0_p16box_ce67 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce68 = 1'b1;
    end else begin
        cipher_0_p16box_ce68 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce69 = 1'b1;
    end else begin
        cipher_0_p16box_ce69 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce7 = 1'b1;
    end else begin
        cipher_0_p16box_ce7 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce70 = 1'b1;
    end else begin
        cipher_0_p16box_ce70 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce71 = 1'b1;
    end else begin
        cipher_0_p16box_ce71 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce72 = 1'b1;
    end else begin
        cipher_0_p16box_ce72 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce73 = 1'b1;
    end else begin
        cipher_0_p16box_ce73 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce74 = 1'b1;
    end else begin
        cipher_0_p16box_ce74 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce75 = 1'b1;
    end else begin
        cipher_0_p16box_ce75 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce76 = 1'b1;
    end else begin
        cipher_0_p16box_ce76 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce77 = 1'b1;
    end else begin
        cipher_0_p16box_ce77 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce78 = 1'b1;
    end else begin
        cipher_0_p16box_ce78 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce79 = 1'b1;
    end else begin
        cipher_0_p16box_ce79 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce8 = 1'b1;
    end else begin
        cipher_0_p16box_ce8 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce80 = 1'b1;
    end else begin
        cipher_0_p16box_ce80 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce81 = 1'b1;
    end else begin
        cipher_0_p16box_ce81 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce82 = 1'b1;
    end else begin
        cipher_0_p16box_ce82 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce83 = 1'b1;
    end else begin
        cipher_0_p16box_ce83 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce84 = 1'b1;
    end else begin
        cipher_0_p16box_ce84 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce85 = 1'b1;
    end else begin
        cipher_0_p16box_ce85 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce86 = 1'b1;
    end else begin
        cipher_0_p16box_ce86 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce87 = 1'b1;
    end else begin
        cipher_0_p16box_ce87 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce88 = 1'b1;
    end else begin
        cipher_0_p16box_ce88 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce89 = 1'b1;
    end else begin
        cipher_0_p16box_ce89 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce9 = 1'b1;
    end else begin
        cipher_0_p16box_ce9 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce90 = 1'b1;
    end else begin
        cipher_0_p16box_ce90 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce91 = 1'b1;
    end else begin
        cipher_0_p16box_ce91 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce92 = 1'b1;
    end else begin
        cipher_0_p16box_ce92 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce93 = 1'b1;
    end else begin
        cipher_0_p16box_ce93 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce94 = 1'b1;
    end else begin
        cipher_0_p16box_ce94 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce95 = 1'b1;
    end else begin
        cipher_0_p16box_ce95 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce96 = 1'b1;
    end else begin
        cipher_0_p16box_ce96 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce97 = 1'b1;
    end else begin
        cipher_0_p16box_ce97 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce98 = 1'b1;
    end else begin
        cipher_0_p16box_ce98 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce99 = 1'b1;
    end else begin
        cipher_0_p16box_ce99 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce0 = 1'b1;
    end else begin
        cipher_0_ssbox_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce1 = 1'b1;
    end else begin
        cipher_0_ssbox_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce10 = 1'b1;
    end else begin
        cipher_0_ssbox_ce10 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce100 = 1'b1;
    end else begin
        cipher_0_ssbox_ce100 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce101 = 1'b1;
    end else begin
        cipher_0_ssbox_ce101 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce102 = 1'b1;
    end else begin
        cipher_0_ssbox_ce102 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce103 = 1'b1;
    end else begin
        cipher_0_ssbox_ce103 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce104 = 1'b1;
    end else begin
        cipher_0_ssbox_ce104 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce105 = 1'b1;
    end else begin
        cipher_0_ssbox_ce105 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce106 = 1'b1;
    end else begin
        cipher_0_ssbox_ce106 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce107 = 1'b1;
    end else begin
        cipher_0_ssbox_ce107 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce108 = 1'b1;
    end else begin
        cipher_0_ssbox_ce108 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce109 = 1'b1;
    end else begin
        cipher_0_ssbox_ce109 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce11 = 1'b1;
    end else begin
        cipher_0_ssbox_ce11 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce110 = 1'b1;
    end else begin
        cipher_0_ssbox_ce110 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce111 = 1'b1;
    end else begin
        cipher_0_ssbox_ce111 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce112 = 1'b1;
    end else begin
        cipher_0_ssbox_ce112 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce113 = 1'b1;
    end else begin
        cipher_0_ssbox_ce113 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce114 = 1'b1;
    end else begin
        cipher_0_ssbox_ce114 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce115 = 1'b1;
    end else begin
        cipher_0_ssbox_ce115 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce116 = 1'b1;
    end else begin
        cipher_0_ssbox_ce116 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce117 = 1'b1;
    end else begin
        cipher_0_ssbox_ce117 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce118 = 1'b1;
    end else begin
        cipher_0_ssbox_ce118 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce119 = 1'b1;
    end else begin
        cipher_0_ssbox_ce119 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce12 = 1'b1;
    end else begin
        cipher_0_ssbox_ce12 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce120 = 1'b1;
    end else begin
        cipher_0_ssbox_ce120 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce121 = 1'b1;
    end else begin
        cipher_0_ssbox_ce121 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce122 = 1'b1;
    end else begin
        cipher_0_ssbox_ce122 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce123 = 1'b1;
    end else begin
        cipher_0_ssbox_ce123 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce124 = 1'b1;
    end else begin
        cipher_0_ssbox_ce124 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce125 = 1'b1;
    end else begin
        cipher_0_ssbox_ce125 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce126 = 1'b1;
    end else begin
        cipher_0_ssbox_ce126 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce127 = 1'b1;
    end else begin
        cipher_0_ssbox_ce127 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce128 = 1'b1;
    end else begin
        cipher_0_ssbox_ce128 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce129 = 1'b1;
    end else begin
        cipher_0_ssbox_ce129 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce13 = 1'b1;
    end else begin
        cipher_0_ssbox_ce13 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce130 = 1'b1;
    end else begin
        cipher_0_ssbox_ce130 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce131 = 1'b1;
    end else begin
        cipher_0_ssbox_ce131 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce132 = 1'b1;
    end else begin
        cipher_0_ssbox_ce132 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce133 = 1'b1;
    end else begin
        cipher_0_ssbox_ce133 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce134 = 1'b1;
    end else begin
        cipher_0_ssbox_ce134 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce135 = 1'b1;
    end else begin
        cipher_0_ssbox_ce135 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce136 = 1'b1;
    end else begin
        cipher_0_ssbox_ce136 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce137 = 1'b1;
    end else begin
        cipher_0_ssbox_ce137 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce138 = 1'b1;
    end else begin
        cipher_0_ssbox_ce138 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce139 = 1'b1;
    end else begin
        cipher_0_ssbox_ce139 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce14 = 1'b1;
    end else begin
        cipher_0_ssbox_ce14 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce140 = 1'b1;
    end else begin
        cipher_0_ssbox_ce140 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce141 = 1'b1;
    end else begin
        cipher_0_ssbox_ce141 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce142 = 1'b1;
    end else begin
        cipher_0_ssbox_ce142 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce143 = 1'b1;
    end else begin
        cipher_0_ssbox_ce143 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce144 = 1'b1;
    end else begin
        cipher_0_ssbox_ce144 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce145 = 1'b1;
    end else begin
        cipher_0_ssbox_ce145 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce146 = 1'b1;
    end else begin
        cipher_0_ssbox_ce146 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce147 = 1'b1;
    end else begin
        cipher_0_ssbox_ce147 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce148 = 1'b1;
    end else begin
        cipher_0_ssbox_ce148 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce149 = 1'b1;
    end else begin
        cipher_0_ssbox_ce149 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce15 = 1'b1;
    end else begin
        cipher_0_ssbox_ce15 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce150 = 1'b1;
    end else begin
        cipher_0_ssbox_ce150 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce151 = 1'b1;
    end else begin
        cipher_0_ssbox_ce151 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce152 = 1'b1;
    end else begin
        cipher_0_ssbox_ce152 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce153 = 1'b1;
    end else begin
        cipher_0_ssbox_ce153 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce154 = 1'b1;
    end else begin
        cipher_0_ssbox_ce154 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce155 = 1'b1;
    end else begin
        cipher_0_ssbox_ce155 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce156 = 1'b1;
    end else begin
        cipher_0_ssbox_ce156 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce157 = 1'b1;
    end else begin
        cipher_0_ssbox_ce157 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce158 = 1'b1;
    end else begin
        cipher_0_ssbox_ce158 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce159 = 1'b1;
    end else begin
        cipher_0_ssbox_ce159 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce16 = 1'b1;
    end else begin
        cipher_0_ssbox_ce16 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce160 = 1'b1;
    end else begin
        cipher_0_ssbox_ce160 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce161 = 1'b1;
    end else begin
        cipher_0_ssbox_ce161 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce162 = 1'b1;
    end else begin
        cipher_0_ssbox_ce162 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce163 = 1'b1;
    end else begin
        cipher_0_ssbox_ce163 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce164 = 1'b1;
    end else begin
        cipher_0_ssbox_ce164 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce165 = 1'b1;
    end else begin
        cipher_0_ssbox_ce165 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce166 = 1'b1;
    end else begin
        cipher_0_ssbox_ce166 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce167 = 1'b1;
    end else begin
        cipher_0_ssbox_ce167 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce168 = 1'b1;
    end else begin
        cipher_0_ssbox_ce168 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce169 = 1'b1;
    end else begin
        cipher_0_ssbox_ce169 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce17 = 1'b1;
    end else begin
        cipher_0_ssbox_ce17 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce170 = 1'b1;
    end else begin
        cipher_0_ssbox_ce170 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce171 = 1'b1;
    end else begin
        cipher_0_ssbox_ce171 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce172 = 1'b1;
    end else begin
        cipher_0_ssbox_ce172 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce173 = 1'b1;
    end else begin
        cipher_0_ssbox_ce173 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce174 = 1'b1;
    end else begin
        cipher_0_ssbox_ce174 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce175 = 1'b1;
    end else begin
        cipher_0_ssbox_ce175 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce176 = 1'b1;
    end else begin
        cipher_0_ssbox_ce176 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce177 = 1'b1;
    end else begin
        cipher_0_ssbox_ce177 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce178 = 1'b1;
    end else begin
        cipher_0_ssbox_ce178 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce179 = 1'b1;
    end else begin
        cipher_0_ssbox_ce179 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce18 = 1'b1;
    end else begin
        cipher_0_ssbox_ce18 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce180 = 1'b1;
    end else begin
        cipher_0_ssbox_ce180 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce181 = 1'b1;
    end else begin
        cipher_0_ssbox_ce181 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce182 = 1'b1;
    end else begin
        cipher_0_ssbox_ce182 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce183 = 1'b1;
    end else begin
        cipher_0_ssbox_ce183 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce184 = 1'b1;
    end else begin
        cipher_0_ssbox_ce184 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce185 = 1'b1;
    end else begin
        cipher_0_ssbox_ce185 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce186 = 1'b1;
    end else begin
        cipher_0_ssbox_ce186 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce187 = 1'b1;
    end else begin
        cipher_0_ssbox_ce187 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce188 = 1'b1;
    end else begin
        cipher_0_ssbox_ce188 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce189 = 1'b1;
    end else begin
        cipher_0_ssbox_ce189 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce19 = 1'b1;
    end else begin
        cipher_0_ssbox_ce19 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce190 = 1'b1;
    end else begin
        cipher_0_ssbox_ce190 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce191 = 1'b1;
    end else begin
        cipher_0_ssbox_ce191 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce2 = 1'b1;
    end else begin
        cipher_0_ssbox_ce2 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce20 = 1'b1;
    end else begin
        cipher_0_ssbox_ce20 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce21 = 1'b1;
    end else begin
        cipher_0_ssbox_ce21 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce22 = 1'b1;
    end else begin
        cipher_0_ssbox_ce22 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce23 = 1'b1;
    end else begin
        cipher_0_ssbox_ce23 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce24 = 1'b1;
    end else begin
        cipher_0_ssbox_ce24 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce25 = 1'b1;
    end else begin
        cipher_0_ssbox_ce25 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce26 = 1'b1;
    end else begin
        cipher_0_ssbox_ce26 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce27 = 1'b1;
    end else begin
        cipher_0_ssbox_ce27 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce28 = 1'b1;
    end else begin
        cipher_0_ssbox_ce28 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce29 = 1'b1;
    end else begin
        cipher_0_ssbox_ce29 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce3 = 1'b1;
    end else begin
        cipher_0_ssbox_ce3 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce30 = 1'b1;
    end else begin
        cipher_0_ssbox_ce30 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce31 = 1'b1;
    end else begin
        cipher_0_ssbox_ce31 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce32 = 1'b1;
    end else begin
        cipher_0_ssbox_ce32 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce33 = 1'b1;
    end else begin
        cipher_0_ssbox_ce33 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce34 = 1'b1;
    end else begin
        cipher_0_ssbox_ce34 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce35 = 1'b1;
    end else begin
        cipher_0_ssbox_ce35 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce36 = 1'b1;
    end else begin
        cipher_0_ssbox_ce36 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce37 = 1'b1;
    end else begin
        cipher_0_ssbox_ce37 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce38 = 1'b1;
    end else begin
        cipher_0_ssbox_ce38 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce39 = 1'b1;
    end else begin
        cipher_0_ssbox_ce39 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce4 = 1'b1;
    end else begin
        cipher_0_ssbox_ce4 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce40 = 1'b1;
    end else begin
        cipher_0_ssbox_ce40 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce41 = 1'b1;
    end else begin
        cipher_0_ssbox_ce41 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce42 = 1'b1;
    end else begin
        cipher_0_ssbox_ce42 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce43 = 1'b1;
    end else begin
        cipher_0_ssbox_ce43 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce44 = 1'b1;
    end else begin
        cipher_0_ssbox_ce44 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce45 = 1'b1;
    end else begin
        cipher_0_ssbox_ce45 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce46 = 1'b1;
    end else begin
        cipher_0_ssbox_ce46 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce47 = 1'b1;
    end else begin
        cipher_0_ssbox_ce47 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce48 = 1'b1;
    end else begin
        cipher_0_ssbox_ce48 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce49 = 1'b1;
    end else begin
        cipher_0_ssbox_ce49 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce5 = 1'b1;
    end else begin
        cipher_0_ssbox_ce5 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce50 = 1'b1;
    end else begin
        cipher_0_ssbox_ce50 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce51 = 1'b1;
    end else begin
        cipher_0_ssbox_ce51 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce52 = 1'b1;
    end else begin
        cipher_0_ssbox_ce52 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce53 = 1'b1;
    end else begin
        cipher_0_ssbox_ce53 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce54 = 1'b1;
    end else begin
        cipher_0_ssbox_ce54 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce55 = 1'b1;
    end else begin
        cipher_0_ssbox_ce55 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce56 = 1'b1;
    end else begin
        cipher_0_ssbox_ce56 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce57 = 1'b1;
    end else begin
        cipher_0_ssbox_ce57 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce58 = 1'b1;
    end else begin
        cipher_0_ssbox_ce58 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce59 = 1'b1;
    end else begin
        cipher_0_ssbox_ce59 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce6 = 1'b1;
    end else begin
        cipher_0_ssbox_ce6 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce60 = 1'b1;
    end else begin
        cipher_0_ssbox_ce60 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce61 = 1'b1;
    end else begin
        cipher_0_ssbox_ce61 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce62 = 1'b1;
    end else begin
        cipher_0_ssbox_ce62 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce63 = 1'b1;
    end else begin
        cipher_0_ssbox_ce63 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce64 = 1'b1;
    end else begin
        cipher_0_ssbox_ce64 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce65 = 1'b1;
    end else begin
        cipher_0_ssbox_ce65 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce66 = 1'b1;
    end else begin
        cipher_0_ssbox_ce66 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce67 = 1'b1;
    end else begin
        cipher_0_ssbox_ce67 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce68 = 1'b1;
    end else begin
        cipher_0_ssbox_ce68 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce69 = 1'b1;
    end else begin
        cipher_0_ssbox_ce69 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce7 = 1'b1;
    end else begin
        cipher_0_ssbox_ce7 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce70 = 1'b1;
    end else begin
        cipher_0_ssbox_ce70 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce71 = 1'b1;
    end else begin
        cipher_0_ssbox_ce71 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce72 = 1'b1;
    end else begin
        cipher_0_ssbox_ce72 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce73 = 1'b1;
    end else begin
        cipher_0_ssbox_ce73 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce74 = 1'b1;
    end else begin
        cipher_0_ssbox_ce74 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce75 = 1'b1;
    end else begin
        cipher_0_ssbox_ce75 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce76 = 1'b1;
    end else begin
        cipher_0_ssbox_ce76 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce77 = 1'b1;
    end else begin
        cipher_0_ssbox_ce77 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce78 = 1'b1;
    end else begin
        cipher_0_ssbox_ce78 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce79 = 1'b1;
    end else begin
        cipher_0_ssbox_ce79 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce8 = 1'b1;
    end else begin
        cipher_0_ssbox_ce8 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce80 = 1'b1;
    end else begin
        cipher_0_ssbox_ce80 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce81 = 1'b1;
    end else begin
        cipher_0_ssbox_ce81 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce82 = 1'b1;
    end else begin
        cipher_0_ssbox_ce82 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce83 = 1'b1;
    end else begin
        cipher_0_ssbox_ce83 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce84 = 1'b1;
    end else begin
        cipher_0_ssbox_ce84 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce85 = 1'b1;
    end else begin
        cipher_0_ssbox_ce85 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce86 = 1'b1;
    end else begin
        cipher_0_ssbox_ce86 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce87 = 1'b1;
    end else begin
        cipher_0_ssbox_ce87 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce88 = 1'b1;
    end else begin
        cipher_0_ssbox_ce88 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce89 = 1'b1;
    end else begin
        cipher_0_ssbox_ce89 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce9 = 1'b1;
    end else begin
        cipher_0_ssbox_ce9 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce90 = 1'b1;
    end else begin
        cipher_0_ssbox_ce90 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce91 = 1'b1;
    end else begin
        cipher_0_ssbox_ce91 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce92 = 1'b1;
    end else begin
        cipher_0_ssbox_ce92 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce93 = 1'b1;
    end else begin
        cipher_0_ssbox_ce93 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce94 = 1'b1;
    end else begin
        cipher_0_ssbox_ce94 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce95 = 1'b1;
    end else begin
        cipher_0_ssbox_ce95 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce96 = 1'b1;
    end else begin
        cipher_0_ssbox_ce96 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce97 = 1'b1;
    end else begin
        cipher_0_ssbox_ce97 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce98 = 1'b1;
    end else begin
        cipher_0_ssbox_ce98 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce99 = 1'b1;
    end else begin
        cipher_0_ssbox_ce99 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_state10_pp0_stage0_iter9 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage0_iter10 = ~(1'b1 == 1'b1);

assign ap_block_state12_pp0_stage0_iter11 = ~(1'b1 == 1'b1);

assign ap_block_state13_pp0_stage0_iter12 = ~(1'b1 == 1'b1);

assign ap_block_state14_pp0_stage0_iter13 = ~(1'b1 == 1'b1);

assign ap_block_state15_pp0_stage0_iter14 = ~(1'b1 == 1'b1);

assign ap_block_state16_pp0_stage0_iter15 = ~(1'b1 == 1'b1);

assign ap_block_state17_pp0_stage0_iter16 = ~(1'b1 == 1'b1);

assign ap_block_state18_pp0_stage0_iter17 = ~(1'b1 == 1'b1);

assign ap_block_state19_pp0_stage0_iter18 = ~(1'b1 == 1'b1);

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state20_pp0_stage0_iter19 = ~(1'b1 == 1'b1);

assign ap_block_state21_pp0_stage0_iter20 = ~(1'b1 == 1'b1);

assign ap_block_state22_pp0_stage0_iter21 = ~(1'b1 == 1'b1);

assign ap_block_state23_pp0_stage0_iter22 = ~(1'b1 == 1'b1);

assign ap_block_state24_pp0_stage0_iter23 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter8 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_enable_reg_pp0_iter0 = ap_start;

assign ap_return = (p_read_1_reg_14078_pp0_iter22_reg ^ p_Result_35_fu_14037_p17);

assign cipher_0_p16box_address0 = zext_ln587_175_fu_13277_p1;

assign cipher_0_p16box_address1 = zext_ln587_174_fu_13272_p1;

assign cipher_0_p16box_address10 = zext_ln587_165_fu_13227_p1;

assign cipher_0_p16box_address100 = zext_ln587_75_fu_8247_p1;

assign cipher_0_p16box_address101 = zext_ln587_74_fu_8242_p1;

assign cipher_0_p16box_address102 = zext_ln587_73_fu_8237_p1;

assign cipher_0_p16box_address103 = zext_ln587_72_fu_8232_p1;

assign cipher_0_p16box_address104 = zext_ln587_71_fu_8227_p1;

assign cipher_0_p16box_address105 = zext_ln587_70_fu_8222_p1;

assign cipher_0_p16box_address106 = zext_ln587_69_fu_8217_p1;

assign cipher_0_p16box_address107 = zext_ln587_68_fu_8212_p1;

assign cipher_0_p16box_address108 = zext_ln587_67_fu_8207_p1;

assign cipher_0_p16box_address109 = zext_ln587_66_fu_8202_p1;

assign cipher_0_p16box_address11 = zext_ln587_164_fu_13222_p1;

assign cipher_0_p16box_address110 = zext_ln587_65_fu_8197_p1;

assign cipher_0_p16box_address111 = zext_ln587_64_fu_8192_p1;

assign cipher_0_p16box_address112 = zext_ln587_63_fu_7432_p1;

assign cipher_0_p16box_address113 = zext_ln587_62_fu_7427_p1;

assign cipher_0_p16box_address114 = zext_ln587_61_fu_7422_p1;

assign cipher_0_p16box_address115 = zext_ln587_60_fu_7417_p1;

assign cipher_0_p16box_address116 = zext_ln587_59_fu_7412_p1;

assign cipher_0_p16box_address117 = zext_ln587_58_fu_7407_p1;

assign cipher_0_p16box_address118 = zext_ln587_57_fu_7402_p1;

assign cipher_0_p16box_address119 = zext_ln587_56_fu_7397_p1;

assign cipher_0_p16box_address12 = zext_ln587_163_fu_13217_p1;

assign cipher_0_p16box_address120 = zext_ln587_55_fu_7392_p1;

assign cipher_0_p16box_address121 = zext_ln587_54_fu_7387_p1;

assign cipher_0_p16box_address122 = zext_ln587_53_fu_7382_p1;

assign cipher_0_p16box_address123 = zext_ln587_52_fu_7377_p1;

assign cipher_0_p16box_address124 = zext_ln587_51_fu_7372_p1;

assign cipher_0_p16box_address125 = zext_ln587_50_fu_7367_p1;

assign cipher_0_p16box_address126 = zext_ln587_49_fu_7362_p1;

assign cipher_0_p16box_address127 = zext_ln587_48_fu_7357_p1;

assign cipher_0_p16box_address128 = zext_ln587_47_fu_6597_p1;

assign cipher_0_p16box_address129 = zext_ln587_46_fu_6592_p1;

assign cipher_0_p16box_address13 = zext_ln587_162_fu_13212_p1;

assign cipher_0_p16box_address130 = zext_ln587_45_fu_6587_p1;

assign cipher_0_p16box_address131 = zext_ln587_44_fu_6582_p1;

assign cipher_0_p16box_address132 = zext_ln587_43_fu_6577_p1;

assign cipher_0_p16box_address133 = zext_ln587_42_fu_6572_p1;

assign cipher_0_p16box_address134 = zext_ln587_41_fu_6567_p1;

assign cipher_0_p16box_address135 = zext_ln587_40_fu_6562_p1;

assign cipher_0_p16box_address136 = zext_ln587_39_fu_6557_p1;

assign cipher_0_p16box_address137 = zext_ln587_38_fu_6552_p1;

assign cipher_0_p16box_address138 = zext_ln587_37_fu_6547_p1;

assign cipher_0_p16box_address139 = zext_ln587_36_fu_6542_p1;

assign cipher_0_p16box_address14 = zext_ln587_161_fu_13207_p1;

assign cipher_0_p16box_address140 = zext_ln587_35_fu_6537_p1;

assign cipher_0_p16box_address141 = zext_ln587_34_fu_6532_p1;

assign cipher_0_p16box_address142 = zext_ln587_33_fu_6527_p1;

assign cipher_0_p16box_address143 = zext_ln587_32_fu_6522_p1;

assign cipher_0_p16box_address144 = zext_ln587_31_fu_5762_p1;

assign cipher_0_p16box_address145 = zext_ln587_30_fu_5757_p1;

assign cipher_0_p16box_address146 = zext_ln587_29_fu_5752_p1;

assign cipher_0_p16box_address147 = zext_ln587_28_fu_5747_p1;

assign cipher_0_p16box_address148 = zext_ln587_27_fu_5742_p1;

assign cipher_0_p16box_address149 = zext_ln587_26_fu_5737_p1;

assign cipher_0_p16box_address15 = zext_ln587_160_fu_13202_p1;

assign cipher_0_p16box_address150 = zext_ln587_25_fu_5732_p1;

assign cipher_0_p16box_address151 = zext_ln587_24_fu_5727_p1;

assign cipher_0_p16box_address152 = zext_ln587_23_fu_5722_p1;

assign cipher_0_p16box_address153 = zext_ln587_22_fu_5717_p1;

assign cipher_0_p16box_address154 = zext_ln587_21_fu_5712_p1;

assign cipher_0_p16box_address155 = zext_ln587_20_fu_5707_p1;

assign cipher_0_p16box_address156 = zext_ln587_19_fu_5702_p1;

assign cipher_0_p16box_address157 = zext_ln587_18_fu_5697_p1;

assign cipher_0_p16box_address158 = zext_ln587_17_fu_5692_p1;

assign cipher_0_p16box_address159 = zext_ln587_16_fu_5687_p1;

assign cipher_0_p16box_address16 = zext_ln587_159_fu_12442_p1;

assign cipher_0_p16box_address160 = zext_ln587_15_fu_4927_p1;

assign cipher_0_p16box_address161 = zext_ln587_14_fu_4922_p1;

assign cipher_0_p16box_address162 = zext_ln587_13_fu_4917_p1;

assign cipher_0_p16box_address163 = zext_ln587_12_fu_4912_p1;

assign cipher_0_p16box_address164 = zext_ln587_11_fu_4907_p1;

assign cipher_0_p16box_address165 = zext_ln587_10_fu_4902_p1;

assign cipher_0_p16box_address166 = zext_ln587_9_fu_4897_p1;

assign cipher_0_p16box_address167 = zext_ln587_8_fu_4892_p1;

assign cipher_0_p16box_address168 = zext_ln587_7_fu_4887_p1;

assign cipher_0_p16box_address169 = zext_ln587_6_fu_4882_p1;

assign cipher_0_p16box_address17 = zext_ln587_158_fu_12437_p1;

assign cipher_0_p16box_address170 = zext_ln587_5_fu_4877_p1;

assign cipher_0_p16box_address171 = zext_ln587_4_fu_4872_p1;

assign cipher_0_p16box_address172 = zext_ln587_3_fu_4867_p1;

assign cipher_0_p16box_address173 = zext_ln587_2_fu_4862_p1;

assign cipher_0_p16box_address174 = zext_ln587_1_fu_4857_p1;

assign cipher_0_p16box_address175 = zext_ln587_fu_4852_p1;

assign cipher_0_p16box_address18 = zext_ln587_157_fu_12432_p1;

assign cipher_0_p16box_address19 = zext_ln587_156_fu_12427_p1;

assign cipher_0_p16box_address2 = zext_ln587_173_fu_13267_p1;

assign cipher_0_p16box_address20 = zext_ln587_155_fu_12422_p1;

assign cipher_0_p16box_address21 = zext_ln587_154_fu_12417_p1;

assign cipher_0_p16box_address22 = zext_ln587_153_fu_12412_p1;

assign cipher_0_p16box_address23 = zext_ln587_152_fu_12407_p1;

assign cipher_0_p16box_address24 = zext_ln587_151_fu_12402_p1;

assign cipher_0_p16box_address25 = zext_ln587_150_fu_12397_p1;

assign cipher_0_p16box_address26 = zext_ln587_149_fu_12392_p1;

assign cipher_0_p16box_address27 = zext_ln587_148_fu_12387_p1;

assign cipher_0_p16box_address28 = zext_ln587_147_fu_12382_p1;

assign cipher_0_p16box_address29 = zext_ln587_146_fu_12377_p1;

assign cipher_0_p16box_address3 = zext_ln587_172_fu_13262_p1;

assign cipher_0_p16box_address30 = zext_ln587_145_fu_12372_p1;

assign cipher_0_p16box_address31 = zext_ln587_144_fu_12367_p1;

assign cipher_0_p16box_address32 = zext_ln587_143_fu_11607_p1;

assign cipher_0_p16box_address33 = zext_ln587_142_fu_11602_p1;

assign cipher_0_p16box_address34 = zext_ln587_141_fu_11597_p1;

assign cipher_0_p16box_address35 = zext_ln587_140_fu_11592_p1;

assign cipher_0_p16box_address36 = zext_ln587_139_fu_11587_p1;

assign cipher_0_p16box_address37 = zext_ln587_138_fu_11582_p1;

assign cipher_0_p16box_address38 = zext_ln587_137_fu_11577_p1;

assign cipher_0_p16box_address39 = zext_ln587_136_fu_11572_p1;

assign cipher_0_p16box_address4 = zext_ln587_171_fu_13257_p1;

assign cipher_0_p16box_address40 = zext_ln587_135_fu_11567_p1;

assign cipher_0_p16box_address41 = zext_ln587_134_fu_11562_p1;

assign cipher_0_p16box_address42 = zext_ln587_133_fu_11557_p1;

assign cipher_0_p16box_address43 = zext_ln587_132_fu_11552_p1;

assign cipher_0_p16box_address44 = zext_ln587_131_fu_11547_p1;

assign cipher_0_p16box_address45 = zext_ln587_130_fu_11542_p1;

assign cipher_0_p16box_address46 = zext_ln587_129_fu_11537_p1;

assign cipher_0_p16box_address47 = zext_ln587_128_fu_11532_p1;

assign cipher_0_p16box_address48 = zext_ln587_127_fu_10772_p1;

assign cipher_0_p16box_address49 = zext_ln587_126_fu_10767_p1;

assign cipher_0_p16box_address5 = zext_ln587_170_fu_13252_p1;

assign cipher_0_p16box_address50 = zext_ln587_125_fu_10762_p1;

assign cipher_0_p16box_address51 = zext_ln587_124_fu_10757_p1;

assign cipher_0_p16box_address52 = zext_ln587_123_fu_10752_p1;

assign cipher_0_p16box_address53 = zext_ln587_122_fu_10747_p1;

assign cipher_0_p16box_address54 = zext_ln587_121_fu_10742_p1;

assign cipher_0_p16box_address55 = zext_ln587_120_fu_10737_p1;

assign cipher_0_p16box_address56 = zext_ln587_119_fu_10732_p1;

assign cipher_0_p16box_address57 = zext_ln587_118_fu_10727_p1;

assign cipher_0_p16box_address58 = zext_ln587_117_fu_10722_p1;

assign cipher_0_p16box_address59 = zext_ln587_116_fu_10717_p1;

assign cipher_0_p16box_address6 = zext_ln587_169_fu_13247_p1;

assign cipher_0_p16box_address60 = zext_ln587_115_fu_10712_p1;

assign cipher_0_p16box_address61 = zext_ln587_114_fu_10707_p1;

assign cipher_0_p16box_address62 = zext_ln587_113_fu_10702_p1;

assign cipher_0_p16box_address63 = zext_ln587_112_fu_10697_p1;

assign cipher_0_p16box_address64 = zext_ln587_111_fu_9937_p1;

assign cipher_0_p16box_address65 = zext_ln587_110_fu_9932_p1;

assign cipher_0_p16box_address66 = zext_ln587_109_fu_9927_p1;

assign cipher_0_p16box_address67 = zext_ln587_108_fu_9922_p1;

assign cipher_0_p16box_address68 = zext_ln587_107_fu_9917_p1;

assign cipher_0_p16box_address69 = zext_ln587_106_fu_9912_p1;

assign cipher_0_p16box_address7 = zext_ln587_168_fu_13242_p1;

assign cipher_0_p16box_address70 = zext_ln587_105_fu_9907_p1;

assign cipher_0_p16box_address71 = zext_ln587_104_fu_9902_p1;

assign cipher_0_p16box_address72 = zext_ln587_103_fu_9897_p1;

assign cipher_0_p16box_address73 = zext_ln587_102_fu_9892_p1;

assign cipher_0_p16box_address74 = zext_ln587_101_fu_9887_p1;

assign cipher_0_p16box_address75 = zext_ln587_100_fu_9882_p1;

assign cipher_0_p16box_address76 = zext_ln587_99_fu_9877_p1;

assign cipher_0_p16box_address77 = zext_ln587_98_fu_9872_p1;

assign cipher_0_p16box_address78 = zext_ln587_97_fu_9867_p1;

assign cipher_0_p16box_address79 = zext_ln587_96_fu_9862_p1;

assign cipher_0_p16box_address8 = zext_ln587_167_fu_13237_p1;

assign cipher_0_p16box_address80 = zext_ln587_95_fu_9102_p1;

assign cipher_0_p16box_address81 = zext_ln587_94_fu_9097_p1;

assign cipher_0_p16box_address82 = zext_ln587_93_fu_9092_p1;

assign cipher_0_p16box_address83 = zext_ln587_92_fu_9087_p1;

assign cipher_0_p16box_address84 = zext_ln587_91_fu_9082_p1;

assign cipher_0_p16box_address85 = zext_ln587_90_fu_9077_p1;

assign cipher_0_p16box_address86 = zext_ln587_89_fu_9072_p1;

assign cipher_0_p16box_address87 = zext_ln587_88_fu_9067_p1;

assign cipher_0_p16box_address88 = zext_ln587_87_fu_9062_p1;

assign cipher_0_p16box_address89 = zext_ln587_86_fu_9057_p1;

assign cipher_0_p16box_address9 = zext_ln587_166_fu_13232_p1;

assign cipher_0_p16box_address90 = zext_ln587_85_fu_9052_p1;

assign cipher_0_p16box_address91 = zext_ln587_84_fu_9047_p1;

assign cipher_0_p16box_address92 = zext_ln587_83_fu_9042_p1;

assign cipher_0_p16box_address93 = zext_ln587_82_fu_9037_p1;

assign cipher_0_p16box_address94 = zext_ln587_81_fu_9032_p1;

assign cipher_0_p16box_address95 = zext_ln587_80_fu_9027_p1;

assign cipher_0_p16box_address96 = zext_ln587_79_fu_8267_p1;

assign cipher_0_p16box_address97 = zext_ln587_78_fu_8262_p1;

assign cipher_0_p16box_address98 = zext_ln587_77_fu_8257_p1;

assign cipher_0_p16box_address99 = zext_ln587_76_fu_8252_p1;

assign cipher_0_ssbox_address0 = zext_ln708_194_fu_14032_p1;

assign cipher_0_ssbox_address1 = zext_ln708_193_fu_14017_p1;

assign cipher_0_ssbox_address10 = zext_ln708_184_fu_13882_p1;

assign cipher_0_ssbox_address100 = zext_ln708_94_fu_8962_p1;

assign cipher_0_ssbox_address101 = zext_ln708_93_fu_8947_p1;

assign cipher_0_ssbox_address102 = zext_ln708_92_fu_8932_p1;

assign cipher_0_ssbox_address103 = zext_ln708_91_fu_8917_p1;

assign cipher_0_ssbox_address104 = zext_ln708_90_fu_8902_p1;

assign cipher_0_ssbox_address105 = zext_ln708_89_fu_8887_p1;

assign cipher_0_ssbox_address106 = zext_ln708_88_fu_8872_p1;

assign cipher_0_ssbox_address107 = zext_ln708_87_fu_8857_p1;

assign cipher_0_ssbox_address108 = zext_ln708_86_fu_8842_p1;

assign cipher_0_ssbox_address109 = zext_ln708_85_fu_8827_p1;

assign cipher_0_ssbox_address11 = zext_ln708_183_fu_13867_p1;

assign cipher_0_ssbox_address110 = zext_ln708_84_fu_8812_p1;

assign cipher_0_ssbox_address111 = zext_ln708_83_fu_8797_p1;

assign cipher_0_ssbox_address112 = zext_ln708_82_fu_8187_p1;

assign cipher_0_ssbox_address113 = zext_ln708_81_fu_8172_p1;

assign cipher_0_ssbox_address114 = zext_ln708_80_fu_8157_p1;

assign cipher_0_ssbox_address115 = zext_ln708_79_fu_8142_p1;

assign cipher_0_ssbox_address116 = zext_ln708_78_fu_8127_p1;

assign cipher_0_ssbox_address117 = zext_ln708_77_fu_8112_p1;

assign cipher_0_ssbox_address118 = zext_ln708_76_fu_8097_p1;

assign cipher_0_ssbox_address119 = zext_ln708_75_fu_8082_p1;

assign cipher_0_ssbox_address12 = zext_ln708_182_fu_13852_p1;

assign cipher_0_ssbox_address120 = zext_ln708_74_fu_8067_p1;

assign cipher_0_ssbox_address121 = zext_ln708_73_fu_8052_p1;

assign cipher_0_ssbox_address122 = zext_ln708_72_fu_8037_p1;

assign cipher_0_ssbox_address123 = zext_ln708_71_fu_8022_p1;

assign cipher_0_ssbox_address124 = zext_ln708_70_fu_8007_p1;

assign cipher_0_ssbox_address125 = zext_ln708_69_fu_7992_p1;

assign cipher_0_ssbox_address126 = zext_ln708_68_fu_7977_p1;

assign cipher_0_ssbox_address127 = zext_ln708_67_fu_7962_p1;

assign cipher_0_ssbox_address128 = zext_ln708_66_fu_7352_p1;

assign cipher_0_ssbox_address129 = zext_ln708_65_fu_7337_p1;

assign cipher_0_ssbox_address13 = zext_ln708_181_fu_13837_p1;

assign cipher_0_ssbox_address130 = zext_ln708_64_fu_7322_p1;

assign cipher_0_ssbox_address131 = zext_ln708_63_fu_7307_p1;

assign cipher_0_ssbox_address132 = zext_ln708_62_fu_7292_p1;

assign cipher_0_ssbox_address133 = zext_ln708_61_fu_7277_p1;

assign cipher_0_ssbox_address134 = zext_ln708_60_fu_7262_p1;

assign cipher_0_ssbox_address135 = zext_ln708_59_fu_7247_p1;

assign cipher_0_ssbox_address136 = zext_ln708_58_fu_7232_p1;

assign cipher_0_ssbox_address137 = zext_ln708_57_fu_7217_p1;

assign cipher_0_ssbox_address138 = zext_ln708_56_fu_7202_p1;

assign cipher_0_ssbox_address139 = zext_ln708_55_fu_7187_p1;

assign cipher_0_ssbox_address14 = zext_ln708_180_fu_13822_p1;

assign cipher_0_ssbox_address140 = zext_ln708_54_fu_7172_p1;

assign cipher_0_ssbox_address141 = zext_ln708_53_fu_7157_p1;

assign cipher_0_ssbox_address142 = zext_ln708_52_fu_7142_p1;

assign cipher_0_ssbox_address143 = zext_ln708_51_fu_7127_p1;

assign cipher_0_ssbox_address144 = zext_ln708_50_fu_6517_p1;

assign cipher_0_ssbox_address145 = zext_ln708_49_fu_6502_p1;

assign cipher_0_ssbox_address146 = zext_ln708_48_fu_6487_p1;

assign cipher_0_ssbox_address147 = zext_ln708_47_fu_6472_p1;

assign cipher_0_ssbox_address148 = zext_ln708_46_fu_6457_p1;

assign cipher_0_ssbox_address149 = zext_ln708_45_fu_6442_p1;

assign cipher_0_ssbox_address15 = zext_ln708_179_fu_13807_p1;

assign cipher_0_ssbox_address150 = zext_ln708_44_fu_6427_p1;

assign cipher_0_ssbox_address151 = zext_ln708_43_fu_6412_p1;

assign cipher_0_ssbox_address152 = zext_ln708_42_fu_6397_p1;

assign cipher_0_ssbox_address153 = zext_ln708_41_fu_6382_p1;

assign cipher_0_ssbox_address154 = zext_ln708_40_fu_6367_p1;

assign cipher_0_ssbox_address155 = zext_ln708_39_fu_6352_p1;

assign cipher_0_ssbox_address156 = zext_ln708_38_fu_6337_p1;

assign cipher_0_ssbox_address157 = zext_ln708_37_fu_6322_p1;

assign cipher_0_ssbox_address158 = zext_ln708_36_fu_6307_p1;

assign cipher_0_ssbox_address159 = zext_ln708_35_fu_6292_p1;

assign cipher_0_ssbox_address16 = zext_ln708_178_fu_13197_p1;

assign cipher_0_ssbox_address160 = zext_ln708_34_fu_5682_p1;

assign cipher_0_ssbox_address161 = zext_ln708_33_fu_5667_p1;

assign cipher_0_ssbox_address162 = zext_ln708_32_fu_5652_p1;

assign cipher_0_ssbox_address163 = zext_ln708_31_fu_5637_p1;

assign cipher_0_ssbox_address164 = zext_ln708_30_fu_5622_p1;

assign cipher_0_ssbox_address165 = zext_ln708_29_fu_5607_p1;

assign cipher_0_ssbox_address166 = zext_ln708_28_fu_5592_p1;

assign cipher_0_ssbox_address167 = zext_ln708_27_fu_5577_p1;

assign cipher_0_ssbox_address168 = zext_ln708_26_fu_5562_p1;

assign cipher_0_ssbox_address169 = zext_ln708_25_fu_5547_p1;

assign cipher_0_ssbox_address17 = zext_ln708_177_fu_13182_p1;

assign cipher_0_ssbox_address170 = zext_ln708_24_fu_5532_p1;

assign cipher_0_ssbox_address171 = zext_ln708_23_fu_5517_p1;

assign cipher_0_ssbox_address172 = zext_ln708_22_fu_5502_p1;

assign cipher_0_ssbox_address173 = zext_ln708_21_fu_5487_p1;

assign cipher_0_ssbox_address174 = zext_ln708_20_fu_5472_p1;

assign cipher_0_ssbox_address175 = zext_ln708_19_fu_5457_p1;

assign cipher_0_ssbox_address176 = zext_ln708_18_fu_4847_p1;

assign cipher_0_ssbox_address177 = zext_ln708_17_fu_4832_p1;

assign cipher_0_ssbox_address178 = zext_ln708_16_fu_4817_p1;

assign cipher_0_ssbox_address179 = zext_ln708_15_fu_4802_p1;

assign cipher_0_ssbox_address18 = zext_ln708_176_fu_13167_p1;

assign cipher_0_ssbox_address180 = zext_ln708_14_fu_4787_p1;

assign cipher_0_ssbox_address181 = zext_ln708_13_fu_4772_p1;

assign cipher_0_ssbox_address182 = zext_ln708_12_fu_4757_p1;

assign cipher_0_ssbox_address183 = zext_ln708_11_fu_4742_p1;

assign cipher_0_ssbox_address184 = zext_ln708_10_fu_4727_p1;

assign cipher_0_ssbox_address185 = zext_ln708_9_fu_4712_p1;

assign cipher_0_ssbox_address186 = zext_ln708_8_fu_4697_p1;

assign cipher_0_ssbox_address187 = zext_ln708_7_fu_4682_p1;

assign cipher_0_ssbox_address188 = zext_ln708_6_fu_4667_p1;

assign cipher_0_ssbox_address189 = zext_ln708_5_fu_4652_p1;

assign cipher_0_ssbox_address19 = zext_ln708_175_fu_13152_p1;

assign cipher_0_ssbox_address190 = zext_ln708_4_fu_4637_p1;

assign cipher_0_ssbox_address191 = zext_ln708_fu_4622_p1;

assign cipher_0_ssbox_address2 = zext_ln708_192_fu_14002_p1;

assign cipher_0_ssbox_address20 = zext_ln708_174_fu_13137_p1;

assign cipher_0_ssbox_address21 = zext_ln708_173_fu_13122_p1;

assign cipher_0_ssbox_address22 = zext_ln708_172_fu_13107_p1;

assign cipher_0_ssbox_address23 = zext_ln708_171_fu_13092_p1;

assign cipher_0_ssbox_address24 = zext_ln708_170_fu_13077_p1;

assign cipher_0_ssbox_address25 = zext_ln708_169_fu_13062_p1;

assign cipher_0_ssbox_address26 = zext_ln708_168_fu_13047_p1;

assign cipher_0_ssbox_address27 = zext_ln708_167_fu_13032_p1;

assign cipher_0_ssbox_address28 = zext_ln708_166_fu_13017_p1;

assign cipher_0_ssbox_address29 = zext_ln708_165_fu_13002_p1;

assign cipher_0_ssbox_address3 = zext_ln708_191_fu_13987_p1;

assign cipher_0_ssbox_address30 = zext_ln708_164_fu_12987_p1;

assign cipher_0_ssbox_address31 = zext_ln708_163_fu_12972_p1;

assign cipher_0_ssbox_address32 = zext_ln708_162_fu_12362_p1;

assign cipher_0_ssbox_address33 = zext_ln708_161_fu_12347_p1;

assign cipher_0_ssbox_address34 = zext_ln708_160_fu_12332_p1;

assign cipher_0_ssbox_address35 = zext_ln708_159_fu_12317_p1;

assign cipher_0_ssbox_address36 = zext_ln708_158_fu_12302_p1;

assign cipher_0_ssbox_address37 = zext_ln708_157_fu_12287_p1;

assign cipher_0_ssbox_address38 = zext_ln708_156_fu_12272_p1;

assign cipher_0_ssbox_address39 = zext_ln708_155_fu_12257_p1;

assign cipher_0_ssbox_address4 = zext_ln708_190_fu_13972_p1;

assign cipher_0_ssbox_address40 = zext_ln708_154_fu_12242_p1;

assign cipher_0_ssbox_address41 = zext_ln708_153_fu_12227_p1;

assign cipher_0_ssbox_address42 = zext_ln708_152_fu_12212_p1;

assign cipher_0_ssbox_address43 = zext_ln708_151_fu_12197_p1;

assign cipher_0_ssbox_address44 = zext_ln708_150_fu_12182_p1;

assign cipher_0_ssbox_address45 = zext_ln708_149_fu_12167_p1;

assign cipher_0_ssbox_address46 = zext_ln708_148_fu_12152_p1;

assign cipher_0_ssbox_address47 = zext_ln708_147_fu_12137_p1;

assign cipher_0_ssbox_address48 = zext_ln708_146_fu_11527_p1;

assign cipher_0_ssbox_address49 = zext_ln708_145_fu_11512_p1;

assign cipher_0_ssbox_address5 = zext_ln708_189_fu_13957_p1;

assign cipher_0_ssbox_address50 = zext_ln708_144_fu_11497_p1;

assign cipher_0_ssbox_address51 = zext_ln708_143_fu_11482_p1;

assign cipher_0_ssbox_address52 = zext_ln708_142_fu_11467_p1;

assign cipher_0_ssbox_address53 = zext_ln708_141_fu_11452_p1;

assign cipher_0_ssbox_address54 = zext_ln708_140_fu_11437_p1;

assign cipher_0_ssbox_address55 = zext_ln708_139_fu_11422_p1;

assign cipher_0_ssbox_address56 = zext_ln708_138_fu_11407_p1;

assign cipher_0_ssbox_address57 = zext_ln708_137_fu_11392_p1;

assign cipher_0_ssbox_address58 = zext_ln708_136_fu_11377_p1;

assign cipher_0_ssbox_address59 = zext_ln708_135_fu_11362_p1;

assign cipher_0_ssbox_address6 = zext_ln708_188_fu_13942_p1;

assign cipher_0_ssbox_address60 = zext_ln708_134_fu_11347_p1;

assign cipher_0_ssbox_address61 = zext_ln708_133_fu_11332_p1;

assign cipher_0_ssbox_address62 = zext_ln708_132_fu_11317_p1;

assign cipher_0_ssbox_address63 = zext_ln708_131_fu_11302_p1;

assign cipher_0_ssbox_address64 = zext_ln708_130_fu_10692_p1;

assign cipher_0_ssbox_address65 = zext_ln708_129_fu_10677_p1;

assign cipher_0_ssbox_address66 = zext_ln708_128_fu_10662_p1;

assign cipher_0_ssbox_address67 = zext_ln708_127_fu_10647_p1;

assign cipher_0_ssbox_address68 = zext_ln708_126_fu_10632_p1;

assign cipher_0_ssbox_address69 = zext_ln708_125_fu_10617_p1;

assign cipher_0_ssbox_address7 = zext_ln708_187_fu_13927_p1;

assign cipher_0_ssbox_address70 = zext_ln708_124_fu_10602_p1;

assign cipher_0_ssbox_address71 = zext_ln708_123_fu_10587_p1;

assign cipher_0_ssbox_address72 = zext_ln708_122_fu_10572_p1;

assign cipher_0_ssbox_address73 = zext_ln708_121_fu_10557_p1;

assign cipher_0_ssbox_address74 = zext_ln708_120_fu_10542_p1;

assign cipher_0_ssbox_address75 = zext_ln708_119_fu_10527_p1;

assign cipher_0_ssbox_address76 = zext_ln708_118_fu_10512_p1;

assign cipher_0_ssbox_address77 = zext_ln708_117_fu_10497_p1;

assign cipher_0_ssbox_address78 = zext_ln708_116_fu_10482_p1;

assign cipher_0_ssbox_address79 = zext_ln708_115_fu_10467_p1;

assign cipher_0_ssbox_address8 = zext_ln708_186_fu_13912_p1;

assign cipher_0_ssbox_address80 = zext_ln708_114_fu_9857_p1;

assign cipher_0_ssbox_address81 = zext_ln708_113_fu_9842_p1;

assign cipher_0_ssbox_address82 = zext_ln708_112_fu_9827_p1;

assign cipher_0_ssbox_address83 = zext_ln708_111_fu_9812_p1;

assign cipher_0_ssbox_address84 = zext_ln708_110_fu_9797_p1;

assign cipher_0_ssbox_address85 = zext_ln708_109_fu_9782_p1;

assign cipher_0_ssbox_address86 = zext_ln708_108_fu_9767_p1;

assign cipher_0_ssbox_address87 = zext_ln708_107_fu_9752_p1;

assign cipher_0_ssbox_address88 = zext_ln708_106_fu_9737_p1;

assign cipher_0_ssbox_address89 = zext_ln708_105_fu_9722_p1;

assign cipher_0_ssbox_address9 = zext_ln708_185_fu_13897_p1;

assign cipher_0_ssbox_address90 = zext_ln708_104_fu_9707_p1;

assign cipher_0_ssbox_address91 = zext_ln708_103_fu_9692_p1;

assign cipher_0_ssbox_address92 = zext_ln708_102_fu_9677_p1;

assign cipher_0_ssbox_address93 = zext_ln708_101_fu_9662_p1;

assign cipher_0_ssbox_address94 = zext_ln708_100_fu_9647_p1;

assign cipher_0_ssbox_address95 = zext_ln708_99_fu_9632_p1;

assign cipher_0_ssbox_address96 = zext_ln708_98_fu_9022_p1;

assign cipher_0_ssbox_address97 = zext_ln708_97_fu_9007_p1;

assign cipher_0_ssbox_address98 = zext_ln708_96_fu_8992_p1;

assign cipher_0_ssbox_address99 = zext_ln708_95_fu_8977_p1;

assign p_Result_25_fu_6247_p17 = {{{{{{{{{{{{{{{{xor_ln1545_100_fu_6241_p2}, {xor_ln1545_97_fu_6225_p2}}, {xor_ln1545_94_fu_6209_p2}}, {xor_ln1545_91_fu_6193_p2}}, {xor_ln1545_88_fu_6177_p2}}, {xor_ln1545_85_fu_6161_p2}}, {xor_ln1545_82_fu_6145_p2}}, {xor_ln1545_79_fu_6129_p2}}, {xor_ln1545_76_fu_6113_p2}}, {xor_ln1545_73_fu_6097_p2}}, {xor_ln1545_70_fu_6081_p2}}, {xor_ln1545_67_fu_6065_p2}}, {xor_ln1545_64_fu_6049_p2}}, {xor_ln1545_61_fu_6033_p2}}, {xor_ln1545_58_fu_6017_p2}}, {xor_ln1545_55_fu_6001_p2}};

assign p_Result_26_fu_7082_p17 = {{{{{{{{{{{{{{{{xor_ln1545_148_fu_7076_p2}, {xor_ln1545_145_fu_7060_p2}}, {xor_ln1545_142_fu_7044_p2}}, {xor_ln1545_139_fu_7028_p2}}, {xor_ln1545_136_fu_7012_p2}}, {xor_ln1545_133_fu_6996_p2}}, {xor_ln1545_130_fu_6980_p2}}, {xor_ln1545_127_fu_6964_p2}}, {xor_ln1545_124_fu_6948_p2}}, {xor_ln1545_121_fu_6932_p2}}, {xor_ln1545_118_fu_6916_p2}}, {xor_ln1545_115_fu_6900_p2}}, {xor_ln1545_112_fu_6884_p2}}, {xor_ln1545_109_fu_6868_p2}}, {xor_ln1545_106_fu_6852_p2}}, {xor_ln1545_103_fu_6836_p2}};

assign p_Result_27_fu_7917_p17 = {{{{{{{{{{{{{{{{xor_ln1545_196_fu_7911_p2}, {xor_ln1545_193_fu_7895_p2}}, {xor_ln1545_190_fu_7879_p2}}, {xor_ln1545_187_fu_7863_p2}}, {xor_ln1545_184_fu_7847_p2}}, {xor_ln1545_181_fu_7831_p2}}, {xor_ln1545_178_fu_7815_p2}}, {xor_ln1545_175_fu_7799_p2}}, {xor_ln1545_172_fu_7783_p2}}, {xor_ln1545_169_fu_7767_p2}}, {xor_ln1545_166_fu_7751_p2}}, {xor_ln1545_163_fu_7735_p2}}, {xor_ln1545_160_fu_7719_p2}}, {xor_ln1545_157_fu_7703_p2}}, {xor_ln1545_154_fu_7687_p2}}, {xor_ln1545_151_fu_7671_p2}};

assign p_Result_28_fu_8752_p17 = {{{{{{{{{{{{{{{{xor_ln1545_244_fu_8746_p2}, {xor_ln1545_241_fu_8730_p2}}, {xor_ln1545_238_fu_8714_p2}}, {xor_ln1545_235_fu_8698_p2}}, {xor_ln1545_232_fu_8682_p2}}, {xor_ln1545_229_fu_8666_p2}}, {xor_ln1545_226_fu_8650_p2}}, {xor_ln1545_223_fu_8634_p2}}, {xor_ln1545_220_fu_8618_p2}}, {xor_ln1545_217_fu_8602_p2}}, {xor_ln1545_214_fu_8586_p2}}, {xor_ln1545_211_fu_8570_p2}}, {xor_ln1545_208_fu_8554_p2}}, {xor_ln1545_205_fu_8538_p2}}, {xor_ln1545_202_fu_8522_p2}}, {xor_ln1545_199_fu_8506_p2}};

assign p_Result_29_fu_9587_p17 = {{{{{{{{{{{{{{{{xor_ln1545_292_fu_9581_p2}, {xor_ln1545_289_fu_9565_p2}}, {xor_ln1545_286_fu_9549_p2}}, {xor_ln1545_283_fu_9533_p2}}, {xor_ln1545_280_fu_9517_p2}}, {xor_ln1545_277_fu_9501_p2}}, {xor_ln1545_274_fu_9485_p2}}, {xor_ln1545_271_fu_9469_p2}}, {xor_ln1545_268_fu_9453_p2}}, {xor_ln1545_265_fu_9437_p2}}, {xor_ln1545_262_fu_9421_p2}}, {xor_ln1545_259_fu_9405_p2}}, {xor_ln1545_256_fu_9389_p2}}, {xor_ln1545_253_fu_9373_p2}}, {xor_ln1545_250_fu_9357_p2}}, {xor_ln1545_247_fu_9341_p2}};

assign p_Result_30_fu_10422_p17 = {{{{{{{{{{{{{{{{xor_ln1545_340_fu_10416_p2}, {xor_ln1545_337_fu_10400_p2}}, {xor_ln1545_334_fu_10384_p2}}, {xor_ln1545_331_fu_10368_p2}}, {xor_ln1545_328_fu_10352_p2}}, {xor_ln1545_325_fu_10336_p2}}, {xor_ln1545_322_fu_10320_p2}}, {xor_ln1545_319_fu_10304_p2}}, {xor_ln1545_316_fu_10288_p2}}, {xor_ln1545_313_fu_10272_p2}}, {xor_ln1545_310_fu_10256_p2}}, {xor_ln1545_307_fu_10240_p2}}, {xor_ln1545_304_fu_10224_p2}}, {xor_ln1545_301_fu_10208_p2}}, {xor_ln1545_298_fu_10192_p2}}, {xor_ln1545_295_fu_10176_p2}};

assign p_Result_31_fu_11257_p17 = {{{{{{{{{{{{{{{{xor_ln1545_388_fu_11251_p2}, {xor_ln1545_385_fu_11235_p2}}, {xor_ln1545_382_fu_11219_p2}}, {xor_ln1545_379_fu_11203_p2}}, {xor_ln1545_376_fu_11187_p2}}, {xor_ln1545_373_fu_11171_p2}}, {xor_ln1545_370_fu_11155_p2}}, {xor_ln1545_367_fu_11139_p2}}, {xor_ln1545_364_fu_11123_p2}}, {xor_ln1545_361_fu_11107_p2}}, {xor_ln1545_358_fu_11091_p2}}, {xor_ln1545_355_fu_11075_p2}}, {xor_ln1545_352_fu_11059_p2}}, {xor_ln1545_349_fu_11043_p2}}, {xor_ln1545_346_fu_11027_p2}}, {xor_ln1545_343_fu_11011_p2}};

assign p_Result_32_fu_12092_p17 = {{{{{{{{{{{{{{{{xor_ln1545_436_fu_12086_p2}, {xor_ln1545_433_fu_12070_p2}}, {xor_ln1545_430_fu_12054_p2}}, {xor_ln1545_427_fu_12038_p2}}, {xor_ln1545_424_fu_12022_p2}}, {xor_ln1545_421_fu_12006_p2}}, {xor_ln1545_418_fu_11990_p2}}, {xor_ln1545_415_fu_11974_p2}}, {xor_ln1545_412_fu_11958_p2}}, {xor_ln1545_409_fu_11942_p2}}, {xor_ln1545_406_fu_11926_p2}}, {xor_ln1545_403_fu_11910_p2}}, {xor_ln1545_400_fu_11894_p2}}, {xor_ln1545_397_fu_11878_p2}}, {xor_ln1545_394_fu_11862_p2}}, {xor_ln1545_391_fu_11846_p2}};

assign p_Result_33_fu_12927_p17 = {{{{{{{{{{{{{{{{xor_ln1545_484_fu_12921_p2}, {xor_ln1545_481_fu_12905_p2}}, {xor_ln1545_478_fu_12889_p2}}, {xor_ln1545_475_fu_12873_p2}}, {xor_ln1545_472_fu_12857_p2}}, {xor_ln1545_469_fu_12841_p2}}, {xor_ln1545_466_fu_12825_p2}}, {xor_ln1545_463_fu_12809_p2}}, {xor_ln1545_460_fu_12793_p2}}, {xor_ln1545_457_fu_12777_p2}}, {xor_ln1545_454_fu_12761_p2}}, {xor_ln1545_451_fu_12745_p2}}, {xor_ln1545_448_fu_12729_p2}}, {xor_ln1545_445_fu_12713_p2}}, {xor_ln1545_442_fu_12697_p2}}, {xor_ln1545_439_fu_12681_p2}};

assign p_Result_34_fu_13762_p17 = {{{{{{{{{{{{{{{{xor_ln1545_532_fu_13756_p2}, {xor_ln1545_529_fu_13740_p2}}, {xor_ln1545_526_fu_13724_p2}}, {xor_ln1545_523_fu_13708_p2}}, {xor_ln1545_520_fu_13692_p2}}, {xor_ln1545_517_fu_13676_p2}}, {xor_ln1545_514_fu_13660_p2}}, {xor_ln1545_511_fu_13644_p2}}, {xor_ln1545_508_fu_13628_p2}}, {xor_ln1545_505_fu_13612_p2}}, {xor_ln1545_502_fu_13596_p2}}, {xor_ln1545_499_fu_13580_p2}}, {xor_ln1545_496_fu_13564_p2}}, {xor_ln1545_493_fu_13548_p2}}, {xor_ln1545_490_fu_13532_p2}}, {xor_ln1545_487_fu_13516_p2}};

assign p_Result_35_fu_14037_p17 = {{{{{{{{{{{{{{{{cipher_0_ssbox_q4}, {cipher_0_ssbox_q9}}, {cipher_0_ssbox_q14}}, {cipher_0_ssbox_q3}}, {cipher_0_ssbox_q8}}, {cipher_0_ssbox_q13}}, {cipher_0_ssbox_q2}}, {cipher_0_ssbox_q7}}, {cipher_0_ssbox_q12}}, {cipher_0_ssbox_q1}}, {cipher_0_ssbox_q6}}, {cipher_0_ssbox_q11}}, {cipher_0_ssbox_q0}}, {cipher_0_ssbox_q5}}, {cipher_0_ssbox_q10}}, {cipher_0_ssbox_q15}};

assign p_Result_s_fu_5412_p17 = {{{{{{{{{{{{{{{{xor_ln1545_52_fu_5406_p2}, {xor_ln1545_49_fu_5390_p2}}, {xor_ln1545_46_fu_5374_p2}}, {xor_ln1545_43_fu_5358_p2}}, {xor_ln1545_40_fu_5342_p2}}, {xor_ln1545_37_fu_5326_p2}}, {xor_ln1545_34_fu_5310_p2}}, {xor_ln1545_31_fu_5294_p2}}, {xor_ln1545_28_fu_5278_p2}}, {xor_ln1545_25_fu_5262_p2}}, {xor_ln1545_22_fu_5246_p2}}, {xor_ln1545_19_fu_5230_p2}}, {xor_ln1545_16_fu_5214_p2}}, {xor_ln1545_13_fu_5198_p2}}, {xor_ln1545_10_fu_5182_p2}}, {xor_ln1545_7_fu_5166_p2}};

assign ret_V_fu_4612_p2 = (plaintext ^ p_read);

assign state_V_24_fu_5448_p2 = (p_read_12_reg_14133_pp0_iter1_reg ^ p_Result_s_fu_5412_p17);

assign state_V_25_fu_6283_p2 = (p_read_11_reg_14128_pp0_iter3_reg ^ p_Result_25_fu_6247_p17);

assign state_V_26_fu_7118_p2 = (p_read_10_reg_14123_pp0_iter5_reg ^ p_Result_26_fu_7082_p17);

assign state_V_27_fu_7953_p2 = (p_read_9_reg_14118_pp0_iter7_reg ^ p_Result_27_fu_7917_p17);

assign state_V_28_fu_8788_p2 = (p_read_8_reg_14113_pp0_iter9_reg ^ p_Result_28_fu_8752_p17);

assign state_V_29_fu_9623_p2 = (p_read_7_reg_14108_pp0_iter11_reg ^ p_Result_29_fu_9587_p17);

assign state_V_30_fu_11293_p2 = (p_read_5_reg_14098_pp0_iter15_reg ^ p_Result_31_fu_11257_p17);

assign state_V_31_fu_12128_p2 = (p_read_4_reg_14093_pp0_iter17_reg ^ p_Result_32_fu_12092_p17);

assign state_V_32_fu_12963_p2 = (p_read_3_reg_14088_pp0_iter19_reg ^ p_Result_33_fu_12927_p17);

assign state_V_33_fu_13798_p2 = (p_read_2_reg_14083_pp0_iter21_reg ^ p_Result_34_fu_13762_p17);

assign state_V_fu_10458_p2 = (p_read_6_reg_14103_pp0_iter13_reg ^ p_Result_30_fu_10422_p17);

assign tmp_100_fu_6746_p4 = {{cipher_0_p16box_q133[15:8]}};

assign tmp_101_fu_6760_p4 = {{cipher_0_p16box_q132[15:8]}};

assign tmp_102_fu_6774_p4 = {{cipher_0_p16box_q131[15:8]}};

assign tmp_103_fu_6788_p4 = {{cipher_0_p16box_q130[15:8]}};

assign tmp_104_fu_6802_p4 = {{cipher_0_p16box_q129[15:8]}};

assign tmp_105_fu_6816_p4 = {{cipher_0_p16box_q128[15:8]}};

assign tmp_106_fu_7132_p4 = {{state_V_26_fu_7118_p2[15:8]}};

assign tmp_107_fu_7147_p4 = {{state_V_26_fu_7118_p2[23:16]}};

assign tmp_108_fu_7162_p4 = {{state_V_26_fu_7118_p2[31:24]}};

assign tmp_109_fu_7177_p4 = {{state_V_26_fu_7118_p2[39:32]}};

assign tmp_110_fu_7192_p4 = {{state_V_26_fu_7118_p2[47:40]}};

assign tmp_111_fu_7207_p4 = {{state_V_26_fu_7118_p2[55:48]}};

assign tmp_112_fu_7222_p4 = {{state_V_26_fu_7118_p2[63:56]}};

assign tmp_113_fu_7237_p4 = {{state_V_26_fu_7118_p2[71:64]}};

assign tmp_114_fu_7252_p4 = {{state_V_26_fu_7118_p2[79:72]}};

assign tmp_115_fu_7267_p4 = {{state_V_26_fu_7118_p2[87:80]}};

assign tmp_116_fu_7282_p4 = {{state_V_26_fu_7118_p2[95:88]}};

assign tmp_117_fu_7297_p4 = {{state_V_26_fu_7118_p2[103:96]}};

assign tmp_118_fu_7312_p4 = {{state_V_26_fu_7118_p2[111:104]}};

assign tmp_119_fu_7327_p4 = {{state_V_26_fu_7118_p2[119:112]}};

assign tmp_120_fu_7342_p4 = {{state_V_26_fu_7118_p2[127:120]}};

assign tmp_121_fu_7441_p4 = {{cipher_0_p16box_q127[15:8]}};

assign tmp_122_fu_7455_p4 = {{cipher_0_p16box_q126[15:8]}};

assign tmp_123_fu_7469_p4 = {{cipher_0_p16box_q125[15:8]}};

assign tmp_124_fu_7483_p4 = {{cipher_0_p16box_q124[15:8]}};

assign tmp_125_fu_7497_p4 = {{cipher_0_p16box_q123[15:8]}};

assign tmp_126_fu_7511_p4 = {{cipher_0_p16box_q122[15:8]}};

assign tmp_127_fu_7525_p4 = {{cipher_0_p16box_q121[15:8]}};

assign tmp_128_fu_7539_p4 = {{cipher_0_p16box_q120[15:8]}};

assign tmp_129_fu_7553_p4 = {{cipher_0_p16box_q119[15:8]}};

assign tmp_130_fu_7567_p4 = {{cipher_0_p16box_q118[15:8]}};

assign tmp_131_fu_7581_p4 = {{cipher_0_p16box_q117[15:8]}};

assign tmp_132_fu_7595_p4 = {{cipher_0_p16box_q116[15:8]}};

assign tmp_133_fu_7609_p4 = {{cipher_0_p16box_q115[15:8]}};

assign tmp_134_fu_7623_p4 = {{cipher_0_p16box_q114[15:8]}};

assign tmp_135_fu_7637_p4 = {{cipher_0_p16box_q113[15:8]}};

assign tmp_136_fu_7651_p4 = {{cipher_0_p16box_q112[15:8]}};

assign tmp_137_fu_7967_p4 = {{state_V_27_fu_7953_p2[15:8]}};

assign tmp_138_fu_7982_p4 = {{state_V_27_fu_7953_p2[23:16]}};

assign tmp_139_fu_7997_p4 = {{state_V_27_fu_7953_p2[31:24]}};

assign tmp_140_fu_8012_p4 = {{state_V_27_fu_7953_p2[39:32]}};

assign tmp_141_fu_8027_p4 = {{state_V_27_fu_7953_p2[47:40]}};

assign tmp_142_fu_8042_p4 = {{state_V_27_fu_7953_p2[55:48]}};

assign tmp_143_fu_8057_p4 = {{state_V_27_fu_7953_p2[63:56]}};

assign tmp_144_fu_8072_p4 = {{state_V_27_fu_7953_p2[71:64]}};

assign tmp_145_fu_8087_p4 = {{state_V_27_fu_7953_p2[79:72]}};

assign tmp_146_fu_8102_p4 = {{state_V_27_fu_7953_p2[87:80]}};

assign tmp_147_fu_8117_p4 = {{state_V_27_fu_7953_p2[95:88]}};

assign tmp_148_fu_8132_p4 = {{state_V_27_fu_7953_p2[103:96]}};

assign tmp_149_fu_8147_p4 = {{state_V_27_fu_7953_p2[111:104]}};

assign tmp_14_fu_4642_p4 = {{ret_V_fu_4612_p2[23:16]}};

assign tmp_150_fu_8162_p4 = {{state_V_27_fu_7953_p2[119:112]}};

assign tmp_151_fu_8177_p4 = {{state_V_27_fu_7953_p2[127:120]}};

assign tmp_152_fu_8276_p4 = {{cipher_0_p16box_q111[15:8]}};

assign tmp_153_fu_8290_p4 = {{cipher_0_p16box_q110[15:8]}};

assign tmp_154_fu_8304_p4 = {{cipher_0_p16box_q109[15:8]}};

assign tmp_155_fu_8318_p4 = {{cipher_0_p16box_q108[15:8]}};

assign tmp_156_fu_8332_p4 = {{cipher_0_p16box_q107[15:8]}};

assign tmp_157_fu_8346_p4 = {{cipher_0_p16box_q106[15:8]}};

assign tmp_158_fu_8360_p4 = {{cipher_0_p16box_q105[15:8]}};

assign tmp_159_fu_8374_p4 = {{cipher_0_p16box_q104[15:8]}};

assign tmp_15_fu_4657_p4 = {{ret_V_fu_4612_p2[31:24]}};

assign tmp_160_fu_8388_p4 = {{cipher_0_p16box_q103[15:8]}};

assign tmp_161_fu_8402_p4 = {{cipher_0_p16box_q102[15:8]}};

assign tmp_162_fu_8416_p4 = {{cipher_0_p16box_q101[15:8]}};

assign tmp_163_fu_8430_p4 = {{cipher_0_p16box_q100[15:8]}};

assign tmp_164_fu_8444_p4 = {{cipher_0_p16box_q99[15:8]}};

assign tmp_165_fu_8458_p4 = {{cipher_0_p16box_q98[15:8]}};

assign tmp_166_fu_8472_p4 = {{cipher_0_p16box_q97[15:8]}};

assign tmp_167_fu_8486_p4 = {{cipher_0_p16box_q96[15:8]}};

assign tmp_168_fu_8802_p4 = {{state_V_28_fu_8788_p2[15:8]}};

assign tmp_169_fu_8817_p4 = {{state_V_28_fu_8788_p2[23:16]}};

assign tmp_16_fu_4672_p4 = {{ret_V_fu_4612_p2[39:32]}};

assign tmp_170_fu_8832_p4 = {{state_V_28_fu_8788_p2[31:24]}};

assign tmp_171_fu_8847_p4 = {{state_V_28_fu_8788_p2[39:32]}};

assign tmp_172_fu_8862_p4 = {{state_V_28_fu_8788_p2[47:40]}};

assign tmp_173_fu_8877_p4 = {{state_V_28_fu_8788_p2[55:48]}};

assign tmp_174_fu_8892_p4 = {{state_V_28_fu_8788_p2[63:56]}};

assign tmp_175_fu_8907_p4 = {{state_V_28_fu_8788_p2[71:64]}};

assign tmp_176_fu_8922_p4 = {{state_V_28_fu_8788_p2[79:72]}};

assign tmp_177_fu_8937_p4 = {{state_V_28_fu_8788_p2[87:80]}};

assign tmp_178_fu_8952_p4 = {{state_V_28_fu_8788_p2[95:88]}};

assign tmp_179_fu_8967_p4 = {{state_V_28_fu_8788_p2[103:96]}};

assign tmp_17_fu_4687_p4 = {{ret_V_fu_4612_p2[47:40]}};

assign tmp_180_fu_8982_p4 = {{state_V_28_fu_8788_p2[111:104]}};

assign tmp_181_fu_8997_p4 = {{state_V_28_fu_8788_p2[119:112]}};

assign tmp_182_fu_9012_p4 = {{state_V_28_fu_8788_p2[127:120]}};

assign tmp_183_fu_9111_p4 = {{cipher_0_p16box_q95[15:8]}};

assign tmp_184_fu_9125_p4 = {{cipher_0_p16box_q94[15:8]}};

assign tmp_185_fu_9139_p4 = {{cipher_0_p16box_q93[15:8]}};

assign tmp_186_fu_9153_p4 = {{cipher_0_p16box_q92[15:8]}};

assign tmp_187_fu_9167_p4 = {{cipher_0_p16box_q91[15:8]}};

assign tmp_188_fu_9181_p4 = {{cipher_0_p16box_q90[15:8]}};

assign tmp_189_fu_9195_p4 = {{cipher_0_p16box_q89[15:8]}};

assign tmp_18_fu_4702_p4 = {{ret_V_fu_4612_p2[55:48]}};

assign tmp_190_fu_9209_p4 = {{cipher_0_p16box_q88[15:8]}};

assign tmp_191_fu_9223_p4 = {{cipher_0_p16box_q87[15:8]}};

assign tmp_192_fu_9237_p4 = {{cipher_0_p16box_q86[15:8]}};

assign tmp_193_fu_9251_p4 = {{cipher_0_p16box_q85[15:8]}};

assign tmp_194_fu_9265_p4 = {{cipher_0_p16box_q84[15:8]}};

assign tmp_195_fu_9279_p4 = {{cipher_0_p16box_q83[15:8]}};

assign tmp_196_fu_9293_p4 = {{cipher_0_p16box_q82[15:8]}};

assign tmp_197_fu_9307_p4 = {{cipher_0_p16box_q81[15:8]}};

assign tmp_198_fu_9321_p4 = {{cipher_0_p16box_q80[15:8]}};

assign tmp_199_fu_9637_p4 = {{state_V_29_fu_9623_p2[15:8]}};

assign tmp_19_fu_4717_p4 = {{ret_V_fu_4612_p2[63:56]}};

assign tmp_200_fu_9652_p4 = {{state_V_29_fu_9623_p2[23:16]}};

assign tmp_201_fu_9667_p4 = {{state_V_29_fu_9623_p2[31:24]}};

assign tmp_202_fu_9682_p4 = {{state_V_29_fu_9623_p2[39:32]}};

assign tmp_203_fu_9697_p4 = {{state_V_29_fu_9623_p2[47:40]}};

assign tmp_204_fu_9712_p4 = {{state_V_29_fu_9623_p2[55:48]}};

assign tmp_205_fu_9727_p4 = {{state_V_29_fu_9623_p2[63:56]}};

assign tmp_206_fu_9742_p4 = {{state_V_29_fu_9623_p2[71:64]}};

assign tmp_207_fu_9757_p4 = {{state_V_29_fu_9623_p2[79:72]}};

assign tmp_208_fu_9772_p4 = {{state_V_29_fu_9623_p2[87:80]}};

assign tmp_209_fu_9787_p4 = {{state_V_29_fu_9623_p2[95:88]}};

assign tmp_20_fu_4732_p4 = {{ret_V_fu_4612_p2[71:64]}};

assign tmp_210_fu_9802_p4 = {{state_V_29_fu_9623_p2[103:96]}};

assign tmp_211_fu_9817_p4 = {{state_V_29_fu_9623_p2[111:104]}};

assign tmp_212_fu_9832_p4 = {{state_V_29_fu_9623_p2[119:112]}};

assign tmp_213_fu_9847_p4 = {{state_V_29_fu_9623_p2[127:120]}};

assign tmp_214_fu_9946_p4 = {{cipher_0_p16box_q79[15:8]}};

assign tmp_215_fu_9960_p4 = {{cipher_0_p16box_q78[15:8]}};

assign tmp_216_fu_9974_p4 = {{cipher_0_p16box_q77[15:8]}};

assign tmp_217_fu_9988_p4 = {{cipher_0_p16box_q76[15:8]}};

assign tmp_218_fu_10002_p4 = {{cipher_0_p16box_q75[15:8]}};

assign tmp_219_fu_10016_p4 = {{cipher_0_p16box_q74[15:8]}};

assign tmp_21_fu_4747_p4 = {{ret_V_fu_4612_p2[79:72]}};

assign tmp_220_fu_10030_p4 = {{cipher_0_p16box_q73[15:8]}};

assign tmp_221_fu_10044_p4 = {{cipher_0_p16box_q72[15:8]}};

assign tmp_222_fu_10058_p4 = {{cipher_0_p16box_q71[15:8]}};

assign tmp_223_fu_10072_p4 = {{cipher_0_p16box_q70[15:8]}};

assign tmp_224_fu_10086_p4 = {{cipher_0_p16box_q69[15:8]}};

assign tmp_225_fu_10100_p4 = {{cipher_0_p16box_q68[15:8]}};

assign tmp_226_fu_10114_p4 = {{cipher_0_p16box_q67[15:8]}};

assign tmp_227_fu_10128_p4 = {{cipher_0_p16box_q66[15:8]}};

assign tmp_228_fu_10142_p4 = {{cipher_0_p16box_q65[15:8]}};

assign tmp_229_fu_10156_p4 = {{cipher_0_p16box_q64[15:8]}};

assign tmp_22_fu_4762_p4 = {{ret_V_fu_4612_p2[87:80]}};

assign tmp_230_fu_10472_p4 = {{state_V_fu_10458_p2[15:8]}};

assign tmp_231_fu_10487_p4 = {{state_V_fu_10458_p2[23:16]}};

assign tmp_232_fu_10502_p4 = {{state_V_fu_10458_p2[31:24]}};

assign tmp_233_fu_10517_p4 = {{state_V_fu_10458_p2[39:32]}};

assign tmp_234_fu_10532_p4 = {{state_V_fu_10458_p2[47:40]}};

assign tmp_235_fu_10547_p4 = {{state_V_fu_10458_p2[55:48]}};

assign tmp_236_fu_10562_p4 = {{state_V_fu_10458_p2[63:56]}};

assign tmp_237_fu_10577_p4 = {{state_V_fu_10458_p2[71:64]}};

assign tmp_238_fu_10592_p4 = {{state_V_fu_10458_p2[79:72]}};

assign tmp_239_fu_10607_p4 = {{state_V_fu_10458_p2[87:80]}};

assign tmp_23_fu_4777_p4 = {{ret_V_fu_4612_p2[95:88]}};

assign tmp_240_fu_10622_p4 = {{state_V_fu_10458_p2[95:88]}};

assign tmp_241_fu_10637_p4 = {{state_V_fu_10458_p2[103:96]}};

assign tmp_242_fu_10652_p4 = {{state_V_fu_10458_p2[111:104]}};

assign tmp_243_fu_10667_p4 = {{state_V_fu_10458_p2[119:112]}};

assign tmp_244_fu_10682_p4 = {{state_V_fu_10458_p2[127:120]}};

assign tmp_245_fu_10781_p4 = {{cipher_0_p16box_q63[15:8]}};

assign tmp_246_fu_10795_p4 = {{cipher_0_p16box_q62[15:8]}};

assign tmp_247_fu_10809_p4 = {{cipher_0_p16box_q61[15:8]}};

assign tmp_248_fu_10823_p4 = {{cipher_0_p16box_q60[15:8]}};

assign tmp_249_fu_10837_p4 = {{cipher_0_p16box_q59[15:8]}};

assign tmp_24_fu_4792_p4 = {{ret_V_fu_4612_p2[103:96]}};

assign tmp_250_fu_10851_p4 = {{cipher_0_p16box_q58[15:8]}};

assign tmp_251_fu_10865_p4 = {{cipher_0_p16box_q57[15:8]}};

assign tmp_252_fu_10879_p4 = {{cipher_0_p16box_q56[15:8]}};

assign tmp_253_fu_10893_p4 = {{cipher_0_p16box_q55[15:8]}};

assign tmp_254_fu_10907_p4 = {{cipher_0_p16box_q54[15:8]}};

assign tmp_255_fu_10921_p4 = {{cipher_0_p16box_q53[15:8]}};

assign tmp_256_fu_10935_p4 = {{cipher_0_p16box_q52[15:8]}};

assign tmp_257_fu_10949_p4 = {{cipher_0_p16box_q51[15:8]}};

assign tmp_258_fu_10963_p4 = {{cipher_0_p16box_q50[15:8]}};

assign tmp_259_fu_10977_p4 = {{cipher_0_p16box_q49[15:8]}};

assign tmp_25_fu_4807_p4 = {{ret_V_fu_4612_p2[111:104]}};

assign tmp_260_fu_10991_p4 = {{cipher_0_p16box_q48[15:8]}};

assign tmp_261_fu_11307_p4 = {{state_V_30_fu_11293_p2[15:8]}};

assign tmp_262_fu_11322_p4 = {{state_V_30_fu_11293_p2[23:16]}};

assign tmp_263_fu_11337_p4 = {{state_V_30_fu_11293_p2[31:24]}};

assign tmp_264_fu_11352_p4 = {{state_V_30_fu_11293_p2[39:32]}};

assign tmp_265_fu_11367_p4 = {{state_V_30_fu_11293_p2[47:40]}};

assign tmp_266_fu_11382_p4 = {{state_V_30_fu_11293_p2[55:48]}};

assign tmp_267_fu_11397_p4 = {{state_V_30_fu_11293_p2[63:56]}};

assign tmp_268_fu_11412_p4 = {{state_V_30_fu_11293_p2[71:64]}};

assign tmp_269_fu_11427_p4 = {{state_V_30_fu_11293_p2[79:72]}};

assign tmp_26_fu_4822_p4 = {{ret_V_fu_4612_p2[119:112]}};

assign tmp_270_fu_11442_p4 = {{state_V_30_fu_11293_p2[87:80]}};

assign tmp_271_fu_11457_p4 = {{state_V_30_fu_11293_p2[95:88]}};

assign tmp_272_fu_11472_p4 = {{state_V_30_fu_11293_p2[103:96]}};

assign tmp_273_fu_11487_p4 = {{state_V_30_fu_11293_p2[111:104]}};

assign tmp_274_fu_11502_p4 = {{state_V_30_fu_11293_p2[119:112]}};

assign tmp_275_fu_11517_p4 = {{state_V_30_fu_11293_p2[127:120]}};

assign tmp_276_fu_11616_p4 = {{cipher_0_p16box_q47[15:8]}};

assign tmp_277_fu_11630_p4 = {{cipher_0_p16box_q46[15:8]}};

assign tmp_278_fu_11644_p4 = {{cipher_0_p16box_q45[15:8]}};

assign tmp_279_fu_11658_p4 = {{cipher_0_p16box_q44[15:8]}};

assign tmp_27_fu_4837_p4 = {{ret_V_fu_4612_p2[127:120]}};

assign tmp_280_fu_11672_p4 = {{cipher_0_p16box_q43[15:8]}};

assign tmp_281_fu_11686_p4 = {{cipher_0_p16box_q42[15:8]}};

assign tmp_282_fu_11700_p4 = {{cipher_0_p16box_q41[15:8]}};

assign tmp_283_fu_11714_p4 = {{cipher_0_p16box_q40[15:8]}};

assign tmp_284_fu_11728_p4 = {{cipher_0_p16box_q39[15:8]}};

assign tmp_285_fu_11742_p4 = {{cipher_0_p16box_q38[15:8]}};

assign tmp_286_fu_11756_p4 = {{cipher_0_p16box_q37[15:8]}};

assign tmp_287_fu_11770_p4 = {{cipher_0_p16box_q36[15:8]}};

assign tmp_288_fu_11784_p4 = {{cipher_0_p16box_q35[15:8]}};

assign tmp_289_fu_11798_p4 = {{cipher_0_p16box_q34[15:8]}};

assign tmp_28_fu_4936_p4 = {{cipher_0_p16box_q175[15:8]}};

assign tmp_290_fu_11812_p4 = {{cipher_0_p16box_q33[15:8]}};

assign tmp_291_fu_11826_p4 = {{cipher_0_p16box_q32[15:8]}};

assign tmp_292_fu_12142_p4 = {{state_V_31_fu_12128_p2[15:8]}};

assign tmp_293_fu_12157_p4 = {{state_V_31_fu_12128_p2[23:16]}};

assign tmp_294_fu_12172_p4 = {{state_V_31_fu_12128_p2[31:24]}};

assign tmp_295_fu_12187_p4 = {{state_V_31_fu_12128_p2[39:32]}};

assign tmp_296_fu_12202_p4 = {{state_V_31_fu_12128_p2[47:40]}};

assign tmp_297_fu_12217_p4 = {{state_V_31_fu_12128_p2[55:48]}};

assign tmp_298_fu_12232_p4 = {{state_V_31_fu_12128_p2[63:56]}};

assign tmp_299_fu_12247_p4 = {{state_V_31_fu_12128_p2[71:64]}};

assign tmp_29_fu_4950_p4 = {{cipher_0_p16box_q174[15:8]}};

assign tmp_300_fu_12262_p4 = {{state_V_31_fu_12128_p2[79:72]}};

assign tmp_301_fu_12277_p4 = {{state_V_31_fu_12128_p2[87:80]}};

assign tmp_302_fu_12292_p4 = {{state_V_31_fu_12128_p2[95:88]}};

assign tmp_303_fu_12307_p4 = {{state_V_31_fu_12128_p2[103:96]}};

assign tmp_304_fu_12322_p4 = {{state_V_31_fu_12128_p2[111:104]}};

assign tmp_305_fu_12337_p4 = {{state_V_31_fu_12128_p2[119:112]}};

assign tmp_306_fu_12352_p4 = {{state_V_31_fu_12128_p2[127:120]}};

assign tmp_307_fu_12451_p4 = {{cipher_0_p16box_q31[15:8]}};

assign tmp_308_fu_12465_p4 = {{cipher_0_p16box_q30[15:8]}};

assign tmp_309_fu_12479_p4 = {{cipher_0_p16box_q29[15:8]}};

assign tmp_30_fu_4964_p4 = {{cipher_0_p16box_q173[15:8]}};

assign tmp_310_fu_12493_p4 = {{cipher_0_p16box_q28[15:8]}};

assign tmp_311_fu_12507_p4 = {{cipher_0_p16box_q27[15:8]}};

assign tmp_312_fu_12521_p4 = {{cipher_0_p16box_q26[15:8]}};

assign tmp_313_fu_12535_p4 = {{cipher_0_p16box_q25[15:8]}};

assign tmp_314_fu_12549_p4 = {{cipher_0_p16box_q24[15:8]}};

assign tmp_315_fu_12563_p4 = {{cipher_0_p16box_q23[15:8]}};

assign tmp_316_fu_12577_p4 = {{cipher_0_p16box_q22[15:8]}};

assign tmp_317_fu_12591_p4 = {{cipher_0_p16box_q21[15:8]}};

assign tmp_318_fu_12605_p4 = {{cipher_0_p16box_q20[15:8]}};

assign tmp_319_fu_12619_p4 = {{cipher_0_p16box_q19[15:8]}};

assign tmp_31_fu_4978_p4 = {{cipher_0_p16box_q172[15:8]}};

assign tmp_320_fu_12633_p4 = {{cipher_0_p16box_q18[15:8]}};

assign tmp_321_fu_12647_p4 = {{cipher_0_p16box_q17[15:8]}};

assign tmp_322_fu_12661_p4 = {{cipher_0_p16box_q16[15:8]}};

assign tmp_323_fu_12977_p4 = {{state_V_32_fu_12963_p2[15:8]}};

assign tmp_324_fu_12992_p4 = {{state_V_32_fu_12963_p2[23:16]}};

assign tmp_325_fu_13007_p4 = {{state_V_32_fu_12963_p2[31:24]}};

assign tmp_326_fu_13022_p4 = {{state_V_32_fu_12963_p2[39:32]}};

assign tmp_327_fu_13037_p4 = {{state_V_32_fu_12963_p2[47:40]}};

assign tmp_328_fu_13052_p4 = {{state_V_32_fu_12963_p2[55:48]}};

assign tmp_329_fu_13067_p4 = {{state_V_32_fu_12963_p2[63:56]}};

assign tmp_32_fu_4992_p4 = {{cipher_0_p16box_q171[15:8]}};

assign tmp_330_fu_13082_p4 = {{state_V_32_fu_12963_p2[71:64]}};

assign tmp_331_fu_13097_p4 = {{state_V_32_fu_12963_p2[79:72]}};

assign tmp_332_fu_13112_p4 = {{state_V_32_fu_12963_p2[87:80]}};

assign tmp_333_fu_13127_p4 = {{state_V_32_fu_12963_p2[95:88]}};

assign tmp_334_fu_13142_p4 = {{state_V_32_fu_12963_p2[103:96]}};

assign tmp_335_fu_13157_p4 = {{state_V_32_fu_12963_p2[111:104]}};

assign tmp_336_fu_13172_p4 = {{state_V_32_fu_12963_p2[119:112]}};

assign tmp_337_fu_13187_p4 = {{state_V_32_fu_12963_p2[127:120]}};

assign tmp_338_fu_13286_p4 = {{cipher_0_p16box_q15[15:8]}};

assign tmp_339_fu_13300_p4 = {{cipher_0_p16box_q14[15:8]}};

assign tmp_33_fu_5006_p4 = {{cipher_0_p16box_q170[15:8]}};

assign tmp_340_fu_13314_p4 = {{cipher_0_p16box_q13[15:8]}};

assign tmp_341_fu_13328_p4 = {{cipher_0_p16box_q12[15:8]}};

assign tmp_342_fu_13342_p4 = {{cipher_0_p16box_q11[15:8]}};

assign tmp_343_fu_13356_p4 = {{cipher_0_p16box_q10[15:8]}};

assign tmp_344_fu_13370_p4 = {{cipher_0_p16box_q9[15:8]}};

assign tmp_345_fu_13384_p4 = {{cipher_0_p16box_q8[15:8]}};

assign tmp_346_fu_13398_p4 = {{cipher_0_p16box_q7[15:8]}};

assign tmp_347_fu_13412_p4 = {{cipher_0_p16box_q6[15:8]}};

assign tmp_348_fu_13426_p4 = {{cipher_0_p16box_q5[15:8]}};

assign tmp_349_fu_13440_p4 = {{cipher_0_p16box_q4[15:8]}};

assign tmp_34_fu_5020_p4 = {{cipher_0_p16box_q169[15:8]}};

assign tmp_350_fu_13454_p4 = {{cipher_0_p16box_q3[15:8]}};

assign tmp_351_fu_13468_p4 = {{cipher_0_p16box_q2[15:8]}};

assign tmp_352_fu_13482_p4 = {{cipher_0_p16box_q1[15:8]}};

assign tmp_353_fu_13496_p4 = {{cipher_0_p16box_q0[15:8]}};

assign tmp_354_fu_13812_p4 = {{state_V_33_fu_13798_p2[15:8]}};

assign tmp_355_fu_13827_p4 = {{state_V_33_fu_13798_p2[23:16]}};

assign tmp_356_fu_13842_p4 = {{state_V_33_fu_13798_p2[31:24]}};

assign tmp_357_fu_13857_p4 = {{state_V_33_fu_13798_p2[39:32]}};

assign tmp_358_fu_13872_p4 = {{state_V_33_fu_13798_p2[47:40]}};

assign tmp_359_fu_13887_p4 = {{state_V_33_fu_13798_p2[55:48]}};

assign tmp_35_fu_5034_p4 = {{cipher_0_p16box_q168[15:8]}};

assign tmp_360_fu_13902_p4 = {{state_V_33_fu_13798_p2[63:56]}};

assign tmp_361_fu_13917_p4 = {{state_V_33_fu_13798_p2[71:64]}};

assign tmp_362_fu_13932_p4 = {{state_V_33_fu_13798_p2[79:72]}};

assign tmp_363_fu_13947_p4 = {{state_V_33_fu_13798_p2[87:80]}};

assign tmp_364_fu_13962_p4 = {{state_V_33_fu_13798_p2[95:88]}};

assign tmp_365_fu_13977_p4 = {{state_V_33_fu_13798_p2[103:96]}};

assign tmp_366_fu_13992_p4 = {{state_V_33_fu_13798_p2[111:104]}};

assign tmp_367_fu_14007_p4 = {{state_V_33_fu_13798_p2[119:112]}};

assign tmp_368_fu_14022_p4 = {{state_V_33_fu_13798_p2[127:120]}};

assign tmp_36_fu_5048_p4 = {{cipher_0_p16box_q167[15:8]}};

assign tmp_37_fu_5062_p4 = {{cipher_0_p16box_q166[15:8]}};

assign tmp_38_fu_5076_p4 = {{cipher_0_p16box_q165[15:8]}};

assign tmp_39_fu_5090_p4 = {{cipher_0_p16box_q164[15:8]}};

assign tmp_40_fu_5104_p4 = {{cipher_0_p16box_q163[15:8]}};

assign tmp_41_fu_5118_p4 = {{cipher_0_p16box_q162[15:8]}};

assign tmp_42_fu_5132_p4 = {{cipher_0_p16box_q161[15:8]}};

assign tmp_43_fu_5146_p4 = {{cipher_0_p16box_q160[15:8]}};

assign tmp_44_fu_5462_p4 = {{state_V_24_fu_5448_p2[15:8]}};

assign tmp_45_fu_5477_p4 = {{state_V_24_fu_5448_p2[23:16]}};

assign tmp_46_fu_5492_p4 = {{state_V_24_fu_5448_p2[31:24]}};

assign tmp_47_fu_5507_p4 = {{state_V_24_fu_5448_p2[39:32]}};

assign tmp_48_fu_5522_p4 = {{state_V_24_fu_5448_p2[47:40]}};

assign tmp_49_fu_5537_p4 = {{state_V_24_fu_5448_p2[55:48]}};

assign tmp_50_fu_5552_p4 = {{state_V_24_fu_5448_p2[63:56]}};

assign tmp_51_fu_5567_p4 = {{state_V_24_fu_5448_p2[71:64]}};

assign tmp_52_fu_5582_p4 = {{state_V_24_fu_5448_p2[79:72]}};

assign tmp_53_fu_5597_p4 = {{state_V_24_fu_5448_p2[87:80]}};

assign tmp_54_fu_5612_p4 = {{state_V_24_fu_5448_p2[95:88]}};

assign tmp_55_fu_5627_p4 = {{state_V_24_fu_5448_p2[103:96]}};

assign tmp_56_fu_5642_p4 = {{state_V_24_fu_5448_p2[111:104]}};

assign tmp_57_fu_5657_p4 = {{state_V_24_fu_5448_p2[119:112]}};

assign tmp_58_fu_5672_p4 = {{state_V_24_fu_5448_p2[127:120]}};

assign tmp_59_fu_5771_p4 = {{cipher_0_p16box_q159[15:8]}};

assign tmp_60_fu_5785_p4 = {{cipher_0_p16box_q158[15:8]}};

assign tmp_61_fu_5799_p4 = {{cipher_0_p16box_q157[15:8]}};

assign tmp_62_fu_5813_p4 = {{cipher_0_p16box_q156[15:8]}};

assign tmp_63_fu_5827_p4 = {{cipher_0_p16box_q155[15:8]}};

assign tmp_64_fu_5841_p4 = {{cipher_0_p16box_q154[15:8]}};

assign tmp_65_fu_5855_p4 = {{cipher_0_p16box_q153[15:8]}};

assign tmp_66_fu_5869_p4 = {{cipher_0_p16box_q152[15:8]}};

assign tmp_67_fu_5883_p4 = {{cipher_0_p16box_q151[15:8]}};

assign tmp_68_fu_5897_p4 = {{cipher_0_p16box_q150[15:8]}};

assign tmp_69_fu_5911_p4 = {{cipher_0_p16box_q149[15:8]}};

assign tmp_70_fu_5925_p4 = {{cipher_0_p16box_q148[15:8]}};

assign tmp_71_fu_5939_p4 = {{cipher_0_p16box_q147[15:8]}};

assign tmp_72_fu_5953_p4 = {{cipher_0_p16box_q146[15:8]}};

assign tmp_73_fu_5967_p4 = {{cipher_0_p16box_q145[15:8]}};

assign tmp_74_fu_5981_p4 = {{cipher_0_p16box_q144[15:8]}};

assign tmp_75_fu_6297_p4 = {{state_V_25_fu_6283_p2[15:8]}};

assign tmp_76_fu_6312_p4 = {{state_V_25_fu_6283_p2[23:16]}};

assign tmp_77_fu_6327_p4 = {{state_V_25_fu_6283_p2[31:24]}};

assign tmp_78_fu_6342_p4 = {{state_V_25_fu_6283_p2[39:32]}};

assign tmp_79_fu_6357_p4 = {{state_V_25_fu_6283_p2[47:40]}};

assign tmp_80_fu_6372_p4 = {{state_V_25_fu_6283_p2[55:48]}};

assign tmp_81_fu_6387_p4 = {{state_V_25_fu_6283_p2[63:56]}};

assign tmp_82_fu_6402_p4 = {{state_V_25_fu_6283_p2[71:64]}};

assign tmp_83_fu_6417_p4 = {{state_V_25_fu_6283_p2[79:72]}};

assign tmp_84_fu_6432_p4 = {{state_V_25_fu_6283_p2[87:80]}};

assign tmp_85_fu_6447_p4 = {{state_V_25_fu_6283_p2[95:88]}};

assign tmp_86_fu_6462_p4 = {{state_V_25_fu_6283_p2[103:96]}};

assign tmp_87_fu_6477_p4 = {{state_V_25_fu_6283_p2[111:104]}};

assign tmp_88_fu_6492_p4 = {{state_V_25_fu_6283_p2[119:112]}};

assign tmp_89_fu_6507_p4 = {{state_V_25_fu_6283_p2[127:120]}};

assign tmp_90_fu_6606_p4 = {{cipher_0_p16box_q143[15:8]}};

assign tmp_91_fu_6620_p4 = {{cipher_0_p16box_q142[15:8]}};

assign tmp_92_fu_6634_p4 = {{cipher_0_p16box_q141[15:8]}};

assign tmp_93_fu_6648_p4 = {{cipher_0_p16box_q140[15:8]}};

assign tmp_94_fu_6662_p4 = {{cipher_0_p16box_q139[15:8]}};

assign tmp_95_fu_6676_p4 = {{cipher_0_p16box_q138[15:8]}};

assign tmp_96_fu_6690_p4 = {{cipher_0_p16box_q137[15:8]}};

assign tmp_97_fu_6704_p4 = {{cipher_0_p16box_q136[15:8]}};

assign tmp_98_fu_6718_p4 = {{cipher_0_p16box_q135[15:8]}};

assign tmp_99_fu_6732_p4 = {{cipher_0_p16box_q134[15:8]}};

assign tmp_s_fu_4627_p4 = {{ret_V_fu_4612_p2[15:8]}};

assign trunc_ln674_100_fu_9984_p1 = cipher_0_p16box_q76[7:0];

assign trunc_ln674_101_fu_9998_p1 = cipher_0_p16box_q75[7:0];

assign trunc_ln674_102_fu_10012_p1 = cipher_0_p16box_q74[7:0];

assign trunc_ln674_103_fu_10026_p1 = cipher_0_p16box_q73[7:0];

assign trunc_ln674_104_fu_10040_p1 = cipher_0_p16box_q72[7:0];

assign trunc_ln674_105_fu_10054_p1 = cipher_0_p16box_q71[7:0];

assign trunc_ln674_106_fu_10068_p1 = cipher_0_p16box_q70[7:0];

assign trunc_ln674_107_fu_10082_p1 = cipher_0_p16box_q69[7:0];

assign trunc_ln674_108_fu_10096_p1 = cipher_0_p16box_q68[7:0];

assign trunc_ln674_109_fu_10110_p1 = cipher_0_p16box_q67[7:0];

assign trunc_ln674_10_fu_5058_p1 = cipher_0_p16box_q166[7:0];

assign trunc_ln674_110_fu_10124_p1 = cipher_0_p16box_q66[7:0];

assign trunc_ln674_111_fu_10138_p1 = cipher_0_p16box_q65[7:0];

assign trunc_ln674_112_fu_10152_p1 = cipher_0_p16box_q64[7:0];

assign trunc_ln674_113_fu_10777_p1 = cipher_0_p16box_q63[7:0];

assign trunc_ln674_114_fu_10791_p1 = cipher_0_p16box_q62[7:0];

assign trunc_ln674_115_fu_10805_p1 = cipher_0_p16box_q61[7:0];

assign trunc_ln674_116_fu_10819_p1 = cipher_0_p16box_q60[7:0];

assign trunc_ln674_117_fu_10833_p1 = cipher_0_p16box_q59[7:0];

assign trunc_ln674_118_fu_10847_p1 = cipher_0_p16box_q58[7:0];

assign trunc_ln674_119_fu_10861_p1 = cipher_0_p16box_q57[7:0];

assign trunc_ln674_11_fu_5072_p1 = cipher_0_p16box_q165[7:0];

assign trunc_ln674_120_fu_10875_p1 = cipher_0_p16box_q56[7:0];

assign trunc_ln674_121_fu_10889_p1 = cipher_0_p16box_q55[7:0];

assign trunc_ln674_122_fu_10903_p1 = cipher_0_p16box_q54[7:0];

assign trunc_ln674_123_fu_10917_p1 = cipher_0_p16box_q53[7:0];

assign trunc_ln674_124_fu_10931_p1 = cipher_0_p16box_q52[7:0];

assign trunc_ln674_125_fu_10945_p1 = cipher_0_p16box_q51[7:0];

assign trunc_ln674_126_fu_10959_p1 = cipher_0_p16box_q50[7:0];

assign trunc_ln674_127_fu_10973_p1 = cipher_0_p16box_q49[7:0];

assign trunc_ln674_128_fu_10987_p1 = cipher_0_p16box_q48[7:0];

assign trunc_ln674_129_fu_11612_p1 = cipher_0_p16box_q47[7:0];

assign trunc_ln674_12_fu_5086_p1 = cipher_0_p16box_q164[7:0];

assign trunc_ln674_130_fu_11626_p1 = cipher_0_p16box_q46[7:0];

assign trunc_ln674_131_fu_11640_p1 = cipher_0_p16box_q45[7:0];

assign trunc_ln674_132_fu_11654_p1 = cipher_0_p16box_q44[7:0];

assign trunc_ln674_133_fu_11668_p1 = cipher_0_p16box_q43[7:0];

assign trunc_ln674_134_fu_11682_p1 = cipher_0_p16box_q42[7:0];

assign trunc_ln674_135_fu_11696_p1 = cipher_0_p16box_q41[7:0];

assign trunc_ln674_136_fu_11710_p1 = cipher_0_p16box_q40[7:0];

assign trunc_ln674_137_fu_11724_p1 = cipher_0_p16box_q39[7:0];

assign trunc_ln674_138_fu_11738_p1 = cipher_0_p16box_q38[7:0];

assign trunc_ln674_139_fu_11752_p1 = cipher_0_p16box_q37[7:0];

assign trunc_ln674_13_fu_5100_p1 = cipher_0_p16box_q163[7:0];

assign trunc_ln674_140_fu_11766_p1 = cipher_0_p16box_q36[7:0];

assign trunc_ln674_141_fu_11780_p1 = cipher_0_p16box_q35[7:0];

assign trunc_ln674_142_fu_11794_p1 = cipher_0_p16box_q34[7:0];

assign trunc_ln674_143_fu_11808_p1 = cipher_0_p16box_q33[7:0];

assign trunc_ln674_144_fu_11822_p1 = cipher_0_p16box_q32[7:0];

assign trunc_ln674_145_fu_12447_p1 = cipher_0_p16box_q31[7:0];

assign trunc_ln674_146_fu_12461_p1 = cipher_0_p16box_q30[7:0];

assign trunc_ln674_147_fu_12475_p1 = cipher_0_p16box_q29[7:0];

assign trunc_ln674_148_fu_12489_p1 = cipher_0_p16box_q28[7:0];

assign trunc_ln674_149_fu_12503_p1 = cipher_0_p16box_q27[7:0];

assign trunc_ln674_14_fu_5114_p1 = cipher_0_p16box_q162[7:0];

assign trunc_ln674_150_fu_12517_p1 = cipher_0_p16box_q26[7:0];

assign trunc_ln674_151_fu_12531_p1 = cipher_0_p16box_q25[7:0];

assign trunc_ln674_152_fu_12545_p1 = cipher_0_p16box_q24[7:0];

assign trunc_ln674_153_fu_12559_p1 = cipher_0_p16box_q23[7:0];

assign trunc_ln674_154_fu_12573_p1 = cipher_0_p16box_q22[7:0];

assign trunc_ln674_155_fu_12587_p1 = cipher_0_p16box_q21[7:0];

assign trunc_ln674_156_fu_12601_p1 = cipher_0_p16box_q20[7:0];

assign trunc_ln674_157_fu_12615_p1 = cipher_0_p16box_q19[7:0];

assign trunc_ln674_158_fu_12629_p1 = cipher_0_p16box_q18[7:0];

assign trunc_ln674_159_fu_12643_p1 = cipher_0_p16box_q17[7:0];

assign trunc_ln674_15_fu_5128_p1 = cipher_0_p16box_q161[7:0];

assign trunc_ln674_160_fu_12657_p1 = cipher_0_p16box_q16[7:0];

assign trunc_ln674_161_fu_13282_p1 = cipher_0_p16box_q15[7:0];

assign trunc_ln674_162_fu_13296_p1 = cipher_0_p16box_q14[7:0];

assign trunc_ln674_163_fu_13310_p1 = cipher_0_p16box_q13[7:0];

assign trunc_ln674_164_fu_13324_p1 = cipher_0_p16box_q12[7:0];

assign trunc_ln674_165_fu_13338_p1 = cipher_0_p16box_q11[7:0];

assign trunc_ln674_166_fu_13352_p1 = cipher_0_p16box_q10[7:0];

assign trunc_ln674_167_fu_13366_p1 = cipher_0_p16box_q9[7:0];

assign trunc_ln674_168_fu_13380_p1 = cipher_0_p16box_q8[7:0];

assign trunc_ln674_169_fu_13394_p1 = cipher_0_p16box_q7[7:0];

assign trunc_ln674_16_fu_5142_p1 = cipher_0_p16box_q160[7:0];

assign trunc_ln674_170_fu_13408_p1 = cipher_0_p16box_q6[7:0];

assign trunc_ln674_171_fu_13422_p1 = cipher_0_p16box_q5[7:0];

assign trunc_ln674_172_fu_13436_p1 = cipher_0_p16box_q4[7:0];

assign trunc_ln674_173_fu_13450_p1 = cipher_0_p16box_q3[7:0];

assign trunc_ln674_174_fu_13464_p1 = cipher_0_p16box_q2[7:0];

assign trunc_ln674_175_fu_13478_p1 = cipher_0_p16box_q1[7:0];

assign trunc_ln674_176_fu_13492_p1 = cipher_0_p16box_q0[7:0];

assign trunc_ln674_17_fu_5767_p1 = cipher_0_p16box_q159[7:0];

assign trunc_ln674_18_fu_5781_p1 = cipher_0_p16box_q158[7:0];

assign trunc_ln674_19_fu_5795_p1 = cipher_0_p16box_q157[7:0];

assign trunc_ln674_20_fu_5809_p1 = cipher_0_p16box_q156[7:0];

assign trunc_ln674_21_fu_5823_p1 = cipher_0_p16box_q155[7:0];

assign trunc_ln674_22_fu_5837_p1 = cipher_0_p16box_q154[7:0];

assign trunc_ln674_23_fu_5851_p1 = cipher_0_p16box_q153[7:0];

assign trunc_ln674_24_fu_5865_p1 = cipher_0_p16box_q152[7:0];

assign trunc_ln674_25_fu_5879_p1 = cipher_0_p16box_q151[7:0];

assign trunc_ln674_26_fu_5893_p1 = cipher_0_p16box_q150[7:0];

assign trunc_ln674_27_fu_5907_p1 = cipher_0_p16box_q149[7:0];

assign trunc_ln674_28_fu_5921_p1 = cipher_0_p16box_q148[7:0];

assign trunc_ln674_29_fu_5935_p1 = cipher_0_p16box_q147[7:0];

assign trunc_ln674_2_fu_4946_p1 = cipher_0_p16box_q174[7:0];

assign trunc_ln674_30_fu_5949_p1 = cipher_0_p16box_q146[7:0];

assign trunc_ln674_31_fu_5963_p1 = cipher_0_p16box_q145[7:0];

assign trunc_ln674_32_fu_5977_p1 = cipher_0_p16box_q144[7:0];

assign trunc_ln674_33_fu_6602_p1 = cipher_0_p16box_q143[7:0];

assign trunc_ln674_34_fu_6616_p1 = cipher_0_p16box_q142[7:0];

assign trunc_ln674_35_fu_6630_p1 = cipher_0_p16box_q141[7:0];

assign trunc_ln674_36_fu_6644_p1 = cipher_0_p16box_q140[7:0];

assign trunc_ln674_37_fu_6658_p1 = cipher_0_p16box_q139[7:0];

assign trunc_ln674_38_fu_6672_p1 = cipher_0_p16box_q138[7:0];

assign trunc_ln674_39_fu_6686_p1 = cipher_0_p16box_q137[7:0];

assign trunc_ln674_3_fu_4960_p1 = cipher_0_p16box_q173[7:0];

assign trunc_ln674_40_fu_6700_p1 = cipher_0_p16box_q136[7:0];

assign trunc_ln674_41_fu_6714_p1 = cipher_0_p16box_q135[7:0];

assign trunc_ln674_42_fu_6728_p1 = cipher_0_p16box_q134[7:0];

assign trunc_ln674_43_fu_6742_p1 = cipher_0_p16box_q133[7:0];

assign trunc_ln674_44_fu_6756_p1 = cipher_0_p16box_q132[7:0];

assign trunc_ln674_45_fu_6770_p1 = cipher_0_p16box_q131[7:0];

assign trunc_ln674_46_fu_6784_p1 = cipher_0_p16box_q130[7:0];

assign trunc_ln674_47_fu_6798_p1 = cipher_0_p16box_q129[7:0];

assign trunc_ln674_48_fu_6812_p1 = cipher_0_p16box_q128[7:0];

assign trunc_ln674_49_fu_7437_p1 = cipher_0_p16box_q127[7:0];

assign trunc_ln674_4_fu_4974_p1 = cipher_0_p16box_q172[7:0];

assign trunc_ln674_50_fu_7451_p1 = cipher_0_p16box_q126[7:0];

assign trunc_ln674_51_fu_7465_p1 = cipher_0_p16box_q125[7:0];

assign trunc_ln674_52_fu_7479_p1 = cipher_0_p16box_q124[7:0];

assign trunc_ln674_53_fu_7493_p1 = cipher_0_p16box_q123[7:0];

assign trunc_ln674_54_fu_7507_p1 = cipher_0_p16box_q122[7:0];

assign trunc_ln674_55_fu_7521_p1 = cipher_0_p16box_q121[7:0];

assign trunc_ln674_56_fu_7535_p1 = cipher_0_p16box_q120[7:0];

assign trunc_ln674_57_fu_7549_p1 = cipher_0_p16box_q119[7:0];

assign trunc_ln674_58_fu_7563_p1 = cipher_0_p16box_q118[7:0];

assign trunc_ln674_59_fu_7577_p1 = cipher_0_p16box_q117[7:0];

assign trunc_ln674_5_fu_4988_p1 = cipher_0_p16box_q171[7:0];

assign trunc_ln674_60_fu_7591_p1 = cipher_0_p16box_q116[7:0];

assign trunc_ln674_61_fu_7605_p1 = cipher_0_p16box_q115[7:0];

assign trunc_ln674_62_fu_7619_p1 = cipher_0_p16box_q114[7:0];

assign trunc_ln674_63_fu_7633_p1 = cipher_0_p16box_q113[7:0];

assign trunc_ln674_64_fu_7647_p1 = cipher_0_p16box_q112[7:0];

assign trunc_ln674_65_fu_8272_p1 = cipher_0_p16box_q111[7:0];

assign trunc_ln674_66_fu_8286_p1 = cipher_0_p16box_q110[7:0];

assign trunc_ln674_67_fu_8300_p1 = cipher_0_p16box_q109[7:0];

assign trunc_ln674_68_fu_8314_p1 = cipher_0_p16box_q108[7:0];

assign trunc_ln674_69_fu_8328_p1 = cipher_0_p16box_q107[7:0];

assign trunc_ln674_6_fu_5002_p1 = cipher_0_p16box_q170[7:0];

assign trunc_ln674_70_fu_8342_p1 = cipher_0_p16box_q106[7:0];

assign trunc_ln674_71_fu_8356_p1 = cipher_0_p16box_q105[7:0];

assign trunc_ln674_72_fu_8370_p1 = cipher_0_p16box_q104[7:0];

assign trunc_ln674_73_fu_8384_p1 = cipher_0_p16box_q103[7:0];

assign trunc_ln674_74_fu_8398_p1 = cipher_0_p16box_q102[7:0];

assign trunc_ln674_75_fu_8412_p1 = cipher_0_p16box_q101[7:0];

assign trunc_ln674_76_fu_8426_p1 = cipher_0_p16box_q100[7:0];

assign trunc_ln674_77_fu_8440_p1 = cipher_0_p16box_q99[7:0];

assign trunc_ln674_78_fu_8454_p1 = cipher_0_p16box_q98[7:0];

assign trunc_ln674_79_fu_8468_p1 = cipher_0_p16box_q97[7:0];

assign trunc_ln674_7_fu_5016_p1 = cipher_0_p16box_q169[7:0];

assign trunc_ln674_80_fu_8482_p1 = cipher_0_p16box_q96[7:0];

assign trunc_ln674_81_fu_9107_p1 = cipher_0_p16box_q95[7:0];

assign trunc_ln674_82_fu_9121_p1 = cipher_0_p16box_q94[7:0];

assign trunc_ln674_83_fu_9135_p1 = cipher_0_p16box_q93[7:0];

assign trunc_ln674_84_fu_9149_p1 = cipher_0_p16box_q92[7:0];

assign trunc_ln674_85_fu_9163_p1 = cipher_0_p16box_q91[7:0];

assign trunc_ln674_86_fu_9177_p1 = cipher_0_p16box_q90[7:0];

assign trunc_ln674_87_fu_9191_p1 = cipher_0_p16box_q89[7:0];

assign trunc_ln674_88_fu_9205_p1 = cipher_0_p16box_q88[7:0];

assign trunc_ln674_89_fu_9219_p1 = cipher_0_p16box_q87[7:0];

assign trunc_ln674_8_fu_5030_p1 = cipher_0_p16box_q168[7:0];

assign trunc_ln674_90_fu_9233_p1 = cipher_0_p16box_q86[7:0];

assign trunc_ln674_91_fu_9247_p1 = cipher_0_p16box_q85[7:0];

assign trunc_ln674_92_fu_9261_p1 = cipher_0_p16box_q84[7:0];

assign trunc_ln674_93_fu_9275_p1 = cipher_0_p16box_q83[7:0];

assign trunc_ln674_94_fu_9289_p1 = cipher_0_p16box_q82[7:0];

assign trunc_ln674_95_fu_9303_p1 = cipher_0_p16box_q81[7:0];

assign trunc_ln674_96_fu_9317_p1 = cipher_0_p16box_q80[7:0];

assign trunc_ln674_97_fu_9942_p1 = cipher_0_p16box_q79[7:0];

assign trunc_ln674_98_fu_9956_p1 = cipher_0_p16box_q78[7:0];

assign trunc_ln674_99_fu_9970_p1 = cipher_0_p16box_q77[7:0];

assign trunc_ln674_9_fu_5044_p1 = cipher_0_p16box_q167[7:0];

assign trunc_ln674_fu_4932_p1 = cipher_0_p16box_q175[7:0];

assign trunc_ln708_10_fu_12968_p1 = state_V_32_fu_12963_p2[7:0];

assign trunc_ln708_11_fu_13803_p1 = state_V_33_fu_13798_p2[7:0];

assign trunc_ln708_1_fu_5453_p1 = state_V_24_fu_5448_p2[7:0];

assign trunc_ln708_2_fu_6288_p1 = state_V_25_fu_6283_p2[7:0];

assign trunc_ln708_3_fu_7123_p1 = state_V_26_fu_7118_p2[7:0];

assign trunc_ln708_4_fu_7958_p1 = state_V_27_fu_7953_p2[7:0];

assign trunc_ln708_5_fu_8793_p1 = state_V_28_fu_8788_p2[7:0];

assign trunc_ln708_6_fu_9628_p1 = state_V_29_fu_9623_p2[7:0];

assign trunc_ln708_7_fu_10463_p1 = state_V_fu_10458_p2[7:0];

assign trunc_ln708_8_fu_11298_p1 = state_V_30_fu_11293_p2[7:0];

assign trunc_ln708_9_fu_12133_p1 = state_V_31_fu_12128_p2[7:0];

assign trunc_ln708_fu_4618_p1 = ret_V_fu_4612_p2[7:0];

assign xor_ln1545_100_fu_6241_p2 = (xor_ln1545_99_fu_6231_p2 ^ xor_ln1545_101_fu_6235_p2);

assign xor_ln1545_101_fu_6235_p2 = (trunc_ln674_32_fu_5977_p1 ^ tmp_71_fu_5939_p4);

assign xor_ln1545_102_fu_6826_p2 = (tmp_V_34_reg_14790 ^ tmp_3_V_14_reg_14820);

assign xor_ln1545_103_fu_6836_p2 = (xor_ln1545_104_fu_6830_p2 ^ xor_ln1545_102_fu_6826_p2);

assign xor_ln1545_104_fu_6830_p2 = (trunc_ln674_33_fu_6602_p1 ^ tmp_91_fu_6620_p4);

assign xor_ln1545_105_fu_6842_p2 = (tmp_V_32_reg_14730 ^ tmp_3_V_14_reg_14820);

assign xor_ln1545_106_fu_6852_p2 = (xor_ln1545_107_fu_6846_p2 ^ xor_ln1545_105_fu_6842_p2);

assign xor_ln1545_107_fu_6846_p2 = (trunc_ln674_34_fu_6616_p1 ^ tmp_92_fu_6634_p4);

assign xor_ln1545_108_fu_6858_p2 = (tmp_V_33_reg_14760 ^ tmp_V_32_reg_14730);

assign xor_ln1545_109_fu_6868_p2 = (xor_ln1545_110_fu_6862_p2 ^ xor_ln1545_108_fu_6858_p2);

assign xor_ln1545_10_fu_5182_p2 = (xor_ln1545_9_fu_5172_p2 ^ xor_ln1545_11_fu_5176_p2);

assign xor_ln1545_110_fu_6862_p2 = (trunc_ln674_35_fu_6630_p1 ^ tmp_93_fu_6648_p4);

assign xor_ln1545_111_fu_6874_p2 = (tmp_V_34_reg_14790 ^ tmp_V_33_reg_14760);

assign xor_ln1545_112_fu_6884_p2 = (xor_ln1545_113_fu_6878_p2 ^ xor_ln1545_111_fu_6874_p2);

assign xor_ln1545_113_fu_6878_p2 = (trunc_ln674_36_fu_6644_p1 ^ tmp_90_fu_6606_p4);

assign xor_ln1545_114_fu_6890_p2 = (tmp_V_39_reg_14748 ^ tmp_V_38_reg_14814);

assign xor_ln1545_115_fu_6900_p2 = (xor_ln1545_116_fu_6894_p2 ^ xor_ln1545_114_fu_6890_p2);

assign xor_ln1545_116_fu_6894_p2 = (trunc_ln674_37_fu_6658_p1 ^ tmp_95_fu_6676_p4);

assign xor_ln1545_117_fu_6906_p2 = (tmp_V_39_reg_14748 ^ tmp_V_36_reg_14754);

assign xor_ln1545_118_fu_6916_p2 = (xor_ln1545_119_fu_6910_p2 ^ xor_ln1545_117_fu_6906_p2);

assign xor_ln1545_119_fu_6910_p2 = (trunc_ln674_38_fu_6672_p1 ^ tmp_96_fu_6690_p4);

assign xor_ln1545_11_fu_5176_p2 = (trunc_ln674_2_fu_4946_p1 ^ tmp_30_fu_4964_p4);

assign xor_ln1545_120_fu_6922_p2 = (tmp_V_37_reg_14784 ^ tmp_V_36_reg_14754);

assign xor_ln1545_121_fu_6932_p2 = (xor_ln1545_122_fu_6926_p2 ^ xor_ln1545_120_fu_6922_p2);

assign xor_ln1545_122_fu_6926_p2 = (trunc_ln674_39_fu_6686_p1 ^ tmp_97_fu_6704_p4);

assign xor_ln1545_123_fu_6938_p2 = (tmp_V_38_reg_14814 ^ tmp_V_37_reg_14784);

assign xor_ln1545_124_fu_6948_p2 = (xor_ln1545_125_fu_6942_p2 ^ xor_ln1545_123_fu_6938_p2);

assign xor_ln1545_125_fu_6942_p2 = (trunc_ln674_40_fu_6700_p1 ^ tmp_94_fu_6662_p4);

assign xor_ln1545_126_fu_6954_p2 = (tmp_V_43_reg_14772 ^ tmp_2_1_V_14_reg_14742);

assign xor_ln1545_127_fu_6964_p2 = (xor_ln1545_128_fu_6958_p2 ^ xor_ln1545_126_fu_6954_p2);

assign xor_ln1545_128_fu_6958_p2 = (trunc_ln674_41_fu_6714_p1 ^ tmp_99_fu_6732_p4);

assign xor_ln1545_129_fu_6970_p2 = (tmp_V_43_reg_14772 ^ tmp_V_40_reg_14778);

assign xor_ln1545_12_fu_5188_p2 = (tmp_V_reg_14218 ^ tmp_V_1_reg_14248);

assign xor_ln1545_130_fu_6980_p2 = (xor_ln1545_131_fu_6974_p2 ^ xor_ln1545_129_fu_6970_p2);

assign xor_ln1545_131_fu_6974_p2 = (trunc_ln674_42_fu_6728_p1 ^ tmp_100_fu_6746_p4);

assign xor_ln1545_132_fu_6986_p2 = (tmp_V_41_reg_14808 ^ tmp_V_40_reg_14778);

assign xor_ln1545_133_fu_6996_p2 = (xor_ln1545_134_fu_6990_p2 ^ xor_ln1545_132_fu_6986_p2);

assign xor_ln1545_134_fu_6990_p2 = (trunc_ln674_43_fu_6742_p1 ^ tmp_101_fu_6760_p4);

assign xor_ln1545_135_fu_7002_p2 = (tmp_V_41_reg_14808 ^ tmp_2_1_V_14_reg_14742);

assign xor_ln1545_136_fu_7012_p2 = (xor_ln1545_137_fu_7006_p2 ^ xor_ln1545_135_fu_7002_p2);

assign xor_ln1545_137_fu_7006_p2 = (trunc_ln674_44_fu_6756_p1 ^ tmp_98_fu_6718_p4);

assign xor_ln1545_138_fu_7018_p2 = (tmp_V_47_reg_14796 ^ tmp_2_2_V_14_reg_14766);

assign xor_ln1545_139_fu_7028_p2 = (xor_ln1545_140_fu_7022_p2 ^ xor_ln1545_138_fu_7018_p2);

assign xor_ln1545_13_fu_5198_p2 = (xor_ln1545_14_fu_5192_p2 ^ xor_ln1545_12_fu_5188_p2);

assign xor_ln1545_140_fu_7022_p2 = (trunc_ln674_45_fu_6770_p1 ^ tmp_103_fu_6788_p4);

assign xor_ln1545_141_fu_7034_p2 = (tmp_V_47_reg_14796 ^ tmp_V_44_reg_14802);

assign xor_ln1545_142_fu_7044_p2 = (xor_ln1545_143_fu_7038_p2 ^ xor_ln1545_141_fu_7034_p2);

assign xor_ln1545_143_fu_7038_p2 = (trunc_ln674_46_fu_6784_p1 ^ tmp_104_fu_6802_p4);

assign xor_ln1545_144_fu_7050_p2 = (tmp_V_44_reg_14802 ^ tmp_1_V_14_reg_14736);

assign xor_ln1545_145_fu_7060_p2 = (xor_ln1545_146_fu_7054_p2 ^ xor_ln1545_144_fu_7050_p2);

assign xor_ln1545_146_fu_7054_p2 = (trunc_ln674_47_fu_6798_p1 ^ tmp_105_fu_6816_p4);

assign xor_ln1545_147_fu_7066_p2 = (tmp_2_2_V_14_reg_14766 ^ tmp_1_V_14_reg_14736);

assign xor_ln1545_148_fu_7076_p2 = (xor_ln1545_149_fu_7070_p2 ^ xor_ln1545_147_fu_7066_p2);

assign xor_ln1545_149_fu_7070_p2 = (trunc_ln674_48_fu_6812_p1 ^ tmp_102_fu_6774_p4);

assign xor_ln1545_14_fu_5192_p2 = (trunc_ln674_3_fu_4960_p1 ^ tmp_31_fu_4978_p4);

assign xor_ln1545_150_fu_7661_p2 = (tmp_V_50_reg_15046 ^ tmp_3_V_15_reg_15076);

assign xor_ln1545_151_fu_7671_p2 = (xor_ln1545_152_fu_7665_p2 ^ xor_ln1545_150_fu_7661_p2);

assign xor_ln1545_152_fu_7665_p2 = (trunc_ln674_49_fu_7437_p1 ^ tmp_122_fu_7455_p4);

assign xor_ln1545_153_fu_7677_p2 = (tmp_V_48_reg_14986 ^ tmp_3_V_15_reg_15076);

assign xor_ln1545_154_fu_7687_p2 = (xor_ln1545_155_fu_7681_p2 ^ xor_ln1545_153_fu_7677_p2);

assign xor_ln1545_155_fu_7681_p2 = (trunc_ln674_50_fu_7451_p1 ^ tmp_123_fu_7469_p4);

assign xor_ln1545_156_fu_7693_p2 = (tmp_V_49_reg_15016 ^ tmp_V_48_reg_14986);

assign xor_ln1545_157_fu_7703_p2 = (xor_ln1545_158_fu_7697_p2 ^ xor_ln1545_156_fu_7693_p2);

assign xor_ln1545_158_fu_7697_p2 = (trunc_ln674_51_fu_7465_p1 ^ tmp_124_fu_7483_p4);

assign xor_ln1545_159_fu_7709_p2 = (tmp_V_50_reg_15046 ^ tmp_V_49_reg_15016);

assign xor_ln1545_15_fu_5204_p2 = (tmp_V_2_reg_14278 ^ tmp_V_1_reg_14248);

assign xor_ln1545_160_fu_7719_p2 = (xor_ln1545_161_fu_7713_p2 ^ xor_ln1545_159_fu_7709_p2);

assign xor_ln1545_161_fu_7713_p2 = (trunc_ln674_52_fu_7479_p1 ^ tmp_121_fu_7441_p4);

assign xor_ln1545_162_fu_7725_p2 = (tmp_V_55_reg_15004 ^ tmp_V_54_reg_15070);

assign xor_ln1545_163_fu_7735_p2 = (xor_ln1545_164_fu_7729_p2 ^ xor_ln1545_162_fu_7725_p2);

assign xor_ln1545_164_fu_7729_p2 = (trunc_ln674_53_fu_7493_p1 ^ tmp_126_fu_7511_p4);

assign xor_ln1545_165_fu_7741_p2 = (tmp_V_55_reg_15004 ^ tmp_V_52_reg_15010);

assign xor_ln1545_166_fu_7751_p2 = (xor_ln1545_167_fu_7745_p2 ^ xor_ln1545_165_fu_7741_p2);

assign xor_ln1545_167_fu_7745_p2 = (trunc_ln674_54_fu_7507_p1 ^ tmp_127_fu_7525_p4);

assign xor_ln1545_168_fu_7757_p2 = (tmp_V_53_reg_15040 ^ tmp_V_52_reg_15010);

assign xor_ln1545_169_fu_7767_p2 = (xor_ln1545_170_fu_7761_p2 ^ xor_ln1545_168_fu_7757_p2);

assign xor_ln1545_16_fu_5214_p2 = (xor_ln1545_17_fu_5208_p2 ^ xor_ln1545_15_fu_5204_p2);

assign xor_ln1545_170_fu_7761_p2 = (trunc_ln674_55_fu_7521_p1 ^ tmp_128_fu_7539_p4);

assign xor_ln1545_171_fu_7773_p2 = (tmp_V_54_reg_15070 ^ tmp_V_53_reg_15040);

assign xor_ln1545_172_fu_7783_p2 = (xor_ln1545_173_fu_7777_p2 ^ xor_ln1545_171_fu_7773_p2);

assign xor_ln1545_173_fu_7777_p2 = (trunc_ln674_56_fu_7535_p1 ^ tmp_125_fu_7497_p4);

assign xor_ln1545_174_fu_7789_p2 = (tmp_V_59_reg_15028 ^ tmp_2_1_V_15_reg_14998);

assign xor_ln1545_175_fu_7799_p2 = (xor_ln1545_176_fu_7793_p2 ^ xor_ln1545_174_fu_7789_p2);

assign xor_ln1545_176_fu_7793_p2 = (trunc_ln674_57_fu_7549_p1 ^ tmp_130_fu_7567_p4);

assign xor_ln1545_177_fu_7805_p2 = (tmp_V_59_reg_15028 ^ tmp_V_56_reg_15034);

assign xor_ln1545_178_fu_7815_p2 = (xor_ln1545_179_fu_7809_p2 ^ xor_ln1545_177_fu_7805_p2);

assign xor_ln1545_179_fu_7809_p2 = (trunc_ln674_58_fu_7563_p1 ^ tmp_131_fu_7581_p4);

assign xor_ln1545_17_fu_5208_p2 = (trunc_ln674_4_fu_4974_p1 ^ tmp_28_fu_4936_p4);

assign xor_ln1545_180_fu_7821_p2 = (tmp_V_57_reg_15064 ^ tmp_V_56_reg_15034);

assign xor_ln1545_181_fu_7831_p2 = (xor_ln1545_182_fu_7825_p2 ^ xor_ln1545_180_fu_7821_p2);

assign xor_ln1545_182_fu_7825_p2 = (trunc_ln674_59_fu_7577_p1 ^ tmp_132_fu_7595_p4);

assign xor_ln1545_183_fu_7837_p2 = (tmp_V_57_reg_15064 ^ tmp_2_1_V_15_reg_14998);

assign xor_ln1545_184_fu_7847_p2 = (xor_ln1545_185_fu_7841_p2 ^ xor_ln1545_183_fu_7837_p2);

assign xor_ln1545_185_fu_7841_p2 = (trunc_ln674_60_fu_7591_p1 ^ tmp_129_fu_7553_p4);

assign xor_ln1545_186_fu_7853_p2 = (tmp_V_63_reg_15052 ^ tmp_2_2_V_15_reg_15022);

assign xor_ln1545_187_fu_7863_p2 = (xor_ln1545_188_fu_7857_p2 ^ xor_ln1545_186_fu_7853_p2);

assign xor_ln1545_188_fu_7857_p2 = (trunc_ln674_61_fu_7605_p1 ^ tmp_134_fu_7623_p4);

assign xor_ln1545_189_fu_7869_p2 = (tmp_V_63_reg_15052 ^ tmp_V_60_reg_15058);

assign xor_ln1545_18_fu_5220_p2 = (tmp_V_7_reg_14236 ^ tmp_V_6_reg_14302);

assign xor_ln1545_190_fu_7879_p2 = (xor_ln1545_191_fu_7873_p2 ^ xor_ln1545_189_fu_7869_p2);

assign xor_ln1545_191_fu_7873_p2 = (trunc_ln674_62_fu_7619_p1 ^ tmp_135_fu_7637_p4);

assign xor_ln1545_192_fu_7885_p2 = (tmp_V_60_reg_15058 ^ tmp_1_V_15_reg_14992);

assign xor_ln1545_193_fu_7895_p2 = (xor_ln1545_194_fu_7889_p2 ^ xor_ln1545_192_fu_7885_p2);

assign xor_ln1545_194_fu_7889_p2 = (trunc_ln674_63_fu_7633_p1 ^ tmp_136_fu_7651_p4);

assign xor_ln1545_195_fu_7901_p2 = (tmp_2_2_V_15_reg_15022 ^ tmp_1_V_15_reg_14992);

assign xor_ln1545_196_fu_7911_p2 = (xor_ln1545_197_fu_7905_p2 ^ xor_ln1545_195_fu_7901_p2);

assign xor_ln1545_197_fu_7905_p2 = (trunc_ln674_64_fu_7647_p1 ^ tmp_133_fu_7609_p4);

assign xor_ln1545_198_fu_8496_p2 = (tmp_V_66_reg_15302 ^ tmp_3_V_16_reg_15332);

assign xor_ln1545_199_fu_8506_p2 = (xor_ln1545_200_fu_8500_p2 ^ xor_ln1545_198_fu_8496_p2);

assign xor_ln1545_19_fu_5230_p2 = (xor_ln1545_20_fu_5224_p2 ^ xor_ln1545_18_fu_5220_p2);

assign xor_ln1545_200_fu_8500_p2 = (trunc_ln674_65_fu_8272_p1 ^ tmp_153_fu_8290_p4);

assign xor_ln1545_201_fu_8512_p2 = (tmp_V_64_reg_15242 ^ tmp_3_V_16_reg_15332);

assign xor_ln1545_202_fu_8522_p2 = (xor_ln1545_203_fu_8516_p2 ^ xor_ln1545_201_fu_8512_p2);

assign xor_ln1545_203_fu_8516_p2 = (trunc_ln674_66_fu_8286_p1 ^ tmp_154_fu_8304_p4);

assign xor_ln1545_204_fu_8528_p2 = (tmp_V_65_reg_15272 ^ tmp_V_64_reg_15242);

assign xor_ln1545_205_fu_8538_p2 = (xor_ln1545_206_fu_8532_p2 ^ xor_ln1545_204_fu_8528_p2);

assign xor_ln1545_206_fu_8532_p2 = (trunc_ln674_67_fu_8300_p1 ^ tmp_155_fu_8318_p4);

assign xor_ln1545_207_fu_8544_p2 = (tmp_V_66_reg_15302 ^ tmp_V_65_reg_15272);

assign xor_ln1545_208_fu_8554_p2 = (xor_ln1545_209_fu_8548_p2 ^ xor_ln1545_207_fu_8544_p2);

assign xor_ln1545_209_fu_8548_p2 = (trunc_ln674_68_fu_8314_p1 ^ tmp_152_fu_8276_p4);

assign xor_ln1545_20_fu_5224_p2 = (trunc_ln674_5_fu_4988_p1 ^ tmp_33_fu_5006_p4);

assign xor_ln1545_210_fu_8560_p2 = (tmp_V_71_reg_15260 ^ tmp_V_70_reg_15326);

assign xor_ln1545_211_fu_8570_p2 = (xor_ln1545_212_fu_8564_p2 ^ xor_ln1545_210_fu_8560_p2);

assign xor_ln1545_212_fu_8564_p2 = (trunc_ln674_69_fu_8328_p1 ^ tmp_157_fu_8346_p4);

assign xor_ln1545_213_fu_8576_p2 = (tmp_V_71_reg_15260 ^ tmp_V_68_reg_15266);

assign xor_ln1545_214_fu_8586_p2 = (xor_ln1545_215_fu_8580_p2 ^ xor_ln1545_213_fu_8576_p2);

assign xor_ln1545_215_fu_8580_p2 = (trunc_ln674_70_fu_8342_p1 ^ tmp_158_fu_8360_p4);

assign xor_ln1545_216_fu_8592_p2 = (tmp_V_69_reg_15296 ^ tmp_V_68_reg_15266);

assign xor_ln1545_217_fu_8602_p2 = (xor_ln1545_218_fu_8596_p2 ^ xor_ln1545_216_fu_8592_p2);

assign xor_ln1545_218_fu_8596_p2 = (trunc_ln674_71_fu_8356_p1 ^ tmp_159_fu_8374_p4);

assign xor_ln1545_219_fu_8608_p2 = (tmp_V_70_reg_15326 ^ tmp_V_69_reg_15296);

assign xor_ln1545_21_fu_5236_p2 = (tmp_V_7_reg_14236 ^ tmp_V_4_reg_14242);

assign xor_ln1545_220_fu_8618_p2 = (xor_ln1545_221_fu_8612_p2 ^ xor_ln1545_219_fu_8608_p2);

assign xor_ln1545_221_fu_8612_p2 = (trunc_ln674_72_fu_8370_p1 ^ tmp_156_fu_8332_p4);

assign xor_ln1545_222_fu_8624_p2 = (tmp_V_75_reg_15284 ^ tmp_2_1_V_16_reg_15254);

assign xor_ln1545_223_fu_8634_p2 = (xor_ln1545_224_fu_8628_p2 ^ xor_ln1545_222_fu_8624_p2);

assign xor_ln1545_224_fu_8628_p2 = (trunc_ln674_73_fu_8384_p1 ^ tmp_161_fu_8402_p4);

assign xor_ln1545_225_fu_8640_p2 = (tmp_V_75_reg_15284 ^ tmp_V_72_reg_15290);

assign xor_ln1545_226_fu_8650_p2 = (xor_ln1545_227_fu_8644_p2 ^ xor_ln1545_225_fu_8640_p2);

assign xor_ln1545_227_fu_8644_p2 = (trunc_ln674_74_fu_8398_p1 ^ tmp_162_fu_8416_p4);

assign xor_ln1545_228_fu_8656_p2 = (tmp_V_73_reg_15320 ^ tmp_V_72_reg_15290);

assign xor_ln1545_229_fu_8666_p2 = (xor_ln1545_230_fu_8660_p2 ^ xor_ln1545_228_fu_8656_p2);

assign xor_ln1545_22_fu_5246_p2 = (xor_ln1545_23_fu_5240_p2 ^ xor_ln1545_21_fu_5236_p2);

assign xor_ln1545_230_fu_8660_p2 = (trunc_ln674_75_fu_8412_p1 ^ tmp_163_fu_8430_p4);

assign xor_ln1545_231_fu_8672_p2 = (tmp_V_73_reg_15320 ^ tmp_2_1_V_16_reg_15254);

assign xor_ln1545_232_fu_8682_p2 = (xor_ln1545_233_fu_8676_p2 ^ xor_ln1545_231_fu_8672_p2);

assign xor_ln1545_233_fu_8676_p2 = (trunc_ln674_76_fu_8426_p1 ^ tmp_160_fu_8388_p4);

assign xor_ln1545_234_fu_8688_p2 = (tmp_V_79_reg_15308 ^ tmp_2_2_V_16_reg_15278);

assign xor_ln1545_235_fu_8698_p2 = (xor_ln1545_236_fu_8692_p2 ^ xor_ln1545_234_fu_8688_p2);

assign xor_ln1545_236_fu_8692_p2 = (trunc_ln674_77_fu_8440_p1 ^ tmp_165_fu_8458_p4);

assign xor_ln1545_237_fu_8704_p2 = (tmp_V_79_reg_15308 ^ tmp_V_76_reg_15314);

assign xor_ln1545_238_fu_8714_p2 = (xor_ln1545_239_fu_8708_p2 ^ xor_ln1545_237_fu_8704_p2);

assign xor_ln1545_239_fu_8708_p2 = (trunc_ln674_78_fu_8454_p1 ^ tmp_166_fu_8472_p4);

assign xor_ln1545_23_fu_5240_p2 = (trunc_ln674_6_fu_5002_p1 ^ tmp_34_fu_5020_p4);

assign xor_ln1545_240_fu_8720_p2 = (tmp_V_76_reg_15314 ^ tmp_1_V_16_reg_15248);

assign xor_ln1545_241_fu_8730_p2 = (xor_ln1545_242_fu_8724_p2 ^ xor_ln1545_240_fu_8720_p2);

assign xor_ln1545_242_fu_8724_p2 = (trunc_ln674_79_fu_8468_p1 ^ tmp_167_fu_8486_p4);

assign xor_ln1545_243_fu_8736_p2 = (tmp_2_2_V_16_reg_15278 ^ tmp_1_V_16_reg_15248);

assign xor_ln1545_244_fu_8746_p2 = (xor_ln1545_245_fu_8740_p2 ^ xor_ln1545_243_fu_8736_p2);

assign xor_ln1545_245_fu_8740_p2 = (trunc_ln674_80_fu_8482_p1 ^ tmp_164_fu_8444_p4);

assign xor_ln1545_246_fu_9331_p2 = (tmp_V_82_reg_15558 ^ tmp_3_V_17_reg_15588);

assign xor_ln1545_247_fu_9341_p2 = (xor_ln1545_248_fu_9335_p2 ^ xor_ln1545_246_fu_9331_p2);

assign xor_ln1545_248_fu_9335_p2 = (trunc_ln674_81_fu_9107_p1 ^ tmp_184_fu_9125_p4);

assign xor_ln1545_249_fu_9347_p2 = (tmp_V_80_reg_15498 ^ tmp_3_V_17_reg_15588);

assign xor_ln1545_24_fu_5252_p2 = (tmp_V_5_reg_14272 ^ tmp_V_4_reg_14242);

assign xor_ln1545_250_fu_9357_p2 = (xor_ln1545_251_fu_9351_p2 ^ xor_ln1545_249_fu_9347_p2);

assign xor_ln1545_251_fu_9351_p2 = (trunc_ln674_82_fu_9121_p1 ^ tmp_185_fu_9139_p4);

assign xor_ln1545_252_fu_9363_p2 = (tmp_V_81_reg_15528 ^ tmp_V_80_reg_15498);

assign xor_ln1545_253_fu_9373_p2 = (xor_ln1545_254_fu_9367_p2 ^ xor_ln1545_252_fu_9363_p2);

assign xor_ln1545_254_fu_9367_p2 = (trunc_ln674_83_fu_9135_p1 ^ tmp_186_fu_9153_p4);

assign xor_ln1545_255_fu_9379_p2 = (tmp_V_82_reg_15558 ^ tmp_V_81_reg_15528);

assign xor_ln1545_256_fu_9389_p2 = (xor_ln1545_257_fu_9383_p2 ^ xor_ln1545_255_fu_9379_p2);

assign xor_ln1545_257_fu_9383_p2 = (trunc_ln674_84_fu_9149_p1 ^ tmp_183_fu_9111_p4);

assign xor_ln1545_258_fu_9395_p2 = (tmp_V_87_reg_15516 ^ tmp_V_86_reg_15582);

assign xor_ln1545_259_fu_9405_p2 = (xor_ln1545_260_fu_9399_p2 ^ xor_ln1545_258_fu_9395_p2);

assign xor_ln1545_25_fu_5262_p2 = (xor_ln1545_26_fu_5256_p2 ^ xor_ln1545_24_fu_5252_p2);

assign xor_ln1545_260_fu_9399_p2 = (trunc_ln674_85_fu_9163_p1 ^ tmp_188_fu_9181_p4);

assign xor_ln1545_261_fu_9411_p2 = (tmp_V_87_reg_15516 ^ tmp_V_84_reg_15522);

assign xor_ln1545_262_fu_9421_p2 = (xor_ln1545_263_fu_9415_p2 ^ xor_ln1545_261_fu_9411_p2);

assign xor_ln1545_263_fu_9415_p2 = (trunc_ln674_86_fu_9177_p1 ^ tmp_189_fu_9195_p4);

assign xor_ln1545_264_fu_9427_p2 = (tmp_V_85_reg_15552 ^ tmp_V_84_reg_15522);

assign xor_ln1545_265_fu_9437_p2 = (xor_ln1545_266_fu_9431_p2 ^ xor_ln1545_264_fu_9427_p2);

assign xor_ln1545_266_fu_9431_p2 = (trunc_ln674_87_fu_9191_p1 ^ tmp_190_fu_9209_p4);

assign xor_ln1545_267_fu_9443_p2 = (tmp_V_86_reg_15582 ^ tmp_V_85_reg_15552);

assign xor_ln1545_268_fu_9453_p2 = (xor_ln1545_269_fu_9447_p2 ^ xor_ln1545_267_fu_9443_p2);

assign xor_ln1545_269_fu_9447_p2 = (trunc_ln674_88_fu_9205_p1 ^ tmp_187_fu_9167_p4);

assign xor_ln1545_26_fu_5256_p2 = (trunc_ln674_7_fu_5016_p1 ^ tmp_35_fu_5034_p4);

assign xor_ln1545_270_fu_9459_p2 = (tmp_V_91_reg_15540 ^ tmp_2_1_V_17_reg_15510);

assign xor_ln1545_271_fu_9469_p2 = (xor_ln1545_272_fu_9463_p2 ^ xor_ln1545_270_fu_9459_p2);

assign xor_ln1545_272_fu_9463_p2 = (trunc_ln674_89_fu_9219_p1 ^ tmp_192_fu_9237_p4);

assign xor_ln1545_273_fu_9475_p2 = (tmp_V_91_reg_15540 ^ tmp_V_88_reg_15546);

assign xor_ln1545_274_fu_9485_p2 = (xor_ln1545_275_fu_9479_p2 ^ xor_ln1545_273_fu_9475_p2);

assign xor_ln1545_275_fu_9479_p2 = (trunc_ln674_90_fu_9233_p1 ^ tmp_193_fu_9251_p4);

assign xor_ln1545_276_fu_9491_p2 = (tmp_V_89_reg_15576 ^ tmp_V_88_reg_15546);

assign xor_ln1545_277_fu_9501_p2 = (xor_ln1545_278_fu_9495_p2 ^ xor_ln1545_276_fu_9491_p2);

assign xor_ln1545_278_fu_9495_p2 = (trunc_ln674_91_fu_9247_p1 ^ tmp_194_fu_9265_p4);

assign xor_ln1545_279_fu_9507_p2 = (tmp_V_89_reg_15576 ^ tmp_2_1_V_17_reg_15510);

assign xor_ln1545_27_fu_5268_p2 = (tmp_V_6_reg_14302 ^ tmp_V_5_reg_14272);

assign xor_ln1545_280_fu_9517_p2 = (xor_ln1545_281_fu_9511_p2 ^ xor_ln1545_279_fu_9507_p2);

assign xor_ln1545_281_fu_9511_p2 = (trunc_ln674_92_fu_9261_p1 ^ tmp_191_fu_9223_p4);

assign xor_ln1545_282_fu_9523_p2 = (tmp_V_95_reg_15564 ^ tmp_2_2_V_17_reg_15534);

assign xor_ln1545_283_fu_9533_p2 = (xor_ln1545_284_fu_9527_p2 ^ xor_ln1545_282_fu_9523_p2);

assign xor_ln1545_284_fu_9527_p2 = (trunc_ln674_93_fu_9275_p1 ^ tmp_196_fu_9293_p4);

assign xor_ln1545_285_fu_9539_p2 = (tmp_V_95_reg_15564 ^ tmp_V_92_reg_15570);

assign xor_ln1545_286_fu_9549_p2 = (xor_ln1545_287_fu_9543_p2 ^ xor_ln1545_285_fu_9539_p2);

assign xor_ln1545_287_fu_9543_p2 = (trunc_ln674_94_fu_9289_p1 ^ tmp_197_fu_9307_p4);

assign xor_ln1545_288_fu_9555_p2 = (tmp_V_92_reg_15570 ^ tmp_1_V_17_reg_15504);

assign xor_ln1545_289_fu_9565_p2 = (xor_ln1545_290_fu_9559_p2 ^ xor_ln1545_288_fu_9555_p2);

assign xor_ln1545_28_fu_5278_p2 = (xor_ln1545_29_fu_5272_p2 ^ xor_ln1545_27_fu_5268_p2);

assign xor_ln1545_290_fu_9559_p2 = (trunc_ln674_95_fu_9303_p1 ^ tmp_198_fu_9321_p4);

assign xor_ln1545_291_fu_9571_p2 = (tmp_2_2_V_17_reg_15534 ^ tmp_1_V_17_reg_15504);

assign xor_ln1545_292_fu_9581_p2 = (xor_ln1545_293_fu_9575_p2 ^ xor_ln1545_291_fu_9571_p2);

assign xor_ln1545_293_fu_9575_p2 = (trunc_ln674_96_fu_9317_p1 ^ tmp_195_fu_9279_p4);

assign xor_ln1545_294_fu_10166_p2 = (tmp_V_98_reg_15814 ^ tmp_3_V_18_reg_15844);

assign xor_ln1545_295_fu_10176_p2 = (xor_ln1545_296_fu_10170_p2 ^ xor_ln1545_294_fu_10166_p2);

assign xor_ln1545_296_fu_10170_p2 = (trunc_ln674_97_fu_9942_p1 ^ tmp_215_fu_9960_p4);

assign xor_ln1545_297_fu_10182_p2 = (tmp_V_96_reg_15754 ^ tmp_3_V_18_reg_15844);

assign xor_ln1545_298_fu_10192_p2 = (xor_ln1545_299_fu_10186_p2 ^ xor_ln1545_297_fu_10182_p2);

assign xor_ln1545_299_fu_10186_p2 = (trunc_ln674_98_fu_9956_p1 ^ tmp_216_fu_9974_p4);

assign xor_ln1545_29_fu_5272_p2 = (trunc_ln674_8_fu_5030_p1 ^ tmp_32_fu_4992_p4);

assign xor_ln1545_300_fu_10198_p2 = (tmp_V_97_reg_15784 ^ tmp_V_96_reg_15754);

assign xor_ln1545_301_fu_10208_p2 = (xor_ln1545_302_fu_10202_p2 ^ xor_ln1545_300_fu_10198_p2);

assign xor_ln1545_302_fu_10202_p2 = (trunc_ln674_99_fu_9970_p1 ^ tmp_217_fu_9988_p4);

assign xor_ln1545_303_fu_10214_p2 = (tmp_V_98_reg_15814 ^ tmp_V_97_reg_15784);

assign xor_ln1545_304_fu_10224_p2 = (xor_ln1545_305_fu_10218_p2 ^ xor_ln1545_303_fu_10214_p2);

assign xor_ln1545_305_fu_10218_p2 = (trunc_ln674_100_fu_9984_p1 ^ tmp_214_fu_9946_p4);

assign xor_ln1545_306_fu_10230_p2 = (tmp_V_103_reg_15772 ^ tmp_V_102_reg_15838);

assign xor_ln1545_307_fu_10240_p2 = (xor_ln1545_308_fu_10234_p2 ^ xor_ln1545_306_fu_10230_p2);

assign xor_ln1545_308_fu_10234_p2 = (trunc_ln674_101_fu_9998_p1 ^ tmp_219_fu_10016_p4);

assign xor_ln1545_309_fu_10246_p2 = (tmp_V_103_reg_15772 ^ tmp_V_100_reg_15778);

assign xor_ln1545_30_fu_5284_p2 = (tmp_V_11_reg_14260 ^ tmp_2_1_V_12_reg_14230);

assign xor_ln1545_310_fu_10256_p2 = (xor_ln1545_311_fu_10250_p2 ^ xor_ln1545_309_fu_10246_p2);

assign xor_ln1545_311_fu_10250_p2 = (trunc_ln674_102_fu_10012_p1 ^ tmp_220_fu_10030_p4);

assign xor_ln1545_312_fu_10262_p2 = (tmp_V_101_reg_15808 ^ tmp_V_100_reg_15778);

assign xor_ln1545_313_fu_10272_p2 = (xor_ln1545_314_fu_10266_p2 ^ xor_ln1545_312_fu_10262_p2);

assign xor_ln1545_314_fu_10266_p2 = (trunc_ln674_103_fu_10026_p1 ^ tmp_221_fu_10044_p4);

assign xor_ln1545_315_fu_10278_p2 = (tmp_V_102_reg_15838 ^ tmp_V_101_reg_15808);

assign xor_ln1545_316_fu_10288_p2 = (xor_ln1545_317_fu_10282_p2 ^ xor_ln1545_315_fu_10278_p2);

assign xor_ln1545_317_fu_10282_p2 = (trunc_ln674_104_fu_10040_p1 ^ tmp_218_fu_10002_p4);

assign xor_ln1545_318_fu_10294_p2 = (tmp_V_107_reg_15796 ^ tmp_2_1_V_18_reg_15766);

assign xor_ln1545_319_fu_10304_p2 = (xor_ln1545_320_fu_10298_p2 ^ xor_ln1545_318_fu_10294_p2);

assign xor_ln1545_31_fu_5294_p2 = (xor_ln1545_32_fu_5288_p2 ^ xor_ln1545_30_fu_5284_p2);

assign xor_ln1545_320_fu_10298_p2 = (trunc_ln674_105_fu_10054_p1 ^ tmp_223_fu_10072_p4);

assign xor_ln1545_321_fu_10310_p2 = (tmp_V_107_reg_15796 ^ tmp_V_104_reg_15802);

assign xor_ln1545_322_fu_10320_p2 = (xor_ln1545_323_fu_10314_p2 ^ xor_ln1545_321_fu_10310_p2);

assign xor_ln1545_323_fu_10314_p2 = (trunc_ln674_106_fu_10068_p1 ^ tmp_224_fu_10086_p4);

assign xor_ln1545_324_fu_10326_p2 = (tmp_V_105_reg_15832 ^ tmp_V_104_reg_15802);

assign xor_ln1545_325_fu_10336_p2 = (xor_ln1545_326_fu_10330_p2 ^ xor_ln1545_324_fu_10326_p2);

assign xor_ln1545_326_fu_10330_p2 = (trunc_ln674_107_fu_10082_p1 ^ tmp_225_fu_10100_p4);

assign xor_ln1545_327_fu_10342_p2 = (tmp_V_105_reg_15832 ^ tmp_2_1_V_18_reg_15766);

assign xor_ln1545_328_fu_10352_p2 = (xor_ln1545_329_fu_10346_p2 ^ xor_ln1545_327_fu_10342_p2);

assign xor_ln1545_329_fu_10346_p2 = (trunc_ln674_108_fu_10096_p1 ^ tmp_222_fu_10058_p4);

assign xor_ln1545_32_fu_5288_p2 = (trunc_ln674_9_fu_5044_p1 ^ tmp_37_fu_5062_p4);

assign xor_ln1545_330_fu_10358_p2 = (tmp_V_111_reg_15820 ^ tmp_2_2_V_18_reg_15790);

assign xor_ln1545_331_fu_10368_p2 = (xor_ln1545_332_fu_10362_p2 ^ xor_ln1545_330_fu_10358_p2);

assign xor_ln1545_332_fu_10362_p2 = (trunc_ln674_109_fu_10110_p1 ^ tmp_227_fu_10128_p4);

assign xor_ln1545_333_fu_10374_p2 = (tmp_V_111_reg_15820 ^ tmp_V_108_reg_15826);

assign xor_ln1545_334_fu_10384_p2 = (xor_ln1545_335_fu_10378_p2 ^ xor_ln1545_333_fu_10374_p2);

assign xor_ln1545_335_fu_10378_p2 = (trunc_ln674_110_fu_10124_p1 ^ tmp_228_fu_10142_p4);

assign xor_ln1545_336_fu_10390_p2 = (tmp_V_108_reg_15826 ^ tmp_1_V_18_reg_15760);

assign xor_ln1545_337_fu_10400_p2 = (xor_ln1545_338_fu_10394_p2 ^ xor_ln1545_336_fu_10390_p2);

assign xor_ln1545_338_fu_10394_p2 = (trunc_ln674_111_fu_10138_p1 ^ tmp_229_fu_10156_p4);

assign xor_ln1545_339_fu_10406_p2 = (tmp_2_2_V_18_reg_15790 ^ tmp_1_V_18_reg_15760);

assign xor_ln1545_33_fu_5300_p2 = (tmp_V_8_reg_14266 ^ tmp_V_11_reg_14260);

assign xor_ln1545_340_fu_10416_p2 = (xor_ln1545_341_fu_10410_p2 ^ xor_ln1545_339_fu_10406_p2);

assign xor_ln1545_341_fu_10410_p2 = (trunc_ln674_112_fu_10152_p1 ^ tmp_226_fu_10114_p4);

assign xor_ln1545_342_fu_11001_p2 = (tmp_V_114_reg_16070 ^ tmp_3_V_19_reg_16100);

assign xor_ln1545_343_fu_11011_p2 = (xor_ln1545_344_fu_11005_p2 ^ xor_ln1545_342_fu_11001_p2);

assign xor_ln1545_344_fu_11005_p2 = (trunc_ln674_113_fu_10777_p1 ^ tmp_246_fu_10795_p4);

assign xor_ln1545_345_fu_11017_p2 = (tmp_V_112_reg_16010 ^ tmp_3_V_19_reg_16100);

assign xor_ln1545_346_fu_11027_p2 = (xor_ln1545_347_fu_11021_p2 ^ xor_ln1545_345_fu_11017_p2);

assign xor_ln1545_347_fu_11021_p2 = (trunc_ln674_114_fu_10791_p1 ^ tmp_247_fu_10809_p4);

assign xor_ln1545_348_fu_11033_p2 = (tmp_V_113_reg_16040 ^ tmp_V_112_reg_16010);

assign xor_ln1545_349_fu_11043_p2 = (xor_ln1545_350_fu_11037_p2 ^ xor_ln1545_348_fu_11033_p2);

assign xor_ln1545_34_fu_5310_p2 = (xor_ln1545_35_fu_5304_p2 ^ xor_ln1545_33_fu_5300_p2);

assign xor_ln1545_350_fu_11037_p2 = (trunc_ln674_115_fu_10805_p1 ^ tmp_248_fu_10823_p4);

assign xor_ln1545_351_fu_11049_p2 = (tmp_V_114_reg_16070 ^ tmp_V_113_reg_16040);

assign xor_ln1545_352_fu_11059_p2 = (xor_ln1545_353_fu_11053_p2 ^ xor_ln1545_351_fu_11049_p2);

assign xor_ln1545_353_fu_11053_p2 = (trunc_ln674_116_fu_10819_p1 ^ tmp_245_fu_10781_p4);

assign xor_ln1545_354_fu_11065_p2 = (tmp_V_119_reg_16028 ^ tmp_V_118_reg_16094);

assign xor_ln1545_355_fu_11075_p2 = (xor_ln1545_356_fu_11069_p2 ^ xor_ln1545_354_fu_11065_p2);

assign xor_ln1545_356_fu_11069_p2 = (trunc_ln674_117_fu_10833_p1 ^ tmp_250_fu_10851_p4);

assign xor_ln1545_357_fu_11081_p2 = (tmp_V_119_reg_16028 ^ tmp_V_116_reg_16034);

assign xor_ln1545_358_fu_11091_p2 = (xor_ln1545_359_fu_11085_p2 ^ xor_ln1545_357_fu_11081_p2);

assign xor_ln1545_359_fu_11085_p2 = (trunc_ln674_118_fu_10847_p1 ^ tmp_251_fu_10865_p4);

assign xor_ln1545_35_fu_5304_p2 = (trunc_ln674_10_fu_5058_p1 ^ tmp_38_fu_5076_p4);

assign xor_ln1545_360_fu_11097_p2 = (tmp_V_117_reg_16064 ^ tmp_V_116_reg_16034);

assign xor_ln1545_361_fu_11107_p2 = (xor_ln1545_362_fu_11101_p2 ^ xor_ln1545_360_fu_11097_p2);

assign xor_ln1545_362_fu_11101_p2 = (trunc_ln674_119_fu_10861_p1 ^ tmp_252_fu_10879_p4);

assign xor_ln1545_363_fu_11113_p2 = (tmp_V_118_reg_16094 ^ tmp_V_117_reg_16064);

assign xor_ln1545_364_fu_11123_p2 = (xor_ln1545_365_fu_11117_p2 ^ xor_ln1545_363_fu_11113_p2);

assign xor_ln1545_365_fu_11117_p2 = (trunc_ln674_120_fu_10875_p1 ^ tmp_249_fu_10837_p4);

assign xor_ln1545_366_fu_11129_p2 = (tmp_V_123_reg_16052 ^ tmp_2_1_V_19_reg_16022);

assign xor_ln1545_367_fu_11139_p2 = (xor_ln1545_368_fu_11133_p2 ^ xor_ln1545_366_fu_11129_p2);

assign xor_ln1545_368_fu_11133_p2 = (trunc_ln674_121_fu_10889_p1 ^ tmp_254_fu_10907_p4);

assign xor_ln1545_369_fu_11145_p2 = (tmp_V_123_reg_16052 ^ tmp_V_120_reg_16058);

assign xor_ln1545_36_fu_5316_p2 = (tmp_V_9_reg_14296 ^ tmp_V_8_reg_14266);

assign xor_ln1545_370_fu_11155_p2 = (xor_ln1545_371_fu_11149_p2 ^ xor_ln1545_369_fu_11145_p2);

assign xor_ln1545_371_fu_11149_p2 = (trunc_ln674_122_fu_10903_p1 ^ tmp_255_fu_10921_p4);

assign xor_ln1545_372_fu_11161_p2 = (tmp_V_121_reg_16088 ^ tmp_V_120_reg_16058);

assign xor_ln1545_373_fu_11171_p2 = (xor_ln1545_374_fu_11165_p2 ^ xor_ln1545_372_fu_11161_p2);

assign xor_ln1545_374_fu_11165_p2 = (trunc_ln674_123_fu_10917_p1 ^ tmp_256_fu_10935_p4);

assign xor_ln1545_375_fu_11177_p2 = (tmp_V_121_reg_16088 ^ tmp_2_1_V_19_reg_16022);

assign xor_ln1545_376_fu_11187_p2 = (xor_ln1545_377_fu_11181_p2 ^ xor_ln1545_375_fu_11177_p2);

assign xor_ln1545_377_fu_11181_p2 = (trunc_ln674_124_fu_10931_p1 ^ tmp_253_fu_10893_p4);

assign xor_ln1545_378_fu_11193_p2 = (tmp_V_127_reg_16076 ^ tmp_2_2_V_19_reg_16046);

assign xor_ln1545_379_fu_11203_p2 = (xor_ln1545_380_fu_11197_p2 ^ xor_ln1545_378_fu_11193_p2);

assign xor_ln1545_37_fu_5326_p2 = (xor_ln1545_38_fu_5320_p2 ^ xor_ln1545_36_fu_5316_p2);

assign xor_ln1545_380_fu_11197_p2 = (trunc_ln674_125_fu_10945_p1 ^ tmp_258_fu_10963_p4);

assign xor_ln1545_381_fu_11209_p2 = (tmp_V_127_reg_16076 ^ tmp_V_124_reg_16082);

assign xor_ln1545_382_fu_11219_p2 = (xor_ln1545_383_fu_11213_p2 ^ xor_ln1545_381_fu_11209_p2);

assign xor_ln1545_383_fu_11213_p2 = (trunc_ln674_126_fu_10959_p1 ^ tmp_259_fu_10977_p4);

assign xor_ln1545_384_fu_11225_p2 = (tmp_V_124_reg_16082 ^ tmp_1_V_19_reg_16016);

assign xor_ln1545_385_fu_11235_p2 = (xor_ln1545_386_fu_11229_p2 ^ xor_ln1545_384_fu_11225_p2);

assign xor_ln1545_386_fu_11229_p2 = (trunc_ln674_127_fu_10973_p1 ^ tmp_260_fu_10991_p4);

assign xor_ln1545_387_fu_11241_p2 = (tmp_2_2_V_19_reg_16046 ^ tmp_1_V_19_reg_16016);

assign xor_ln1545_388_fu_11251_p2 = (xor_ln1545_389_fu_11245_p2 ^ xor_ln1545_387_fu_11241_p2);

assign xor_ln1545_389_fu_11245_p2 = (trunc_ln674_128_fu_10987_p1 ^ tmp_257_fu_10949_p4);

assign xor_ln1545_38_fu_5320_p2 = (trunc_ln674_11_fu_5072_p1 ^ tmp_39_fu_5090_p4);

assign xor_ln1545_390_fu_11836_p2 = (tmp_V_130_reg_16326 ^ tmp_3_V_20_reg_16356);

assign xor_ln1545_391_fu_11846_p2 = (xor_ln1545_392_fu_11840_p2 ^ xor_ln1545_390_fu_11836_p2);

assign xor_ln1545_392_fu_11840_p2 = (trunc_ln674_129_fu_11612_p1 ^ tmp_277_fu_11630_p4);

assign xor_ln1545_393_fu_11852_p2 = (tmp_V_128_reg_16266 ^ tmp_3_V_20_reg_16356);

assign xor_ln1545_394_fu_11862_p2 = (xor_ln1545_395_fu_11856_p2 ^ xor_ln1545_393_fu_11852_p2);

assign xor_ln1545_395_fu_11856_p2 = (trunc_ln674_130_fu_11626_p1 ^ tmp_278_fu_11644_p4);

assign xor_ln1545_396_fu_11868_p2 = (tmp_V_129_reg_16296 ^ tmp_V_128_reg_16266);

assign xor_ln1545_397_fu_11878_p2 = (xor_ln1545_398_fu_11872_p2 ^ xor_ln1545_396_fu_11868_p2);

assign xor_ln1545_398_fu_11872_p2 = (trunc_ln674_131_fu_11640_p1 ^ tmp_279_fu_11658_p4);

assign xor_ln1545_399_fu_11884_p2 = (tmp_V_130_reg_16326 ^ tmp_V_129_reg_16296);

assign xor_ln1545_39_fu_5332_p2 = (tmp_V_9_reg_14296 ^ tmp_2_1_V_12_reg_14230);

assign xor_ln1545_400_fu_11894_p2 = (xor_ln1545_401_fu_11888_p2 ^ xor_ln1545_399_fu_11884_p2);

assign xor_ln1545_401_fu_11888_p2 = (trunc_ln674_132_fu_11654_p1 ^ tmp_276_fu_11616_p4);

assign xor_ln1545_402_fu_11900_p2 = (tmp_V_135_reg_16284 ^ tmp_V_134_reg_16350);

assign xor_ln1545_403_fu_11910_p2 = (xor_ln1545_404_fu_11904_p2 ^ xor_ln1545_402_fu_11900_p2);

assign xor_ln1545_404_fu_11904_p2 = (trunc_ln674_133_fu_11668_p1 ^ tmp_281_fu_11686_p4);

assign xor_ln1545_405_fu_11916_p2 = (tmp_V_135_reg_16284 ^ tmp_V_132_reg_16290);

assign xor_ln1545_406_fu_11926_p2 = (xor_ln1545_407_fu_11920_p2 ^ xor_ln1545_405_fu_11916_p2);

assign xor_ln1545_407_fu_11920_p2 = (trunc_ln674_134_fu_11682_p1 ^ tmp_282_fu_11700_p4);

assign xor_ln1545_408_fu_11932_p2 = (tmp_V_133_reg_16320 ^ tmp_V_132_reg_16290);

assign xor_ln1545_409_fu_11942_p2 = (xor_ln1545_410_fu_11936_p2 ^ xor_ln1545_408_fu_11932_p2);

assign xor_ln1545_40_fu_5342_p2 = (xor_ln1545_41_fu_5336_p2 ^ xor_ln1545_39_fu_5332_p2);

assign xor_ln1545_410_fu_11936_p2 = (trunc_ln674_135_fu_11696_p1 ^ tmp_283_fu_11714_p4);

assign xor_ln1545_411_fu_11948_p2 = (tmp_V_134_reg_16350 ^ tmp_V_133_reg_16320);

assign xor_ln1545_412_fu_11958_p2 = (xor_ln1545_413_fu_11952_p2 ^ xor_ln1545_411_fu_11948_p2);

assign xor_ln1545_413_fu_11952_p2 = (trunc_ln674_136_fu_11710_p1 ^ tmp_280_fu_11672_p4);

assign xor_ln1545_414_fu_11964_p2 = (tmp_V_139_reg_16308 ^ tmp_2_1_V_20_reg_16278);

assign xor_ln1545_415_fu_11974_p2 = (xor_ln1545_416_fu_11968_p2 ^ xor_ln1545_414_fu_11964_p2);

assign xor_ln1545_416_fu_11968_p2 = (trunc_ln674_137_fu_11724_p1 ^ tmp_285_fu_11742_p4);

assign xor_ln1545_417_fu_11980_p2 = (tmp_V_139_reg_16308 ^ tmp_V_136_reg_16314);

assign xor_ln1545_418_fu_11990_p2 = (xor_ln1545_419_fu_11984_p2 ^ xor_ln1545_417_fu_11980_p2);

assign xor_ln1545_419_fu_11984_p2 = (trunc_ln674_138_fu_11738_p1 ^ tmp_286_fu_11756_p4);

assign xor_ln1545_41_fu_5336_p2 = (trunc_ln674_12_fu_5086_p1 ^ tmp_36_fu_5048_p4);

assign xor_ln1545_420_fu_11996_p2 = (tmp_V_137_reg_16344 ^ tmp_V_136_reg_16314);

assign xor_ln1545_421_fu_12006_p2 = (xor_ln1545_422_fu_12000_p2 ^ xor_ln1545_420_fu_11996_p2);

assign xor_ln1545_422_fu_12000_p2 = (trunc_ln674_139_fu_11752_p1 ^ tmp_287_fu_11770_p4);

assign xor_ln1545_423_fu_12012_p2 = (tmp_V_137_reg_16344 ^ tmp_2_1_V_20_reg_16278);

assign xor_ln1545_424_fu_12022_p2 = (xor_ln1545_425_fu_12016_p2 ^ xor_ln1545_423_fu_12012_p2);

assign xor_ln1545_425_fu_12016_p2 = (trunc_ln674_140_fu_11766_p1 ^ tmp_284_fu_11728_p4);

assign xor_ln1545_426_fu_12028_p2 = (tmp_V_143_reg_16332 ^ tmp_2_2_V_20_reg_16302);

assign xor_ln1545_427_fu_12038_p2 = (xor_ln1545_428_fu_12032_p2 ^ xor_ln1545_426_fu_12028_p2);

assign xor_ln1545_428_fu_12032_p2 = (trunc_ln674_141_fu_11780_p1 ^ tmp_289_fu_11798_p4);

assign xor_ln1545_429_fu_12044_p2 = (tmp_V_143_reg_16332 ^ tmp_V_140_reg_16338);

assign xor_ln1545_42_fu_5348_p2 = (tmp_V_15_reg_14284 ^ tmp_2_2_V_12_reg_14254);

assign xor_ln1545_430_fu_12054_p2 = (xor_ln1545_431_fu_12048_p2 ^ xor_ln1545_429_fu_12044_p2);

assign xor_ln1545_431_fu_12048_p2 = (trunc_ln674_142_fu_11794_p1 ^ tmp_290_fu_11812_p4);

assign xor_ln1545_432_fu_12060_p2 = (tmp_V_140_reg_16338 ^ tmp_1_V_20_reg_16272);

assign xor_ln1545_433_fu_12070_p2 = (xor_ln1545_434_fu_12064_p2 ^ xor_ln1545_432_fu_12060_p2);

assign xor_ln1545_434_fu_12064_p2 = (trunc_ln674_143_fu_11808_p1 ^ tmp_291_fu_11826_p4);

assign xor_ln1545_435_fu_12076_p2 = (tmp_2_2_V_20_reg_16302 ^ tmp_1_V_20_reg_16272);

assign xor_ln1545_436_fu_12086_p2 = (xor_ln1545_437_fu_12080_p2 ^ xor_ln1545_435_fu_12076_p2);

assign xor_ln1545_437_fu_12080_p2 = (trunc_ln674_144_fu_11822_p1 ^ tmp_288_fu_11784_p4);

assign xor_ln1545_438_fu_12671_p2 = (tmp_V_146_reg_16582 ^ tmp_3_V_21_reg_16612);

assign xor_ln1545_439_fu_12681_p2 = (xor_ln1545_440_fu_12675_p2 ^ xor_ln1545_438_fu_12671_p2);

assign xor_ln1545_43_fu_5358_p2 = (xor_ln1545_44_fu_5352_p2 ^ xor_ln1545_42_fu_5348_p2);

assign xor_ln1545_440_fu_12675_p2 = (trunc_ln674_145_fu_12447_p1 ^ tmp_308_fu_12465_p4);

assign xor_ln1545_441_fu_12687_p2 = (tmp_V_144_reg_16522 ^ tmp_3_V_21_reg_16612);

assign xor_ln1545_442_fu_12697_p2 = (xor_ln1545_443_fu_12691_p2 ^ xor_ln1545_441_fu_12687_p2);

assign xor_ln1545_443_fu_12691_p2 = (trunc_ln674_146_fu_12461_p1 ^ tmp_309_fu_12479_p4);

assign xor_ln1545_444_fu_12703_p2 = (tmp_V_145_reg_16552 ^ tmp_V_144_reg_16522);

assign xor_ln1545_445_fu_12713_p2 = (xor_ln1545_446_fu_12707_p2 ^ xor_ln1545_444_fu_12703_p2);

assign xor_ln1545_446_fu_12707_p2 = (trunc_ln674_147_fu_12475_p1 ^ tmp_310_fu_12493_p4);

assign xor_ln1545_447_fu_12719_p2 = (tmp_V_146_reg_16582 ^ tmp_V_145_reg_16552);

assign xor_ln1545_448_fu_12729_p2 = (xor_ln1545_449_fu_12723_p2 ^ xor_ln1545_447_fu_12719_p2);

assign xor_ln1545_449_fu_12723_p2 = (trunc_ln674_148_fu_12489_p1 ^ tmp_307_fu_12451_p4);

assign xor_ln1545_44_fu_5352_p2 = (trunc_ln674_13_fu_5100_p1 ^ tmp_41_fu_5118_p4);

assign xor_ln1545_450_fu_12735_p2 = (tmp_V_151_reg_16540 ^ tmp_V_150_reg_16606);

assign xor_ln1545_451_fu_12745_p2 = (xor_ln1545_452_fu_12739_p2 ^ xor_ln1545_450_fu_12735_p2);

assign xor_ln1545_452_fu_12739_p2 = (trunc_ln674_149_fu_12503_p1 ^ tmp_312_fu_12521_p4);

assign xor_ln1545_453_fu_12751_p2 = (tmp_V_151_reg_16540 ^ tmp_V_148_reg_16546);

assign xor_ln1545_454_fu_12761_p2 = (xor_ln1545_455_fu_12755_p2 ^ xor_ln1545_453_fu_12751_p2);

assign xor_ln1545_455_fu_12755_p2 = (trunc_ln674_150_fu_12517_p1 ^ tmp_313_fu_12535_p4);

assign xor_ln1545_456_fu_12767_p2 = (tmp_V_149_reg_16576 ^ tmp_V_148_reg_16546);

assign xor_ln1545_457_fu_12777_p2 = (xor_ln1545_458_fu_12771_p2 ^ xor_ln1545_456_fu_12767_p2);

assign xor_ln1545_458_fu_12771_p2 = (trunc_ln674_151_fu_12531_p1 ^ tmp_314_fu_12549_p4);

assign xor_ln1545_459_fu_12783_p2 = (tmp_V_150_reg_16606 ^ tmp_V_149_reg_16576);

assign xor_ln1545_45_fu_5364_p2 = (tmp_V_15_reg_14284 ^ tmp_V_12_reg_14290);

assign xor_ln1545_460_fu_12793_p2 = (xor_ln1545_461_fu_12787_p2 ^ xor_ln1545_459_fu_12783_p2);

assign xor_ln1545_461_fu_12787_p2 = (trunc_ln674_152_fu_12545_p1 ^ tmp_311_fu_12507_p4);

assign xor_ln1545_462_fu_12799_p2 = (tmp_V_155_reg_16564 ^ tmp_2_1_V_21_reg_16534);

assign xor_ln1545_463_fu_12809_p2 = (xor_ln1545_464_fu_12803_p2 ^ xor_ln1545_462_fu_12799_p2);

assign xor_ln1545_464_fu_12803_p2 = (trunc_ln674_153_fu_12559_p1 ^ tmp_316_fu_12577_p4);

assign xor_ln1545_465_fu_12815_p2 = (tmp_V_155_reg_16564 ^ tmp_V_152_reg_16570);

assign xor_ln1545_466_fu_12825_p2 = (xor_ln1545_467_fu_12819_p2 ^ xor_ln1545_465_fu_12815_p2);

assign xor_ln1545_467_fu_12819_p2 = (trunc_ln674_154_fu_12573_p1 ^ tmp_317_fu_12591_p4);

assign xor_ln1545_468_fu_12831_p2 = (tmp_V_153_reg_16600 ^ tmp_V_152_reg_16570);

assign xor_ln1545_469_fu_12841_p2 = (xor_ln1545_470_fu_12835_p2 ^ xor_ln1545_468_fu_12831_p2);

assign xor_ln1545_46_fu_5374_p2 = (xor_ln1545_47_fu_5368_p2 ^ xor_ln1545_45_fu_5364_p2);

assign xor_ln1545_470_fu_12835_p2 = (trunc_ln674_155_fu_12587_p1 ^ tmp_318_fu_12605_p4);

assign xor_ln1545_471_fu_12847_p2 = (tmp_V_153_reg_16600 ^ tmp_2_1_V_21_reg_16534);

assign xor_ln1545_472_fu_12857_p2 = (xor_ln1545_473_fu_12851_p2 ^ xor_ln1545_471_fu_12847_p2);

assign xor_ln1545_473_fu_12851_p2 = (trunc_ln674_156_fu_12601_p1 ^ tmp_315_fu_12563_p4);

assign xor_ln1545_474_fu_12863_p2 = (tmp_V_159_reg_16588 ^ tmp_2_2_V_21_reg_16558);

assign xor_ln1545_475_fu_12873_p2 = (xor_ln1545_476_fu_12867_p2 ^ xor_ln1545_474_fu_12863_p2);

assign xor_ln1545_476_fu_12867_p2 = (trunc_ln674_157_fu_12615_p1 ^ tmp_320_fu_12633_p4);

assign xor_ln1545_477_fu_12879_p2 = (tmp_V_159_reg_16588 ^ tmp_V_156_reg_16594);

assign xor_ln1545_478_fu_12889_p2 = (xor_ln1545_479_fu_12883_p2 ^ xor_ln1545_477_fu_12879_p2);

assign xor_ln1545_479_fu_12883_p2 = (trunc_ln674_158_fu_12629_p1 ^ tmp_321_fu_12647_p4);

assign xor_ln1545_47_fu_5368_p2 = (trunc_ln674_14_fu_5114_p1 ^ tmp_42_fu_5132_p4);

assign xor_ln1545_480_fu_12895_p2 = (tmp_V_156_reg_16594 ^ tmp_1_V_21_reg_16528);

assign xor_ln1545_481_fu_12905_p2 = (xor_ln1545_482_fu_12899_p2 ^ xor_ln1545_480_fu_12895_p2);

assign xor_ln1545_482_fu_12899_p2 = (trunc_ln674_159_fu_12643_p1 ^ tmp_322_fu_12661_p4);

assign xor_ln1545_483_fu_12911_p2 = (tmp_2_2_V_21_reg_16558 ^ tmp_1_V_21_reg_16528);

assign xor_ln1545_484_fu_12921_p2 = (xor_ln1545_485_fu_12915_p2 ^ xor_ln1545_483_fu_12911_p2);

assign xor_ln1545_485_fu_12915_p2 = (trunc_ln674_160_fu_12657_p1 ^ tmp_319_fu_12619_p4);

assign xor_ln1545_486_fu_13506_p2 = (tmp_V_162_reg_16838 ^ tmp_3_V_22_reg_16868);

assign xor_ln1545_487_fu_13516_p2 = (xor_ln1545_488_fu_13510_p2 ^ xor_ln1545_486_fu_13506_p2);

assign xor_ln1545_488_fu_13510_p2 = (trunc_ln674_161_fu_13282_p1 ^ tmp_339_fu_13300_p4);

assign xor_ln1545_489_fu_13522_p2 = (tmp_V_160_reg_16778 ^ tmp_3_V_22_reg_16868);

assign xor_ln1545_48_fu_5380_p2 = (tmp_V_12_reg_14290 ^ tmp_1_V_12_reg_14224);

assign xor_ln1545_490_fu_13532_p2 = (xor_ln1545_491_fu_13526_p2 ^ xor_ln1545_489_fu_13522_p2);

assign xor_ln1545_491_fu_13526_p2 = (trunc_ln674_162_fu_13296_p1 ^ tmp_340_fu_13314_p4);

assign xor_ln1545_492_fu_13538_p2 = (tmp_V_161_reg_16808 ^ tmp_V_160_reg_16778);

assign xor_ln1545_493_fu_13548_p2 = (xor_ln1545_494_fu_13542_p2 ^ xor_ln1545_492_fu_13538_p2);

assign xor_ln1545_494_fu_13542_p2 = (trunc_ln674_163_fu_13310_p1 ^ tmp_341_fu_13328_p4);

assign xor_ln1545_495_fu_13554_p2 = (tmp_V_162_reg_16838 ^ tmp_V_161_reg_16808);

assign xor_ln1545_496_fu_13564_p2 = (xor_ln1545_497_fu_13558_p2 ^ xor_ln1545_495_fu_13554_p2);

assign xor_ln1545_497_fu_13558_p2 = (trunc_ln674_164_fu_13324_p1 ^ tmp_338_fu_13286_p4);

assign xor_ln1545_498_fu_13570_p2 = (tmp_V_167_reg_16796 ^ tmp_V_166_reg_16862);

assign xor_ln1545_499_fu_13580_p2 = (xor_ln1545_500_fu_13574_p2 ^ xor_ln1545_498_fu_13570_p2);

assign xor_ln1545_49_fu_5390_p2 = (xor_ln1545_50_fu_5384_p2 ^ xor_ln1545_48_fu_5380_p2);

assign xor_ln1545_500_fu_13574_p2 = (trunc_ln674_165_fu_13338_p1 ^ tmp_343_fu_13356_p4);

assign xor_ln1545_501_fu_13586_p2 = (tmp_V_167_reg_16796 ^ tmp_V_164_reg_16802);

assign xor_ln1545_502_fu_13596_p2 = (xor_ln1545_503_fu_13590_p2 ^ xor_ln1545_501_fu_13586_p2);

assign xor_ln1545_503_fu_13590_p2 = (trunc_ln674_166_fu_13352_p1 ^ tmp_344_fu_13370_p4);

assign xor_ln1545_504_fu_13602_p2 = (tmp_V_165_reg_16832 ^ tmp_V_164_reg_16802);

assign xor_ln1545_505_fu_13612_p2 = (xor_ln1545_506_fu_13606_p2 ^ xor_ln1545_504_fu_13602_p2);

assign xor_ln1545_506_fu_13606_p2 = (trunc_ln674_167_fu_13366_p1 ^ tmp_345_fu_13384_p4);

assign xor_ln1545_507_fu_13618_p2 = (tmp_V_166_reg_16862 ^ tmp_V_165_reg_16832);

assign xor_ln1545_508_fu_13628_p2 = (xor_ln1545_509_fu_13622_p2 ^ xor_ln1545_507_fu_13618_p2);

assign xor_ln1545_509_fu_13622_p2 = (trunc_ln674_168_fu_13380_p1 ^ tmp_342_fu_13342_p4);

assign xor_ln1545_50_fu_5384_p2 = (trunc_ln674_15_fu_5128_p1 ^ tmp_43_fu_5146_p4);

assign xor_ln1545_510_fu_13634_p2 = (tmp_V_171_reg_16820 ^ tmp_2_1_V_22_reg_16790);

assign xor_ln1545_511_fu_13644_p2 = (xor_ln1545_512_fu_13638_p2 ^ xor_ln1545_510_fu_13634_p2);

assign xor_ln1545_512_fu_13638_p2 = (trunc_ln674_169_fu_13394_p1 ^ tmp_347_fu_13412_p4);

assign xor_ln1545_513_fu_13650_p2 = (tmp_V_171_reg_16820 ^ tmp_V_168_reg_16826);

assign xor_ln1545_514_fu_13660_p2 = (xor_ln1545_515_fu_13654_p2 ^ xor_ln1545_513_fu_13650_p2);

assign xor_ln1545_515_fu_13654_p2 = (trunc_ln674_170_fu_13408_p1 ^ tmp_348_fu_13426_p4);

assign xor_ln1545_516_fu_13666_p2 = (tmp_V_169_reg_16856 ^ tmp_V_168_reg_16826);

assign xor_ln1545_517_fu_13676_p2 = (xor_ln1545_518_fu_13670_p2 ^ xor_ln1545_516_fu_13666_p2);

assign xor_ln1545_518_fu_13670_p2 = (trunc_ln674_171_fu_13422_p1 ^ tmp_349_fu_13440_p4);

assign xor_ln1545_519_fu_13682_p2 = (tmp_V_169_reg_16856 ^ tmp_2_1_V_22_reg_16790);

assign xor_ln1545_51_fu_5396_p2 = (tmp_2_2_V_12_reg_14254 ^ tmp_1_V_12_reg_14224);

assign xor_ln1545_520_fu_13692_p2 = (xor_ln1545_521_fu_13686_p2 ^ xor_ln1545_519_fu_13682_p2);

assign xor_ln1545_521_fu_13686_p2 = (trunc_ln674_172_fu_13436_p1 ^ tmp_346_fu_13398_p4);

assign xor_ln1545_522_fu_13698_p2 = (tmp_V_175_reg_16844 ^ tmp_2_2_V_22_reg_16814);

assign xor_ln1545_523_fu_13708_p2 = (xor_ln1545_524_fu_13702_p2 ^ xor_ln1545_522_fu_13698_p2);

assign xor_ln1545_524_fu_13702_p2 = (trunc_ln674_173_fu_13450_p1 ^ tmp_351_fu_13468_p4);

assign xor_ln1545_525_fu_13714_p2 = (tmp_V_175_reg_16844 ^ tmp_V_172_reg_16850);

assign xor_ln1545_526_fu_13724_p2 = (xor_ln1545_527_fu_13718_p2 ^ xor_ln1545_525_fu_13714_p2);

assign xor_ln1545_527_fu_13718_p2 = (trunc_ln674_174_fu_13464_p1 ^ tmp_352_fu_13482_p4);

assign xor_ln1545_528_fu_13730_p2 = (tmp_V_172_reg_16850 ^ tmp_1_V_22_reg_16784);

assign xor_ln1545_529_fu_13740_p2 = (xor_ln1545_530_fu_13734_p2 ^ xor_ln1545_528_fu_13730_p2);

assign xor_ln1545_52_fu_5406_p2 = (xor_ln1545_53_fu_5400_p2 ^ xor_ln1545_51_fu_5396_p2);

assign xor_ln1545_530_fu_13734_p2 = (trunc_ln674_175_fu_13478_p1 ^ tmp_353_fu_13496_p4);

assign xor_ln1545_531_fu_13746_p2 = (tmp_2_2_V_22_reg_16814 ^ tmp_1_V_22_reg_16784);

assign xor_ln1545_532_fu_13756_p2 = (xor_ln1545_533_fu_13750_p2 ^ xor_ln1545_531_fu_13746_p2);

assign xor_ln1545_533_fu_13750_p2 = (trunc_ln674_176_fu_13492_p1 ^ tmp_350_fu_13454_p4);

assign xor_ln1545_53_fu_5400_p2 = (trunc_ln674_16_fu_5142_p1 ^ tmp_40_fu_5104_p4);

assign xor_ln1545_54_fu_5991_p2 = (tmp_V_18_reg_14534 ^ tmp_3_V_13_reg_14564);

assign xor_ln1545_55_fu_6001_p2 = (xor_ln1545_56_fu_5995_p2 ^ xor_ln1545_54_fu_5991_p2);

assign xor_ln1545_56_fu_5995_p2 = (trunc_ln674_17_fu_5767_p1 ^ tmp_60_fu_5785_p4);

assign xor_ln1545_57_fu_6007_p2 = (tmp_V_16_reg_14474 ^ tmp_3_V_13_reg_14564);

assign xor_ln1545_58_fu_6017_p2 = (xor_ln1545_59_fu_6011_p2 ^ xor_ln1545_57_fu_6007_p2);

assign xor_ln1545_59_fu_6011_p2 = (trunc_ln674_18_fu_5781_p1 ^ tmp_61_fu_5799_p4);

assign xor_ln1545_60_fu_6023_p2 = (tmp_V_17_reg_14504 ^ tmp_V_16_reg_14474);

assign xor_ln1545_61_fu_6033_p2 = (xor_ln1545_62_fu_6027_p2 ^ xor_ln1545_60_fu_6023_p2);

assign xor_ln1545_62_fu_6027_p2 = (trunc_ln674_19_fu_5795_p1 ^ tmp_62_fu_5813_p4);

assign xor_ln1545_63_fu_6039_p2 = (tmp_V_18_reg_14534 ^ tmp_V_17_reg_14504);

assign xor_ln1545_64_fu_6049_p2 = (xor_ln1545_65_fu_6043_p2 ^ xor_ln1545_63_fu_6039_p2);

assign xor_ln1545_65_fu_6043_p2 = (trunc_ln674_20_fu_5809_p1 ^ tmp_59_fu_5771_p4);

assign xor_ln1545_66_fu_6055_p2 = (tmp_V_23_reg_14492 ^ tmp_V_22_reg_14558);

assign xor_ln1545_67_fu_6065_p2 = (xor_ln1545_68_fu_6059_p2 ^ xor_ln1545_66_fu_6055_p2);

assign xor_ln1545_68_fu_6059_p2 = (trunc_ln674_21_fu_5823_p1 ^ tmp_64_fu_5841_p4);

assign xor_ln1545_69_fu_6071_p2 = (tmp_V_23_reg_14492 ^ tmp_V_20_reg_14498);

assign xor_ln1545_70_fu_6081_p2 = (xor_ln1545_71_fu_6075_p2 ^ xor_ln1545_69_fu_6071_p2);

assign xor_ln1545_71_fu_6075_p2 = (trunc_ln674_22_fu_5837_p1 ^ tmp_65_fu_5855_p4);

assign xor_ln1545_72_fu_6087_p2 = (tmp_V_21_reg_14528 ^ tmp_V_20_reg_14498);

assign xor_ln1545_73_fu_6097_p2 = (xor_ln1545_74_fu_6091_p2 ^ xor_ln1545_72_fu_6087_p2);

assign xor_ln1545_74_fu_6091_p2 = (trunc_ln674_23_fu_5851_p1 ^ tmp_66_fu_5869_p4);

assign xor_ln1545_75_fu_6103_p2 = (tmp_V_22_reg_14558 ^ tmp_V_21_reg_14528);

assign xor_ln1545_76_fu_6113_p2 = (xor_ln1545_77_fu_6107_p2 ^ xor_ln1545_75_fu_6103_p2);

assign xor_ln1545_77_fu_6107_p2 = (trunc_ln674_24_fu_5865_p1 ^ tmp_63_fu_5827_p4);

assign xor_ln1545_78_fu_6119_p2 = (tmp_V_27_reg_14516 ^ tmp_2_1_V_13_reg_14486);

assign xor_ln1545_79_fu_6129_p2 = (xor_ln1545_80_fu_6123_p2 ^ xor_ln1545_78_fu_6119_p2);

assign xor_ln1545_7_fu_5166_p2 = (xor_ln1545_fu_5156_p2 ^ xor_ln1545_8_fu_5160_p2);

assign xor_ln1545_80_fu_6123_p2 = (trunc_ln674_25_fu_5879_p1 ^ tmp_68_fu_5897_p4);

assign xor_ln1545_81_fu_6135_p2 = (tmp_V_27_reg_14516 ^ tmp_V_24_reg_14522);

assign xor_ln1545_82_fu_6145_p2 = (xor_ln1545_83_fu_6139_p2 ^ xor_ln1545_81_fu_6135_p2);

assign xor_ln1545_83_fu_6139_p2 = (trunc_ln674_26_fu_5893_p1 ^ tmp_69_fu_5911_p4);

assign xor_ln1545_84_fu_6151_p2 = (tmp_V_25_reg_14552 ^ tmp_V_24_reg_14522);

assign xor_ln1545_85_fu_6161_p2 = (xor_ln1545_86_fu_6155_p2 ^ xor_ln1545_84_fu_6151_p2);

assign xor_ln1545_86_fu_6155_p2 = (trunc_ln674_27_fu_5907_p1 ^ tmp_70_fu_5925_p4);

assign xor_ln1545_87_fu_6167_p2 = (tmp_V_25_reg_14552 ^ tmp_2_1_V_13_reg_14486);

assign xor_ln1545_88_fu_6177_p2 = (xor_ln1545_89_fu_6171_p2 ^ xor_ln1545_87_fu_6167_p2);

assign xor_ln1545_89_fu_6171_p2 = (trunc_ln674_28_fu_5921_p1 ^ tmp_67_fu_5883_p4);

assign xor_ln1545_8_fu_5160_p2 = (trunc_ln674_fu_4932_p1 ^ tmp_29_fu_4950_p4);

assign xor_ln1545_90_fu_6183_p2 = (tmp_V_31_reg_14540 ^ tmp_2_2_V_13_reg_14510);

assign xor_ln1545_91_fu_6193_p2 = (xor_ln1545_92_fu_6187_p2 ^ xor_ln1545_90_fu_6183_p2);

assign xor_ln1545_92_fu_6187_p2 = (trunc_ln674_29_fu_5935_p1 ^ tmp_72_fu_5953_p4);

assign xor_ln1545_93_fu_6199_p2 = (tmp_V_31_reg_14540 ^ tmp_V_28_reg_14546);

assign xor_ln1545_94_fu_6209_p2 = (xor_ln1545_95_fu_6203_p2 ^ xor_ln1545_93_fu_6199_p2);

assign xor_ln1545_95_fu_6203_p2 = (trunc_ln674_30_fu_5949_p1 ^ tmp_73_fu_5967_p4);

assign xor_ln1545_96_fu_6215_p2 = (tmp_V_28_reg_14546 ^ tmp_1_V_13_reg_14480);

assign xor_ln1545_97_fu_6225_p2 = (xor_ln1545_98_fu_6219_p2 ^ xor_ln1545_96_fu_6215_p2);

assign xor_ln1545_98_fu_6219_p2 = (trunc_ln674_31_fu_5963_p1 ^ tmp_74_fu_5981_p4);

assign xor_ln1545_99_fu_6231_p2 = (tmp_2_2_V_13_reg_14510 ^ tmp_1_V_13_reg_14480);

assign xor_ln1545_9_fu_5172_p2 = (tmp_V_reg_14218 ^ tmp_3_V_12_reg_14308);

assign xor_ln1545_fu_5156_p2 = (tmp_V_2_reg_14278 ^ tmp_3_V_12_reg_14308);

assign zext_ln587_100_fu_9882_p1 = cipher_0_ssbox_q91;

assign zext_ln587_101_fu_9887_p1 = cipher_0_ssbox_q86;

assign zext_ln587_102_fu_9892_p1 = cipher_0_ssbox_q81;

assign zext_ln587_103_fu_9897_p1 = cipher_0_ssbox_q92;

assign zext_ln587_104_fu_9902_p1 = cipher_0_ssbox_q87;

assign zext_ln587_105_fu_9907_p1 = cipher_0_ssbox_q82;

assign zext_ln587_106_fu_9912_p1 = cipher_0_ssbox_q93;

assign zext_ln587_107_fu_9917_p1 = cipher_0_ssbox_q88;

assign zext_ln587_108_fu_9922_p1 = cipher_0_ssbox_q83;

assign zext_ln587_109_fu_9927_p1 = cipher_0_ssbox_q94;

assign zext_ln587_10_fu_4902_p1 = cipher_0_ssbox_q189;

assign zext_ln587_110_fu_9932_p1 = cipher_0_ssbox_q89;

assign zext_ln587_111_fu_9937_p1 = cipher_0_ssbox_q84;

assign zext_ln587_112_fu_10697_p1 = cipher_0_ssbox_q79;

assign zext_ln587_113_fu_10702_p1 = cipher_0_ssbox_q74;

assign zext_ln587_114_fu_10707_p1 = cipher_0_ssbox_q69;

assign zext_ln587_115_fu_10712_p1 = cipher_0_ssbox_q64;

assign zext_ln587_116_fu_10717_p1 = cipher_0_ssbox_q75;

assign zext_ln587_117_fu_10722_p1 = cipher_0_ssbox_q70;

assign zext_ln587_118_fu_10727_p1 = cipher_0_ssbox_q65;

assign zext_ln587_119_fu_10732_p1 = cipher_0_ssbox_q76;

assign zext_ln587_11_fu_4907_p1 = cipher_0_ssbox_q184;

assign zext_ln587_120_fu_10737_p1 = cipher_0_ssbox_q71;

assign zext_ln587_121_fu_10742_p1 = cipher_0_ssbox_q66;

assign zext_ln587_122_fu_10747_p1 = cipher_0_ssbox_q77;

assign zext_ln587_123_fu_10752_p1 = cipher_0_ssbox_q72;

assign zext_ln587_124_fu_10757_p1 = cipher_0_ssbox_q67;

assign zext_ln587_125_fu_10762_p1 = cipher_0_ssbox_q78;

assign zext_ln587_126_fu_10767_p1 = cipher_0_ssbox_q73;

assign zext_ln587_127_fu_10772_p1 = cipher_0_ssbox_q68;

assign zext_ln587_128_fu_11532_p1 = cipher_0_ssbox_q63;

assign zext_ln587_129_fu_11537_p1 = cipher_0_ssbox_q58;

assign zext_ln587_12_fu_4912_p1 = cipher_0_ssbox_q179;

assign zext_ln587_130_fu_11542_p1 = cipher_0_ssbox_q53;

assign zext_ln587_131_fu_11547_p1 = cipher_0_ssbox_q48;

assign zext_ln587_132_fu_11552_p1 = cipher_0_ssbox_q59;

assign zext_ln587_133_fu_11557_p1 = cipher_0_ssbox_q54;

assign zext_ln587_134_fu_11562_p1 = cipher_0_ssbox_q49;

assign zext_ln587_135_fu_11567_p1 = cipher_0_ssbox_q60;

assign zext_ln587_136_fu_11572_p1 = cipher_0_ssbox_q55;

assign zext_ln587_137_fu_11577_p1 = cipher_0_ssbox_q50;

assign zext_ln587_138_fu_11582_p1 = cipher_0_ssbox_q61;

assign zext_ln587_139_fu_11587_p1 = cipher_0_ssbox_q56;

assign zext_ln587_13_fu_4917_p1 = cipher_0_ssbox_q190;

assign zext_ln587_140_fu_11592_p1 = cipher_0_ssbox_q51;

assign zext_ln587_141_fu_11597_p1 = cipher_0_ssbox_q62;

assign zext_ln587_142_fu_11602_p1 = cipher_0_ssbox_q57;

assign zext_ln587_143_fu_11607_p1 = cipher_0_ssbox_q52;

assign zext_ln587_144_fu_12367_p1 = cipher_0_ssbox_q47;

assign zext_ln587_145_fu_12372_p1 = cipher_0_ssbox_q42;

assign zext_ln587_146_fu_12377_p1 = cipher_0_ssbox_q37;

assign zext_ln587_147_fu_12382_p1 = cipher_0_ssbox_q32;

assign zext_ln587_148_fu_12387_p1 = cipher_0_ssbox_q43;

assign zext_ln587_149_fu_12392_p1 = cipher_0_ssbox_q38;

assign zext_ln587_14_fu_4922_p1 = cipher_0_ssbox_q185;

assign zext_ln587_150_fu_12397_p1 = cipher_0_ssbox_q33;

assign zext_ln587_151_fu_12402_p1 = cipher_0_ssbox_q44;

assign zext_ln587_152_fu_12407_p1 = cipher_0_ssbox_q39;

assign zext_ln587_153_fu_12412_p1 = cipher_0_ssbox_q34;

assign zext_ln587_154_fu_12417_p1 = cipher_0_ssbox_q45;

assign zext_ln587_155_fu_12422_p1 = cipher_0_ssbox_q40;

assign zext_ln587_156_fu_12427_p1 = cipher_0_ssbox_q35;

assign zext_ln587_157_fu_12432_p1 = cipher_0_ssbox_q46;

assign zext_ln587_158_fu_12437_p1 = cipher_0_ssbox_q41;

assign zext_ln587_159_fu_12442_p1 = cipher_0_ssbox_q36;

assign zext_ln587_15_fu_4927_p1 = cipher_0_ssbox_q180;

assign zext_ln587_160_fu_13202_p1 = cipher_0_ssbox_q31;

assign zext_ln587_161_fu_13207_p1 = cipher_0_ssbox_q26;

assign zext_ln587_162_fu_13212_p1 = cipher_0_ssbox_q21;

assign zext_ln587_163_fu_13217_p1 = cipher_0_ssbox_q16;

assign zext_ln587_164_fu_13222_p1 = cipher_0_ssbox_q27;

assign zext_ln587_165_fu_13227_p1 = cipher_0_ssbox_q22;

assign zext_ln587_166_fu_13232_p1 = cipher_0_ssbox_q17;

assign zext_ln587_167_fu_13237_p1 = cipher_0_ssbox_q28;

assign zext_ln587_168_fu_13242_p1 = cipher_0_ssbox_q23;

assign zext_ln587_169_fu_13247_p1 = cipher_0_ssbox_q18;

assign zext_ln587_16_fu_5687_p1 = cipher_0_ssbox_q175;

assign zext_ln587_170_fu_13252_p1 = cipher_0_ssbox_q29;

assign zext_ln587_171_fu_13257_p1 = cipher_0_ssbox_q24;

assign zext_ln587_172_fu_13262_p1 = cipher_0_ssbox_q19;

assign zext_ln587_173_fu_13267_p1 = cipher_0_ssbox_q30;

assign zext_ln587_174_fu_13272_p1 = cipher_0_ssbox_q25;

assign zext_ln587_175_fu_13277_p1 = cipher_0_ssbox_q20;

assign zext_ln587_17_fu_5692_p1 = cipher_0_ssbox_q170;

assign zext_ln587_18_fu_5697_p1 = cipher_0_ssbox_q165;

assign zext_ln587_19_fu_5702_p1 = cipher_0_ssbox_q160;

assign zext_ln587_1_fu_4857_p1 = cipher_0_ssbox_q186;

assign zext_ln587_20_fu_5707_p1 = cipher_0_ssbox_q171;

assign zext_ln587_21_fu_5712_p1 = cipher_0_ssbox_q166;

assign zext_ln587_22_fu_5717_p1 = cipher_0_ssbox_q161;

assign zext_ln587_23_fu_5722_p1 = cipher_0_ssbox_q172;

assign zext_ln587_24_fu_5727_p1 = cipher_0_ssbox_q167;

assign zext_ln587_25_fu_5732_p1 = cipher_0_ssbox_q162;

assign zext_ln587_26_fu_5737_p1 = cipher_0_ssbox_q173;

assign zext_ln587_27_fu_5742_p1 = cipher_0_ssbox_q168;

assign zext_ln587_28_fu_5747_p1 = cipher_0_ssbox_q163;

assign zext_ln587_29_fu_5752_p1 = cipher_0_ssbox_q174;

assign zext_ln587_2_fu_4862_p1 = cipher_0_ssbox_q181;

assign zext_ln587_30_fu_5757_p1 = cipher_0_ssbox_q169;

assign zext_ln587_31_fu_5762_p1 = cipher_0_ssbox_q164;

assign zext_ln587_32_fu_6522_p1 = cipher_0_ssbox_q159;

assign zext_ln587_33_fu_6527_p1 = cipher_0_ssbox_q154;

assign zext_ln587_34_fu_6532_p1 = cipher_0_ssbox_q149;

assign zext_ln587_35_fu_6537_p1 = cipher_0_ssbox_q144;

assign zext_ln587_36_fu_6542_p1 = cipher_0_ssbox_q155;

assign zext_ln587_37_fu_6547_p1 = cipher_0_ssbox_q150;

assign zext_ln587_38_fu_6552_p1 = cipher_0_ssbox_q145;

assign zext_ln587_39_fu_6557_p1 = cipher_0_ssbox_q156;

assign zext_ln587_3_fu_4867_p1 = cipher_0_ssbox_q176;

assign zext_ln587_40_fu_6562_p1 = cipher_0_ssbox_q151;

assign zext_ln587_41_fu_6567_p1 = cipher_0_ssbox_q146;

assign zext_ln587_42_fu_6572_p1 = cipher_0_ssbox_q157;

assign zext_ln587_43_fu_6577_p1 = cipher_0_ssbox_q152;

assign zext_ln587_44_fu_6582_p1 = cipher_0_ssbox_q147;

assign zext_ln587_45_fu_6587_p1 = cipher_0_ssbox_q158;

assign zext_ln587_46_fu_6592_p1 = cipher_0_ssbox_q153;

assign zext_ln587_47_fu_6597_p1 = cipher_0_ssbox_q148;

assign zext_ln587_48_fu_7357_p1 = cipher_0_ssbox_q143;

assign zext_ln587_49_fu_7362_p1 = cipher_0_ssbox_q138;

assign zext_ln587_4_fu_4872_p1 = cipher_0_ssbox_q187;

assign zext_ln587_50_fu_7367_p1 = cipher_0_ssbox_q133;

assign zext_ln587_51_fu_7372_p1 = cipher_0_ssbox_q128;

assign zext_ln587_52_fu_7377_p1 = cipher_0_ssbox_q139;

assign zext_ln587_53_fu_7382_p1 = cipher_0_ssbox_q134;

assign zext_ln587_54_fu_7387_p1 = cipher_0_ssbox_q129;

assign zext_ln587_55_fu_7392_p1 = cipher_0_ssbox_q140;

assign zext_ln587_56_fu_7397_p1 = cipher_0_ssbox_q135;

assign zext_ln587_57_fu_7402_p1 = cipher_0_ssbox_q130;

assign zext_ln587_58_fu_7407_p1 = cipher_0_ssbox_q141;

assign zext_ln587_59_fu_7412_p1 = cipher_0_ssbox_q136;

assign zext_ln587_5_fu_4877_p1 = cipher_0_ssbox_q182;

assign zext_ln587_60_fu_7417_p1 = cipher_0_ssbox_q131;

assign zext_ln587_61_fu_7422_p1 = cipher_0_ssbox_q142;

assign zext_ln587_62_fu_7427_p1 = cipher_0_ssbox_q137;

assign zext_ln587_63_fu_7432_p1 = cipher_0_ssbox_q132;

assign zext_ln587_64_fu_8192_p1 = cipher_0_ssbox_q127;

assign zext_ln587_65_fu_8197_p1 = cipher_0_ssbox_q122;

assign zext_ln587_66_fu_8202_p1 = cipher_0_ssbox_q117;

assign zext_ln587_67_fu_8207_p1 = cipher_0_ssbox_q112;

assign zext_ln587_68_fu_8212_p1 = cipher_0_ssbox_q123;

assign zext_ln587_69_fu_8217_p1 = cipher_0_ssbox_q118;

assign zext_ln587_6_fu_4882_p1 = cipher_0_ssbox_q177;

assign zext_ln587_70_fu_8222_p1 = cipher_0_ssbox_q113;

assign zext_ln587_71_fu_8227_p1 = cipher_0_ssbox_q124;

assign zext_ln587_72_fu_8232_p1 = cipher_0_ssbox_q119;

assign zext_ln587_73_fu_8237_p1 = cipher_0_ssbox_q114;

assign zext_ln587_74_fu_8242_p1 = cipher_0_ssbox_q125;

assign zext_ln587_75_fu_8247_p1 = cipher_0_ssbox_q120;

assign zext_ln587_76_fu_8252_p1 = cipher_0_ssbox_q115;

assign zext_ln587_77_fu_8257_p1 = cipher_0_ssbox_q126;

assign zext_ln587_78_fu_8262_p1 = cipher_0_ssbox_q121;

assign zext_ln587_79_fu_8267_p1 = cipher_0_ssbox_q116;

assign zext_ln587_7_fu_4887_p1 = cipher_0_ssbox_q188;

assign zext_ln587_80_fu_9027_p1 = cipher_0_ssbox_q111;

assign zext_ln587_81_fu_9032_p1 = cipher_0_ssbox_q106;

assign zext_ln587_82_fu_9037_p1 = cipher_0_ssbox_q101;

assign zext_ln587_83_fu_9042_p1 = cipher_0_ssbox_q96;

assign zext_ln587_84_fu_9047_p1 = cipher_0_ssbox_q107;

assign zext_ln587_85_fu_9052_p1 = cipher_0_ssbox_q102;

assign zext_ln587_86_fu_9057_p1 = cipher_0_ssbox_q97;

assign zext_ln587_87_fu_9062_p1 = cipher_0_ssbox_q108;

assign zext_ln587_88_fu_9067_p1 = cipher_0_ssbox_q103;

assign zext_ln587_89_fu_9072_p1 = cipher_0_ssbox_q98;

assign zext_ln587_8_fu_4892_p1 = cipher_0_ssbox_q183;

assign zext_ln587_90_fu_9077_p1 = cipher_0_ssbox_q109;

assign zext_ln587_91_fu_9082_p1 = cipher_0_ssbox_q104;

assign zext_ln587_92_fu_9087_p1 = cipher_0_ssbox_q99;

assign zext_ln587_93_fu_9092_p1 = cipher_0_ssbox_q110;

assign zext_ln587_94_fu_9097_p1 = cipher_0_ssbox_q105;

assign zext_ln587_95_fu_9102_p1 = cipher_0_ssbox_q100;

assign zext_ln587_96_fu_9862_p1 = cipher_0_ssbox_q95;

assign zext_ln587_97_fu_9867_p1 = cipher_0_ssbox_q90;

assign zext_ln587_98_fu_9872_p1 = cipher_0_ssbox_q85;

assign zext_ln587_99_fu_9877_p1 = cipher_0_ssbox_q80;

assign zext_ln587_9_fu_4897_p1 = cipher_0_ssbox_q178;

assign zext_ln587_fu_4852_p1 = cipher_0_ssbox_q191;

assign zext_ln708_100_fu_9647_p1 = tmp_199_fu_9637_p4;

assign zext_ln708_101_fu_9662_p1 = tmp_200_fu_9652_p4;

assign zext_ln708_102_fu_9677_p1 = tmp_201_fu_9667_p4;

assign zext_ln708_103_fu_9692_p1 = tmp_202_fu_9682_p4;

assign zext_ln708_104_fu_9707_p1 = tmp_203_fu_9697_p4;

assign zext_ln708_105_fu_9722_p1 = tmp_204_fu_9712_p4;

assign zext_ln708_106_fu_9737_p1 = tmp_205_fu_9727_p4;

assign zext_ln708_107_fu_9752_p1 = tmp_206_fu_9742_p4;

assign zext_ln708_108_fu_9767_p1 = tmp_207_fu_9757_p4;

assign zext_ln708_109_fu_9782_p1 = tmp_208_fu_9772_p4;

assign zext_ln708_10_fu_4727_p1 = tmp_19_fu_4717_p4;

assign zext_ln708_110_fu_9797_p1 = tmp_209_fu_9787_p4;

assign zext_ln708_111_fu_9812_p1 = tmp_210_fu_9802_p4;

assign zext_ln708_112_fu_9827_p1 = tmp_211_fu_9817_p4;

assign zext_ln708_113_fu_9842_p1 = tmp_212_fu_9832_p4;

assign zext_ln708_114_fu_9857_p1 = tmp_213_fu_9847_p4;

assign zext_ln708_115_fu_10467_p1 = trunc_ln708_7_fu_10463_p1;

assign zext_ln708_116_fu_10482_p1 = tmp_230_fu_10472_p4;

assign zext_ln708_117_fu_10497_p1 = tmp_231_fu_10487_p4;

assign zext_ln708_118_fu_10512_p1 = tmp_232_fu_10502_p4;

assign zext_ln708_119_fu_10527_p1 = tmp_233_fu_10517_p4;

assign zext_ln708_11_fu_4742_p1 = tmp_20_fu_4732_p4;

assign zext_ln708_120_fu_10542_p1 = tmp_234_fu_10532_p4;

assign zext_ln708_121_fu_10557_p1 = tmp_235_fu_10547_p4;

assign zext_ln708_122_fu_10572_p1 = tmp_236_fu_10562_p4;

assign zext_ln708_123_fu_10587_p1 = tmp_237_fu_10577_p4;

assign zext_ln708_124_fu_10602_p1 = tmp_238_fu_10592_p4;

assign zext_ln708_125_fu_10617_p1 = tmp_239_fu_10607_p4;

assign zext_ln708_126_fu_10632_p1 = tmp_240_fu_10622_p4;

assign zext_ln708_127_fu_10647_p1 = tmp_241_fu_10637_p4;

assign zext_ln708_128_fu_10662_p1 = tmp_242_fu_10652_p4;

assign zext_ln708_129_fu_10677_p1 = tmp_243_fu_10667_p4;

assign zext_ln708_12_fu_4757_p1 = tmp_21_fu_4747_p4;

assign zext_ln708_130_fu_10692_p1 = tmp_244_fu_10682_p4;

assign zext_ln708_131_fu_11302_p1 = trunc_ln708_8_fu_11298_p1;

assign zext_ln708_132_fu_11317_p1 = tmp_261_fu_11307_p4;

assign zext_ln708_133_fu_11332_p1 = tmp_262_fu_11322_p4;

assign zext_ln708_134_fu_11347_p1 = tmp_263_fu_11337_p4;

assign zext_ln708_135_fu_11362_p1 = tmp_264_fu_11352_p4;

assign zext_ln708_136_fu_11377_p1 = tmp_265_fu_11367_p4;

assign zext_ln708_137_fu_11392_p1 = tmp_266_fu_11382_p4;

assign zext_ln708_138_fu_11407_p1 = tmp_267_fu_11397_p4;

assign zext_ln708_139_fu_11422_p1 = tmp_268_fu_11412_p4;

assign zext_ln708_13_fu_4772_p1 = tmp_22_fu_4762_p4;

assign zext_ln708_140_fu_11437_p1 = tmp_269_fu_11427_p4;

assign zext_ln708_141_fu_11452_p1 = tmp_270_fu_11442_p4;

assign zext_ln708_142_fu_11467_p1 = tmp_271_fu_11457_p4;

assign zext_ln708_143_fu_11482_p1 = tmp_272_fu_11472_p4;

assign zext_ln708_144_fu_11497_p1 = tmp_273_fu_11487_p4;

assign zext_ln708_145_fu_11512_p1 = tmp_274_fu_11502_p4;

assign zext_ln708_146_fu_11527_p1 = tmp_275_fu_11517_p4;

assign zext_ln708_147_fu_12137_p1 = trunc_ln708_9_fu_12133_p1;

assign zext_ln708_148_fu_12152_p1 = tmp_292_fu_12142_p4;

assign zext_ln708_149_fu_12167_p1 = tmp_293_fu_12157_p4;

assign zext_ln708_14_fu_4787_p1 = tmp_23_fu_4777_p4;

assign zext_ln708_150_fu_12182_p1 = tmp_294_fu_12172_p4;

assign zext_ln708_151_fu_12197_p1 = tmp_295_fu_12187_p4;

assign zext_ln708_152_fu_12212_p1 = tmp_296_fu_12202_p4;

assign zext_ln708_153_fu_12227_p1 = tmp_297_fu_12217_p4;

assign zext_ln708_154_fu_12242_p1 = tmp_298_fu_12232_p4;

assign zext_ln708_155_fu_12257_p1 = tmp_299_fu_12247_p4;

assign zext_ln708_156_fu_12272_p1 = tmp_300_fu_12262_p4;

assign zext_ln708_157_fu_12287_p1 = tmp_301_fu_12277_p4;

assign zext_ln708_158_fu_12302_p1 = tmp_302_fu_12292_p4;

assign zext_ln708_159_fu_12317_p1 = tmp_303_fu_12307_p4;

assign zext_ln708_15_fu_4802_p1 = tmp_24_fu_4792_p4;

assign zext_ln708_160_fu_12332_p1 = tmp_304_fu_12322_p4;

assign zext_ln708_161_fu_12347_p1 = tmp_305_fu_12337_p4;

assign zext_ln708_162_fu_12362_p1 = tmp_306_fu_12352_p4;

assign zext_ln708_163_fu_12972_p1 = trunc_ln708_10_fu_12968_p1;

assign zext_ln708_164_fu_12987_p1 = tmp_323_fu_12977_p4;

assign zext_ln708_165_fu_13002_p1 = tmp_324_fu_12992_p4;

assign zext_ln708_166_fu_13017_p1 = tmp_325_fu_13007_p4;

assign zext_ln708_167_fu_13032_p1 = tmp_326_fu_13022_p4;

assign zext_ln708_168_fu_13047_p1 = tmp_327_fu_13037_p4;

assign zext_ln708_169_fu_13062_p1 = tmp_328_fu_13052_p4;

assign zext_ln708_16_fu_4817_p1 = tmp_25_fu_4807_p4;

assign zext_ln708_170_fu_13077_p1 = tmp_329_fu_13067_p4;

assign zext_ln708_171_fu_13092_p1 = tmp_330_fu_13082_p4;

assign zext_ln708_172_fu_13107_p1 = tmp_331_fu_13097_p4;

assign zext_ln708_173_fu_13122_p1 = tmp_332_fu_13112_p4;

assign zext_ln708_174_fu_13137_p1 = tmp_333_fu_13127_p4;

assign zext_ln708_175_fu_13152_p1 = tmp_334_fu_13142_p4;

assign zext_ln708_176_fu_13167_p1 = tmp_335_fu_13157_p4;

assign zext_ln708_177_fu_13182_p1 = tmp_336_fu_13172_p4;

assign zext_ln708_178_fu_13197_p1 = tmp_337_fu_13187_p4;

assign zext_ln708_179_fu_13807_p1 = trunc_ln708_11_fu_13803_p1;

assign zext_ln708_17_fu_4832_p1 = tmp_26_fu_4822_p4;

assign zext_ln708_180_fu_13822_p1 = tmp_354_fu_13812_p4;

assign zext_ln708_181_fu_13837_p1 = tmp_355_fu_13827_p4;

assign zext_ln708_182_fu_13852_p1 = tmp_356_fu_13842_p4;

assign zext_ln708_183_fu_13867_p1 = tmp_357_fu_13857_p4;

assign zext_ln708_184_fu_13882_p1 = tmp_358_fu_13872_p4;

assign zext_ln708_185_fu_13897_p1 = tmp_359_fu_13887_p4;

assign zext_ln708_186_fu_13912_p1 = tmp_360_fu_13902_p4;

assign zext_ln708_187_fu_13927_p1 = tmp_361_fu_13917_p4;

assign zext_ln708_188_fu_13942_p1 = tmp_362_fu_13932_p4;

assign zext_ln708_189_fu_13957_p1 = tmp_363_fu_13947_p4;

assign zext_ln708_18_fu_4847_p1 = tmp_27_fu_4837_p4;

assign zext_ln708_190_fu_13972_p1 = tmp_364_fu_13962_p4;

assign zext_ln708_191_fu_13987_p1 = tmp_365_fu_13977_p4;

assign zext_ln708_192_fu_14002_p1 = tmp_366_fu_13992_p4;

assign zext_ln708_193_fu_14017_p1 = tmp_367_fu_14007_p4;

assign zext_ln708_194_fu_14032_p1 = tmp_368_fu_14022_p4;

assign zext_ln708_19_fu_5457_p1 = trunc_ln708_1_fu_5453_p1;

assign zext_ln708_20_fu_5472_p1 = tmp_44_fu_5462_p4;

assign zext_ln708_21_fu_5487_p1 = tmp_45_fu_5477_p4;

assign zext_ln708_22_fu_5502_p1 = tmp_46_fu_5492_p4;

assign zext_ln708_23_fu_5517_p1 = tmp_47_fu_5507_p4;

assign zext_ln708_24_fu_5532_p1 = tmp_48_fu_5522_p4;

assign zext_ln708_25_fu_5547_p1 = tmp_49_fu_5537_p4;

assign zext_ln708_26_fu_5562_p1 = tmp_50_fu_5552_p4;

assign zext_ln708_27_fu_5577_p1 = tmp_51_fu_5567_p4;

assign zext_ln708_28_fu_5592_p1 = tmp_52_fu_5582_p4;

assign zext_ln708_29_fu_5607_p1 = tmp_53_fu_5597_p4;

assign zext_ln708_30_fu_5622_p1 = tmp_54_fu_5612_p4;

assign zext_ln708_31_fu_5637_p1 = tmp_55_fu_5627_p4;

assign zext_ln708_32_fu_5652_p1 = tmp_56_fu_5642_p4;

assign zext_ln708_33_fu_5667_p1 = tmp_57_fu_5657_p4;

assign zext_ln708_34_fu_5682_p1 = tmp_58_fu_5672_p4;

assign zext_ln708_35_fu_6292_p1 = trunc_ln708_2_fu_6288_p1;

assign zext_ln708_36_fu_6307_p1 = tmp_75_fu_6297_p4;

assign zext_ln708_37_fu_6322_p1 = tmp_76_fu_6312_p4;

assign zext_ln708_38_fu_6337_p1 = tmp_77_fu_6327_p4;

assign zext_ln708_39_fu_6352_p1 = tmp_78_fu_6342_p4;

assign zext_ln708_40_fu_6367_p1 = tmp_79_fu_6357_p4;

assign zext_ln708_41_fu_6382_p1 = tmp_80_fu_6372_p4;

assign zext_ln708_42_fu_6397_p1 = tmp_81_fu_6387_p4;

assign zext_ln708_43_fu_6412_p1 = tmp_82_fu_6402_p4;

assign zext_ln708_44_fu_6427_p1 = tmp_83_fu_6417_p4;

assign zext_ln708_45_fu_6442_p1 = tmp_84_fu_6432_p4;

assign zext_ln708_46_fu_6457_p1 = tmp_85_fu_6447_p4;

assign zext_ln708_47_fu_6472_p1 = tmp_86_fu_6462_p4;

assign zext_ln708_48_fu_6487_p1 = tmp_87_fu_6477_p4;

assign zext_ln708_49_fu_6502_p1 = tmp_88_fu_6492_p4;

assign zext_ln708_4_fu_4637_p1 = tmp_s_fu_4627_p4;

assign zext_ln708_50_fu_6517_p1 = tmp_89_fu_6507_p4;

assign zext_ln708_51_fu_7127_p1 = trunc_ln708_3_fu_7123_p1;

assign zext_ln708_52_fu_7142_p1 = tmp_106_fu_7132_p4;

assign zext_ln708_53_fu_7157_p1 = tmp_107_fu_7147_p4;

assign zext_ln708_54_fu_7172_p1 = tmp_108_fu_7162_p4;

assign zext_ln708_55_fu_7187_p1 = tmp_109_fu_7177_p4;

assign zext_ln708_56_fu_7202_p1 = tmp_110_fu_7192_p4;

assign zext_ln708_57_fu_7217_p1 = tmp_111_fu_7207_p4;

assign zext_ln708_58_fu_7232_p1 = tmp_112_fu_7222_p4;

assign zext_ln708_59_fu_7247_p1 = tmp_113_fu_7237_p4;

assign zext_ln708_5_fu_4652_p1 = tmp_14_fu_4642_p4;

assign zext_ln708_60_fu_7262_p1 = tmp_114_fu_7252_p4;

assign zext_ln708_61_fu_7277_p1 = tmp_115_fu_7267_p4;

assign zext_ln708_62_fu_7292_p1 = tmp_116_fu_7282_p4;

assign zext_ln708_63_fu_7307_p1 = tmp_117_fu_7297_p4;

assign zext_ln708_64_fu_7322_p1 = tmp_118_fu_7312_p4;

assign zext_ln708_65_fu_7337_p1 = tmp_119_fu_7327_p4;

assign zext_ln708_66_fu_7352_p1 = tmp_120_fu_7342_p4;

assign zext_ln708_67_fu_7962_p1 = trunc_ln708_4_fu_7958_p1;

assign zext_ln708_68_fu_7977_p1 = tmp_137_fu_7967_p4;

assign zext_ln708_69_fu_7992_p1 = tmp_138_fu_7982_p4;

assign zext_ln708_6_fu_4667_p1 = tmp_15_fu_4657_p4;

assign zext_ln708_70_fu_8007_p1 = tmp_139_fu_7997_p4;

assign zext_ln708_71_fu_8022_p1 = tmp_140_fu_8012_p4;

assign zext_ln708_72_fu_8037_p1 = tmp_141_fu_8027_p4;

assign zext_ln708_73_fu_8052_p1 = tmp_142_fu_8042_p4;

assign zext_ln708_74_fu_8067_p1 = tmp_143_fu_8057_p4;

assign zext_ln708_75_fu_8082_p1 = tmp_144_fu_8072_p4;

assign zext_ln708_76_fu_8097_p1 = tmp_145_fu_8087_p4;

assign zext_ln708_77_fu_8112_p1 = tmp_146_fu_8102_p4;

assign zext_ln708_78_fu_8127_p1 = tmp_147_fu_8117_p4;

assign zext_ln708_79_fu_8142_p1 = tmp_148_fu_8132_p4;

assign zext_ln708_7_fu_4682_p1 = tmp_16_fu_4672_p4;

assign zext_ln708_80_fu_8157_p1 = tmp_149_fu_8147_p4;

assign zext_ln708_81_fu_8172_p1 = tmp_150_fu_8162_p4;

assign zext_ln708_82_fu_8187_p1 = tmp_151_fu_8177_p4;

assign zext_ln708_83_fu_8797_p1 = trunc_ln708_5_fu_8793_p1;

assign zext_ln708_84_fu_8812_p1 = tmp_168_fu_8802_p4;

assign zext_ln708_85_fu_8827_p1 = tmp_169_fu_8817_p4;

assign zext_ln708_86_fu_8842_p1 = tmp_170_fu_8832_p4;

assign zext_ln708_87_fu_8857_p1 = tmp_171_fu_8847_p4;

assign zext_ln708_88_fu_8872_p1 = tmp_172_fu_8862_p4;

assign zext_ln708_89_fu_8887_p1 = tmp_173_fu_8877_p4;

assign zext_ln708_8_fu_4697_p1 = tmp_17_fu_4687_p4;

assign zext_ln708_90_fu_8902_p1 = tmp_174_fu_8892_p4;

assign zext_ln708_91_fu_8917_p1 = tmp_175_fu_8907_p4;

assign zext_ln708_92_fu_8932_p1 = tmp_176_fu_8922_p4;

assign zext_ln708_93_fu_8947_p1 = tmp_177_fu_8937_p4;

assign zext_ln708_94_fu_8962_p1 = tmp_178_fu_8952_p4;

assign zext_ln708_95_fu_8977_p1 = tmp_179_fu_8967_p4;

assign zext_ln708_96_fu_8992_p1 = tmp_180_fu_8982_p4;

assign zext_ln708_97_fu_9007_p1 = tmp_181_fu_8997_p4;

assign zext_ln708_98_fu_9022_p1 = tmp_182_fu_9012_p4;

assign zext_ln708_99_fu_9632_p1 = trunc_ln708_6_fu_9628_p1;

assign zext_ln708_9_fu_4712_p1 = tmp_18_fu_4702_p4;

assign zext_ln708_fu_4622_p1 = trunc_ln708_fu_4618_p1;

endmodule //testEnc_process_r
