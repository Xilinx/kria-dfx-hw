-- Copyright (C) 2022, Advanced Micro Devices, Inc. All rights reserved.
-- SPDX-License-Identifier: MIT

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity add_sub_mm is
generic (
    C_M_AXI_GMEM_ADDR_WIDTH : INTEGER := 64;
    C_M_AXI_GMEM_ID_WIDTH : INTEGER := 1;
    C_M_AXI_GMEM_AWUSER_WIDTH : INTEGER := 1;
    C_M_AXI_GMEM_DATA_WIDTH : INTEGER := 128;
    C_M_AXI_GMEM_WUSER_WIDTH : INTEGER := 1;
    C_M_AXI_GMEM_ARUSER_WIDTH : INTEGER := 1;
    C_M_AXI_GMEM_RUSER_WIDTH : INTEGER := 1;
    C_M_AXI_GMEM_BUSER_WIDTH : INTEGER := 1;
    C_S_AXI_CONTROL_ADDR_WIDTH : INTEGER := 7;
    C_S_AXI_CONTROL_DATA_WIDTH : INTEGER := 32;
    C_M_AXI_GMEM_USER_VALUE : INTEGER := 0;
    C_M_AXI_GMEM_PROT_VALUE : INTEGER := 0;
    C_M_AXI_GMEM_CACHE_VALUE : INTEGER := 3 );
port (
    ap_clk : IN STD_LOGIC;
    ap_rst_n : IN STD_LOGIC;
    m_axi_gmem_AWVALID : OUT STD_LOGIC;
    m_axi_gmem_AWREADY : IN STD_LOGIC;
    m_axi_gmem_AWADDR : OUT STD_LOGIC_VECTOR (C_M_AXI_GMEM_ADDR_WIDTH-1 downto 0);
    m_axi_gmem_AWID : OUT STD_LOGIC_VECTOR (C_M_AXI_GMEM_ID_WIDTH-1 downto 0);
    m_axi_gmem_AWLEN : OUT STD_LOGIC_VECTOR (7 downto 0);
    m_axi_gmem_AWSIZE : OUT STD_LOGIC_VECTOR (2 downto 0);
    m_axi_gmem_AWBURST : OUT STD_LOGIC_VECTOR (1 downto 0);
    m_axi_gmem_AWLOCK : OUT STD_LOGIC_VECTOR (1 downto 0);
    m_axi_gmem_AWCACHE : OUT STD_LOGIC_VECTOR (3 downto 0);
    m_axi_gmem_AWPROT : OUT STD_LOGIC_VECTOR (2 downto 0);
    m_axi_gmem_AWQOS : OUT STD_LOGIC_VECTOR (3 downto 0);
    m_axi_gmem_AWREGION : OUT STD_LOGIC_VECTOR (3 downto 0);
    m_axi_gmem_AWUSER : OUT STD_LOGIC_VECTOR (C_M_AXI_GMEM_AWUSER_WIDTH-1 downto 0);
    m_axi_gmem_WVALID : OUT STD_LOGIC;
    m_axi_gmem_WREADY : IN STD_LOGIC;
    m_axi_gmem_WDATA : OUT STD_LOGIC_VECTOR (C_M_AXI_GMEM_DATA_WIDTH-1 downto 0);
    m_axi_gmem_WSTRB : OUT STD_LOGIC_VECTOR (C_M_AXI_GMEM_DATA_WIDTH/8-1 downto 0);
    m_axi_gmem_WLAST : OUT STD_LOGIC;
    m_axi_gmem_WID : OUT STD_LOGIC_VECTOR (C_M_AXI_GMEM_ID_WIDTH-1 downto 0);
    m_axi_gmem_WUSER : OUT STD_LOGIC_VECTOR (C_M_AXI_GMEM_WUSER_WIDTH-1 downto 0);
    m_axi_gmem_ARVALID : OUT STD_LOGIC;
    m_axi_gmem_ARREADY : IN STD_LOGIC;
    m_axi_gmem_ARADDR : OUT STD_LOGIC_VECTOR (C_M_AXI_GMEM_ADDR_WIDTH-1 downto 0);
    m_axi_gmem_ARID : OUT STD_LOGIC_VECTOR (C_M_AXI_GMEM_ID_WIDTH-1 downto 0);
    m_axi_gmem_ARLEN : OUT STD_LOGIC_VECTOR (7 downto 0);
    m_axi_gmem_ARSIZE : OUT STD_LOGIC_VECTOR (2 downto 0);
    m_axi_gmem_ARBURST : OUT STD_LOGIC_VECTOR (1 downto 0);
    m_axi_gmem_ARLOCK : OUT STD_LOGIC_VECTOR (1 downto 0);
    m_axi_gmem_ARCACHE : OUT STD_LOGIC_VECTOR (3 downto 0);
    m_axi_gmem_ARPROT : OUT STD_LOGIC_VECTOR (2 downto 0);
    m_axi_gmem_ARQOS : OUT STD_LOGIC_VECTOR (3 downto 0);
    m_axi_gmem_ARREGION : OUT STD_LOGIC_VECTOR (3 downto 0);
    m_axi_gmem_ARUSER : OUT STD_LOGIC_VECTOR (C_M_AXI_GMEM_ARUSER_WIDTH-1 downto 0);
    m_axi_gmem_RVALID : IN STD_LOGIC;
    m_axi_gmem_RREADY : OUT STD_LOGIC;
    m_axi_gmem_RDATA : IN STD_LOGIC_VECTOR (C_M_AXI_GMEM_DATA_WIDTH-1 downto 0);
    m_axi_gmem_RLAST : IN STD_LOGIC;
    m_axi_gmem_RID : IN STD_LOGIC_VECTOR (C_M_AXI_GMEM_ID_WIDTH-1 downto 0);
    m_axi_gmem_RUSER : IN STD_LOGIC_VECTOR (C_M_AXI_GMEM_RUSER_WIDTH-1 downto 0);
    m_axi_gmem_RRESP : IN STD_LOGIC_VECTOR (1 downto 0);
    m_axi_gmem_BVALID : IN STD_LOGIC;
    m_axi_gmem_BREADY : OUT STD_LOGIC;
    m_axi_gmem_BRESP : IN STD_LOGIC_VECTOR (1 downto 0);
    m_axi_gmem_BID : IN STD_LOGIC_VECTOR (C_M_AXI_GMEM_ID_WIDTH-1 downto 0);
    m_axi_gmem_BUSER : IN STD_LOGIC_VECTOR (C_M_AXI_GMEM_BUSER_WIDTH-1 downto 0);
    s_axi_control_AWVALID : IN STD_LOGIC;
    s_axi_control_AWREADY : OUT STD_LOGIC;
    s_axi_control_AWADDR : IN STD_LOGIC_VECTOR (C_S_AXI_CONTROL_ADDR_WIDTH-1 downto 0);
    s_axi_control_WVALID : IN STD_LOGIC;
    s_axi_control_WREADY : OUT STD_LOGIC;
    s_axi_control_WDATA : IN STD_LOGIC_VECTOR (C_S_AXI_CONTROL_DATA_WIDTH-1 downto 0);
    s_axi_control_WSTRB : IN STD_LOGIC_VECTOR (C_S_AXI_CONTROL_DATA_WIDTH/8-1 downto 0);
    s_axi_control_ARVALID : IN STD_LOGIC;
    s_axi_control_ARREADY : OUT STD_LOGIC;
    s_axi_control_ARADDR : IN STD_LOGIC_VECTOR (C_S_AXI_CONTROL_ADDR_WIDTH-1 downto 0);
    s_axi_control_RVALID : OUT STD_LOGIC;
    s_axi_control_RREADY : IN STD_LOGIC;
    s_axi_control_RDATA : OUT STD_LOGIC_VECTOR (C_S_AXI_CONTROL_DATA_WIDTH-1 downto 0);
    s_axi_control_RRESP : OUT STD_LOGIC_VECTOR (1 downto 0);
    s_axi_control_BVALID : OUT STD_LOGIC;
    s_axi_control_BREADY : IN STD_LOGIC;
    s_axi_control_BRESP : OUT STD_LOGIC_VECTOR (1 downto 0);
    interrupt : OUT STD_LOGIC );
end;


architecture behav of add_sub_mm is 
    attribute CORE_GENERATION_INFO : STRING;
    attribute CORE_GENERATION_INFO of behav : architecture is
    "add_sub_mm_add_sub_mm,hls_ip_2022_1,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=0,HLS_INPUT_PART=xck26-sfvc784-2LV-c,HLS_INPUT_CLOCK=3.000000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=2.190000,HLS_SYN_LAT=-1,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=2638,HLS_SYN_LUT=3654,HLS_VERSION=2022_1}";
    constant ap_const_logic_1 : STD_LOGIC := '1';
    constant ap_const_logic_0 : STD_LOGIC := '0';
    constant ap_ST_fsm_state1 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000001";
    constant ap_ST_fsm_pp0_stage0 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
    constant ap_ST_fsm_pp0_stage1 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000100";
    constant ap_ST_fsm_pp0_stage2 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000001000";
    constant ap_ST_fsm_pp0_stage3 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000010000";
    constant ap_ST_fsm_pp0_stage4 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000100000";
    constant ap_ST_fsm_pp0_stage5 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000001000000";
    constant ap_ST_fsm_pp0_stage6 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000010000000";
    constant ap_ST_fsm_pp0_stage7 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000100000000";
    constant ap_ST_fsm_pp0_stage8 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000001000000000";
    constant ap_ST_fsm_pp0_stage9 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000010000000000";
    constant ap_ST_fsm_pp0_stage10 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000100000000000";
    constant ap_ST_fsm_pp0_stage11 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000001000000000000";
    constant ap_ST_fsm_pp0_stage12 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000010000000000000";
    constant ap_ST_fsm_pp0_stage13 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000100000000000000";
    constant ap_ST_fsm_pp0_stage14 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000001000000000000000";
    constant ap_ST_fsm_pp0_stage15 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000010000000000000000";
    constant ap_ST_fsm_pp0_stage16 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000100000000000000000";
    constant ap_ST_fsm_pp0_stage17 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000001000000000000000000";
    constant ap_ST_fsm_pp0_stage18 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000010000000000000000000";
    constant ap_ST_fsm_pp0_stage19 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000100000000000000000000";
    constant ap_ST_fsm_pp0_stage20 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000000000001000000000000000000000";
    constant ap_ST_fsm_pp0_stage21 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000000000010000000000000000000000";
    constant ap_ST_fsm_pp0_stage22 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000000000100000000000000000000000";
    constant ap_ST_fsm_pp0_stage23 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000000001000000000000000000000000";
    constant ap_ST_fsm_pp0_stage24 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000000010000000000000000000000000";
    constant ap_ST_fsm_pp0_stage25 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000000100000000000000000000000000";
    constant ap_ST_fsm_pp0_stage26 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000001000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage27 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000010000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage28 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000100000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage29 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000001000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage30 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000010000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage31 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000100000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage32 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000001000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage33 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000010000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage34 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000100000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage35 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000001000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage36 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000010000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage37 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000100000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage38 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000001000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage39 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000010000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage40 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000100000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage41 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000001000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage42 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000010000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage43 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000100000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage44 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000001000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage45 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000010000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage46 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000100000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage47 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000001000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage48 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000010000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage49 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000100000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage50 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000001000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage51 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000010000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage52 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000100000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage53 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000001000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage54 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000010000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage55 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000100000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage56 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000001000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage57 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000010000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage58 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000100000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage59 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000001000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage60 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000010000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage61 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000100000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage62 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000001000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage63 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000010000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage64 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000100000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage65 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000001000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage66 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000010000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage67 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage68 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000001000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage69 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000010000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage70 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000100000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage71 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000001000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage72 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000010000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage73 : STD_LOGIC_VECTOR (84 downto 0) := "0000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage74 : STD_LOGIC_VECTOR (84 downto 0) := "0000000001000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage75 : STD_LOGIC_VECTOR (84 downto 0) := "0000000010000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage76 : STD_LOGIC_VECTOR (84 downto 0) := "0000000100000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage77 : STD_LOGIC_VECTOR (84 downto 0) := "0000001000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage78 : STD_LOGIC_VECTOR (84 downto 0) := "0000010000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage79 : STD_LOGIC_VECTOR (84 downto 0) := "0000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage80 : STD_LOGIC_VECTOR (84 downto 0) := "0001000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage81 : STD_LOGIC_VECTOR (84 downto 0) := "0010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_pp0_stage82 : STD_LOGIC_VECTOR (84 downto 0) := "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state100 : STD_LOGIC_VECTOR (84 downto 0) := "1000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_const_lv32_0 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000000";
    constant ap_const_boolean_1 : BOOLEAN := true;
    constant ap_const_lv32_2 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000010";
    constant ap_const_boolean_0 : BOOLEAN := false;
    constant ap_const_lv1_1 : STD_LOGIC_VECTOR (0 downto 0) := "1";
    constant ap_const_lv32_9 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000001001";
    constant ap_const_lv32_33 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000110011";
    constant ap_const_lv32_3A : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000111010";
    constant ap_const_lv32_43 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000001000011";
    constant ap_const_lv32_4A : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000001001010";
    constant ap_const_lv32_53 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000001010011";
    constant ap_const_lv32_7 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000111";
    constant ap_const_lv32_12 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000010010";
    constant ap_const_lv1_0 : STD_LOGIC_VECTOR (0 downto 0) := "0";
    constant ap_const_lv32_19 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000011001";
    constant ap_const_lv32_22 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000100010";
    constant ap_const_lv32_29 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000101001";
    constant ap_const_lv32_32 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000110010";
    constant ap_const_lv32_39 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000111001";
    constant ap_const_lv32_3 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000011";
    constant ap_const_lv32_A : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000001010";
    constant ap_const_lv32_34 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000110100";
    constant ap_const_lv32_3B : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000111011";
    constant ap_const_lv32_44 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000001000100";
    constant ap_const_lv32_4B : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000001001011";
    constant ap_const_lv32_1 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000001";
    constant ap_const_lv32_8 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000001000";
    constant ap_const_lv32_13 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000010011";
    constant ap_const_lv32_1A : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000011010";
    constant ap_const_lv32_23 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000100011";
    constant ap_const_lv32_2A : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000101010";
    constant ap_const_lv32_2D : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000101101";
    constant ap_const_lv32_3D : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000111101";
    constant ap_const_lv32_42 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000001000010";
    constant ap_const_lv32_4 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000100";
    constant ap_const_lv32_4D : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000001001101";
    constant ap_const_lv32_52 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000001010010";
    constant ap_const_lv32_C : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000001100";
    constant ap_const_lv32_11 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000010001";
    constant ap_const_lv32_1C : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000011100";
    constant ap_const_lv32_21 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000100001";
    constant ap_const_lv32_2C : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000101100";
    constant ap_const_lv32_31 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000110001";
    constant ap_const_lv32_B : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000001011";
    constant ap_const_lv32_F : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000001111";
    constant ap_const_lv32_1B : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000011011";
    constant ap_const_lv32_2B : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000101011";
    constant ap_const_lv32_3C : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000111100";
    constant ap_const_lv32_4C : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000001001100";
    constant C_S_AXI_DATA_WIDTH : INTEGER range 63 downto 0 := 20;
    constant C_M_AXI_DATA_WIDTH : INTEGER range 63 downto 0 := 20;
    constant ap_const_lv4_0 : STD_LOGIC_VECTOR (3 downto 0) := "0000";
    constant ap_const_lv16_F : STD_LOGIC_VECTOR (15 downto 0) := "0000000000001111";
    constant ap_const_lv16_FFFF : STD_LOGIC_VECTOR (15 downto 0) := "1111111111111111";
    constant ap_const_lv32_20 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000100000";
    constant ap_const_lv32_3F : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000111111";
    constant ap_const_lv32_40 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000001000000";
    constant ap_const_lv32_5F : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000001011111";
    constant ap_const_lv32_60 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000001100000";
    constant ap_const_lv32_7F : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000001111111";
    constant ap_const_lv32_10 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000010000";
    constant ap_const_lv32_54 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000001010100";

    signal ap_rst_n_inv : STD_LOGIC;
    signal ap_start : STD_LOGIC;
    signal ap_done : STD_LOGIC;
    signal ap_idle : STD_LOGIC;
    signal ap_CS_fsm : STD_LOGIC_VECTOR (84 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000001";
    attribute fsm_encoding : string;
    attribute fsm_encoding of ap_CS_fsm : signal is "none";
    signal ap_CS_fsm_state1 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_state1 : signal is "none";
    signal ap_ready : STD_LOGIC;
    signal arg1 : STD_LOGIC_VECTOR (63 downto 0);
    signal arg2 : STD_LOGIC_VECTOR (63 downto 0);
    signal mem : STD_LOGIC_VECTOR (63 downto 0);
    signal src_addr1 : STD_LOGIC_VECTOR (31 downto 0);
    signal src_addr2 : STD_LOGIC_VECTOR (31 downto 0);
    signal dst_addr : STD_LOGIC_VECTOR (31 downto 0);
    signal size : STD_LOGIC_VECTOR (31 downto 0);
    signal op : STD_LOGIC_VECTOR (0 downto 0);
    signal gmem_blk_n_AR : STD_LOGIC;
    signal ap_CS_fsm_pp0_stage1 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage1 : signal is "none";
    signal ap_enable_reg_pp0_iter0 : STD_LOGIC := '0';
    signal ap_block_pp0_stage1 : BOOLEAN;
    signal icmp_ln1073_reg_676 : STD_LOGIC_VECTOR (0 downto 0);
    signal gmem_blk_n_R : STD_LOGIC;
    signal ap_CS_fsm_pp0_stage8 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage8 : signal is "none";
    signal ap_block_pp0_stage8 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage50 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage50 : signal is "none";
    signal ap_block_pp0_stage50 : BOOLEAN;
    signal op_read_reg_640 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_CS_fsm_pp0_stage57 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage57 : signal is "none";
    signal ap_block_pp0_stage57 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage66 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage66 : signal is "none";
    signal ap_block_pp0_stage66 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage73 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage73 : signal is "none";
    signal ap_block_pp0_stage73 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage82 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage82 : signal is "none";
    signal ap_block_pp0_stage82 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage6 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage6 : signal is "none";
    signal ap_enable_reg_pp0_iter1 : STD_LOGIC := '0';
    signal ap_block_pp0_stage6 : BOOLEAN;
    signal icmp_ln1073_reg_676_pp0_iter1_reg : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_CS_fsm_pp0_stage17 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage17 : signal is "none";
    signal ap_block_pp0_stage17 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage24 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage24 : signal is "none";
    signal ap_block_pp0_stage24 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage33 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage33 : signal is "none";
    signal ap_block_pp0_stage33 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage40 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage40 : signal is "none";
    signal ap_block_pp0_stage40 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage49 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage49 : signal is "none";
    signal ap_block_pp0_stage49 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage56 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage56 : signal is "none";
    signal ap_block_pp0_stage56 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage2 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage2 : signal is "none";
    signal ap_block_pp0_stage2 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage9 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage9 : signal is "none";
    signal ap_block_pp0_stage9 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage51 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage51 : signal is "none";
    signal ap_block_pp0_stage51 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage58 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage58 : signal is "none";
    signal ap_block_pp0_stage58 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage67 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage67 : signal is "none";
    signal ap_block_pp0_stage67 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage74 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage74 : signal is "none";
    signal ap_block_pp0_stage74 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage0 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage0 : signal is "none";
    signal ap_block_pp0_stage0 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage7 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage7 : signal is "none";
    signal ap_block_pp0_stage7 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage18 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage18 : signal is "none";
    signal ap_block_pp0_stage18 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage25 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage25 : signal is "none";
    signal ap_block_pp0_stage25 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage34 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage34 : signal is "none";
    signal ap_block_pp0_stage34 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage41 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage41 : signal is "none";
    signal ap_block_pp0_stage41 : BOOLEAN;
    signal gmem_blk_n_AW : STD_LOGIC;
    signal gmem_blk_n_W : STD_LOGIC;
    signal ap_CS_fsm_pp0_stage44 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage44 : signal is "none";
    signal ap_block_pp0_stage44 : BOOLEAN;
    signal gmem_blk_n_B : STD_LOGIC;
    signal ap_CS_fsm_pp0_stage60 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage60 : signal is "none";
    signal ap_block_pp0_stage60 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage65 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage65 : signal is "none";
    signal ap_block_pp0_stage65 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage3 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage3 : signal is "none";
    signal ap_block_pp0_stage3 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage76 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage76 : signal is "none";
    signal ap_block_pp0_stage76 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage81 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage81 : signal is "none";
    signal ap_block_pp0_stage81 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage11 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage11 : signal is "none";
    signal ap_block_pp0_stage11 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage16 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage16 : signal is "none";
    signal ap_block_pp0_stage16 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage27 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage27 : signal is "none";
    signal ap_block_pp0_stage27 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage32 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage32 : signal is "none";
    signal ap_block_pp0_stage32 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage43 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage43 : signal is "none";
    signal ap_block_pp0_stage43 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage48 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage48 : signal is "none";
    signal ap_block_pp0_stage48 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage10 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage10 : signal is "none";
    signal ap_block_pp0_stage10 : BOOLEAN;
    signal ap_CS_fsm_pp0_stage14 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage14 : signal is "none";
    signal ap_block_pp0_stage14 : BOOLEAN;
    signal reg_320 : STD_LOGIC_VECTOR (31 downto 0);
    signal gmem_AWVALID : STD_LOGIC;
    signal gmem_AWREADY : STD_LOGIC;
    signal gmem_AWADDR : STD_LOGIC_VECTOR (63 downto 0);
    signal gmem_WVALID : STD_LOGIC;
    signal gmem_WREADY : STD_LOGIC;
    signal gmem_WDATA : STD_LOGIC_VECTOR (127 downto 0);
    signal gmem_WSTRB : STD_LOGIC_VECTOR (15 downto 0);
    signal gmem_ARVALID : STD_LOGIC;
    signal gmem_ARREADY : STD_LOGIC;
    signal gmem_ARADDR : STD_LOGIC_VECTOR (63 downto 0);
    signal gmem_RVALID : STD_LOGIC;
    signal gmem_RREADY : STD_LOGIC;
    signal gmem_RDATA : STD_LOGIC_VECTOR (127 downto 0);
    signal gmem_RFIFONUM : STD_LOGIC_VECTOR (8 downto 0);
    signal gmem_BVALID : STD_LOGIC;
    signal gmem_BREADY : STD_LOGIC;
    signal ap_predicate_op213_read_state26 : BOOLEAN;
    signal ap_block_state26_pp0_stage24_iter0 : BOOLEAN;
    signal ap_block_pp0_stage24_11001 : BOOLEAN;
    signal ap_predicate_op290_read_state59 : BOOLEAN;
    signal ap_predicate_op292_read_state59 : BOOLEAN;
    signal ap_block_state59_pp0_stage57_iter0 : BOOLEAN;
    signal ap_block_pp0_stage57_11001 : BOOLEAN;
    signal reg_324 : STD_LOGIC_VECTOR (31 downto 0);
    signal ap_predicate_op216_read_state27 : BOOLEAN;
    signal ap_block_state27_pp0_stage25_iter0 : BOOLEAN;
    signal ap_block_pp0_stage25_11001 : BOOLEAN;
    signal ap_predicate_op298_read_state60 : BOOLEAN;
    signal ap_block_state60_pp0_stage58_iter0 : BOOLEAN;
    signal ap_block_pp0_stage58_11001 : BOOLEAN;
    signal reg_328 : STD_LOGIC_VECTOR (31 downto 0);
    signal ap_predicate_op240_read_state42 : BOOLEAN;
    signal ap_block_state42_pp0_stage40_iter0 : BOOLEAN;
    signal ap_block_pp0_stage40_11001 : BOOLEAN;
    signal ap_predicate_op322_read_state75 : BOOLEAN;
    signal ap_block_state75_pp0_stage73_iter0 : BOOLEAN;
    signal ap_block_pp0_stage73_11001 : BOOLEAN;
    signal reg_332 : STD_LOGIC_VECTOR (31 downto 0);
    signal ap_predicate_op243_read_state43 : BOOLEAN;
    signal ap_block_state43_pp0_stage41_iter0 : BOOLEAN;
    signal ap_block_pp0_stage41_11001 : BOOLEAN;
    signal ap_predicate_op325_read_state76 : BOOLEAN;
    signal ap_block_state76_pp0_stage74_iter0 : BOOLEAN;
    signal ap_block_pp0_stage74_11001 : BOOLEAN;
    signal reg_336 : STD_LOGIC_VECTOR (31 downto 0);
    signal ap_predicate_op285_read_state58 : BOOLEAN;
    signal ap_block_state58_pp0_stage56_iter0 : BOOLEAN;
    signal ap_block_pp0_stage56_11001 : BOOLEAN;
    signal ap_block_state8_pp0_stage6_iter0 : BOOLEAN;
    signal ap_predicate_op351_read_state91 : BOOLEAN;
    signal ap_block_state91_pp0_stage6_iter1 : BOOLEAN;
    signal ap_block_pp0_stage6_11001 : BOOLEAN;
    signal reg_340 : STD_LOGIC_VECTOR (31 downto 0);
    signal ap_block_state9_pp0_stage7_iter0 : BOOLEAN;
    signal ap_predicate_op354_read_state92 : BOOLEAN;
    signal ap_block_state92_pp0_stage7_iter1 : BOOLEAN;
    signal ap_block_pp0_stage7_11001 : BOOLEAN;
    signal size_read_reg_644 : STD_LOGIC_VECTOR (31 downto 0);
    signal mem_read_reg_649 : STD_LOGIC_VECTOR (63 downto 0);
    signal lhs_fu_344_p1 : STD_LOGIC_VECTOR (33 downto 0);
    signal lhs_reg_656 : STD_LOGIC_VECTOR (33 downto 0);
    signal lhs_5_fu_348_p1 : STD_LOGIC_VECTOR (33 downto 0);
    signal lhs_5_reg_661 : STD_LOGIC_VECTOR (33 downto 0);
    signal lhs_6_fu_352_p1 : STD_LOGIC_VECTOR (33 downto 0);
    signal lhs_6_reg_666 : STD_LOGIC_VECTOR (33 downto 0);
    signal i_V_2_reg_671 : STD_LOGIC_VECTOR (31 downto 0);
    signal ap_block_state2_pp0_stage0_iter0 : BOOLEAN;
    signal ap_block_state85_pp0_stage0_iter1 : BOOLEAN;
    signal ap_predicate_op340_readreq_state85 : BOOLEAN;
    signal ap_block_state85_io : BOOLEAN;
    signal ap_block_pp0_stage0_11001 : BOOLEAN;
    signal icmp_ln1073_fu_364_p2 : STD_LOGIC_VECTOR (0 downto 0);
    signal trunc_ln_reg_680 : STD_LOGIC_VECTOR (59 downto 0);
    signal trunc_ln357_1_reg_685 : STD_LOGIC_VECTOR (59 downto 0);
    signal trunc_ln1_reg_690 : STD_LOGIC_VECTOR (59 downto 0);
    signal gmem_addr_reg_695 : STD_LOGIC_VECTOR (63 downto 0);
    signal ap_block_state3_pp0_stage1_iter0 : BOOLEAN;
    signal ap_predicate_op164_writereq_state3 : BOOLEAN;
    signal ap_predicate_op165_writereq_state3 : BOOLEAN;
    signal ap_block_state3_io : BOOLEAN;
    signal ap_block_state86_pp0_stage1_iter1 : BOOLEAN;
    signal ap_block_pp0_stage1_11001 : BOOLEAN;
    signal gmem_addr_2_reg_701 : STD_LOGIC_VECTOR (63 downto 0);
    signal gmem_addr_1_reg_713 : STD_LOGIC_VECTOR (63 downto 0);
    signal ap_block_state4_pp0_stage2_iter0 : BOOLEAN;
    signal ap_predicate_op170_writereq_state4 : BOOLEAN;
    signal ap_predicate_op171_writereq_state4 : BOOLEAN;
    signal ap_block_state4_io : BOOLEAN;
    signal ap_block_state87_pp0_stage2_iter1 : BOOLEAN;
    signal ap_block_pp0_stage2_11001 : BOOLEAN;
    signal trunc_ln357_fu_499_p1 : STD_LOGIC_VECTOR (31 downto 0);
    signal trunc_ln357_reg_719 : STD_LOGIC_VECTOR (31 downto 0);
    signal ap_block_state10_pp0_stage8_iter0 : BOOLEAN;
    signal ap_block_state93_pp0_stage8_iter1 : BOOLEAN;
    signal ap_block_pp0_stage8_11001 : BOOLEAN;
    signal trunc_ln357_2_fu_503_p1 : STD_LOGIC_VECTOR (31 downto 0);
    signal trunc_ln357_2_reg_725 : STD_LOGIC_VECTOR (31 downto 0);
    signal ap_block_state11_pp0_stage9_iter0 : BOOLEAN;
    signal ap_block_state94_pp0_stage9_iter1 : BOOLEAN;
    signal ap_block_pp0_stage9_11001 : BOOLEAN;
    signal sub_ln414_fu_507_p2 : STD_LOGIC_VECTOR (31 downto 0);
    signal sub_ln414_reg_731 : STD_LOGIC_VECTOR (31 downto 0);
    signal ap_block_state12_pp0_stage10_iter0 : BOOLEAN;
    signal ap_block_state12_io : BOOLEAN;
    signal ap_block_state95_pp0_stage10_iter1 : BOOLEAN;
    signal ap_block_pp0_stage10_11001 : BOOLEAN;
    signal add_ln414_1_fu_511_p2 : STD_LOGIC_VECTOR (31 downto 0);
    signal add_ln414_1_reg_739 : STD_LOGIC_VECTOR (31 downto 0);
    signal sub_ln414_1_fu_519_p2 : STD_LOGIC_VECTOR (31 downto 0);
    signal sub_ln414_1_reg_747 : STD_LOGIC_VECTOR (31 downto 0);
    signal ap_CS_fsm_pp0_stage26 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage26 : signal is "none";
    signal ap_block_state28_pp0_stage26_iter0 : BOOLEAN;
    signal ap_block_pp0_stage26_11001 : BOOLEAN;
    signal sub_ln414_2_fu_536_p2 : STD_LOGIC_VECTOR (31 downto 0);
    signal sub_ln414_2_reg_754 : STD_LOGIC_VECTOR (31 downto 0);
    signal ap_CS_fsm_pp0_stage42 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage42 : signal is "none";
    signal ap_block_state44_pp0_stage42_iter0 : BOOLEAN;
    signal ap_block_pp0_stage42_11001 : BOOLEAN;
    signal p_Result_4_fu_564_p5 : STD_LOGIC_VECTOR (127 downto 0);
    signal add_ln414_2_fu_573_p2 : STD_LOGIC_VECTOR (31 downto 0);
    signal add_ln414_2_reg_765 : STD_LOGIC_VECTOR (31 downto 0);
    signal ap_CS_fsm_pp0_stage59 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage59 : signal is "none";
    signal ap_block_state61_pp0_stage59_iter0 : BOOLEAN;
    signal ap_block_pp0_stage59_11001 : BOOLEAN;
    signal add_ln414_3_fu_590_p2 : STD_LOGIC_VECTOR (31 downto 0);
    signal add_ln414_3_reg_772 : STD_LOGIC_VECTOR (31 downto 0);
    signal ap_CS_fsm_pp0_stage75 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_pp0_stage75 : signal is "none";
    signal ap_block_state77_pp0_stage75_iter0 : BOOLEAN;
    signal ap_block_pp0_stage75_11001 : BOOLEAN;
    signal p_Result_s_fu_624_p5 : STD_LOGIC_VECTOR (127 downto 0);
    signal ap_block_pp0_stage0_subdone : BOOLEAN;
    signal ap_condition_pp0_exit_iter0_state2 : STD_LOGIC;
    signal ap_block_state84_pp0_stage82_iter0 : BOOLEAN;
    signal ap_predicate_op336_readreq_state84 : BOOLEAN;
    signal ap_block_state84_io : BOOLEAN;
    signal ap_block_pp0_stage82_subdone : BOOLEAN;
    signal ap_block_state16_pp0_stage14_iter0 : BOOLEAN;
    signal ap_block_state99_pp0_stage14_iter1 : BOOLEAN;
    signal ap_block_pp0_stage14_subdone : BOOLEAN;
    signal ap_phi_reg_pp0_iter0_storemerge_reg_250 : STD_LOGIC_VECTOR (127 downto 0);
    signal ap_phi_reg_pp0_iter1_storemerge_reg_250 : STD_LOGIC_VECTOR (127 downto 0);
    signal ap_block_pp0_stage82_11001 : BOOLEAN;
    signal sext_ln357_fu_469_p1 : STD_LOGIC_VECTOR (63 downto 0);
    signal sext_ln414_fu_479_p1 : STD_LOGIC_VECTOR (63 downto 0);
    signal sext_ln357_1_fu_489_p1 : STD_LOGIC_VECTOR (63 downto 0);
    signal ap_block_state19_pp0_stage17_iter0 : BOOLEAN;
    signal ap_predicate_op200_readreq_state19 : BOOLEAN;
    signal ap_block_state19_io : BOOLEAN;
    signal ap_block_pp0_stage17_11001 : BOOLEAN;
    signal ap_block_state35_pp0_stage33_iter0 : BOOLEAN;
    signal ap_predicate_op227_readreq_state35 : BOOLEAN;
    signal ap_block_state35_io : BOOLEAN;
    signal ap_block_pp0_stage33_11001 : BOOLEAN;
    signal ap_predicate_op261_writeresp_state51 : BOOLEAN;
    signal ap_block_state51_pp0_stage49_iter0 : BOOLEAN;
    signal ap_predicate_op260_readreq_state51 : BOOLEAN;
    signal ap_block_state51_io : BOOLEAN;
    signal ap_block_pp0_stage49_11001 : BOOLEAN;
    signal ap_block_state52_pp0_stage50_iter0 : BOOLEAN;
    signal ap_predicate_op263_readreq_state52 : BOOLEAN;
    signal ap_predicate_op264_readreq_state52 : BOOLEAN;
    signal ap_block_state52_io : BOOLEAN;
    signal ap_block_pp0_stage50_11001 : BOOLEAN;
    signal ap_block_state68_pp0_stage66_iter0 : BOOLEAN;
    signal ap_predicate_op309_readreq_state68 : BOOLEAN;
    signal ap_block_state68_io : BOOLEAN;
    signal ap_block_pp0_stage66_11001 : BOOLEAN;
    signal ap_block_state5_pp0_stage3_iter0 : BOOLEAN;
    signal ap_predicate_op174_writereq_state5 : BOOLEAN;
    signal ap_predicate_op175_writereq_state5 : BOOLEAN;
    signal ap_block_state5_io : BOOLEAN;
    signal ap_block_state88_pp0_stage3_iter1 : BOOLEAN;
    signal ap_block_pp0_stage3_11001 : BOOLEAN;
    signal ap_predicate_op199_writeresp_state18 : BOOLEAN;
    signal ap_block_state18_pp0_stage16_iter0 : BOOLEAN;
    signal ap_block_pp0_stage16_11001 : BOOLEAN;
    signal ap_predicate_op226_writeresp_state34 : BOOLEAN;
    signal ap_block_state34_pp0_stage32_iter0 : BOOLEAN;
    signal ap_block_pp0_stage32_11001 : BOOLEAN;
    signal ap_predicate_op258_writeresp_state50 : BOOLEAN;
    signal ap_block_state50_pp0_stage48_iter0 : BOOLEAN;
    signal ap_block_pp0_stage48_11001 : BOOLEAN;
    signal ap_predicate_op308_writeresp_state67 : BOOLEAN;
    signal ap_block_state67_pp0_stage65_iter0 : BOOLEAN;
    signal ap_block_pp0_stage65_11001 : BOOLEAN;
    signal ap_predicate_op335_writeresp_state83 : BOOLEAN;
    signal ap_block_state83_pp0_stage81_iter0 : BOOLEAN;
    signal ap_block_pp0_stage81_11001 : BOOLEAN;
    signal ap_block_pp0_stage14_11001 : BOOLEAN;
    signal ap_block_state20_pp0_stage18_iter0 : BOOLEAN;
    signal ap_predicate_op202_readreq_state20 : BOOLEAN;
    signal ap_block_state20_io : BOOLEAN;
    signal ap_block_pp0_stage18_11001 : BOOLEAN;
    signal ap_block_state36_pp0_stage34_iter0 : BOOLEAN;
    signal ap_predicate_op229_readreq_state36 : BOOLEAN;
    signal ap_block_state36_io : BOOLEAN;
    signal ap_block_pp0_stage34_11001 : BOOLEAN;
    signal ap_block_state53_pp0_stage51_iter0 : BOOLEAN;
    signal ap_predicate_op268_readreq_state53 : BOOLEAN;
    signal ap_block_state53_io : BOOLEAN;
    signal ap_block_pp0_stage51_11001 : BOOLEAN;
    signal ap_block_state69_pp0_stage67_iter0 : BOOLEAN;
    signal ap_predicate_op311_readreq_state69 : BOOLEAN;
    signal ap_block_state69_io : BOOLEAN;
    signal ap_block_pp0_stage67_11001 : BOOLEAN;
    signal ap_block_state13_pp0_stage11_iter0 : BOOLEAN;
    signal ap_predicate_op194_write_state13 : BOOLEAN;
    signal ap_block_state13_io : BOOLEAN;
    signal ap_block_state96_pp0_stage11_iter1 : BOOLEAN;
    signal ap_block_pp0_stage11_11001 : BOOLEAN;
    signal p_Result_11_fu_515_p1 : STD_LOGIC_VECTOR (127 downto 0);
    signal ap_block_pp0_stage11_01001 : BOOLEAN;
    signal ap_block_state29_pp0_stage27_iter0 : BOOLEAN;
    signal ap_predicate_op221_write_state29 : BOOLEAN;
    signal ap_block_state29_io : BOOLEAN;
    signal ap_block_pp0_stage27_11001 : BOOLEAN;
    signal p_Result_12_fu_531_p1 : STD_LOGIC_VECTOR (127 downto 0);
    signal ap_block_pp0_stage27_01001 : BOOLEAN;
    signal ap_block_state45_pp0_stage43_iter0 : BOOLEAN;
    signal ap_predicate_op248_write_state45 : BOOLEAN;
    signal ap_block_state45_io : BOOLEAN;
    signal ap_block_pp0_stage43_11001 : BOOLEAN;
    signal p_Result_13_fu_549_p1 : STD_LOGIC_VECTOR (127 downto 0);
    signal ap_block_pp0_stage43_01001 : BOOLEAN;
    signal ap_block_state46_pp0_stage44_iter0 : BOOLEAN;
    signal ap_predicate_op251_write_state46 : BOOLEAN;
    signal ap_block_state46_io : BOOLEAN;
    signal ap_block_pp0_stage44_11001 : BOOLEAN;
    signal p_Result_8_fu_554_p1 : STD_LOGIC_VECTOR (127 downto 0);
    signal ap_block_pp0_stage44_01001 : BOOLEAN;
    signal ap_block_state62_pp0_stage60_iter0 : BOOLEAN;
    signal ap_predicate_op303_write_state62 : BOOLEAN;
    signal ap_block_state62_io : BOOLEAN;
    signal ap_block_pp0_stage60_11001 : BOOLEAN;
    signal p_Result_9_fu_585_p1 : STD_LOGIC_VECTOR (127 downto 0);
    signal ap_block_pp0_stage60_01001 : BOOLEAN;
    signal ap_block_state78_pp0_stage76_iter0 : BOOLEAN;
    signal ap_predicate_op330_write_state78 : BOOLEAN;
    signal ap_block_state78_io : BOOLEAN;
    signal ap_block_pp0_stage76_11001 : BOOLEAN;
    signal p_Result_10_fu_603_p1 : STD_LOGIC_VECTOR (127 downto 0);
    signal ap_block_pp0_stage76_01001 : BOOLEAN;
    signal ap_block_pp0_stage9_01001 : BOOLEAN;
    signal rhs_V_fu_122 : STD_LOGIC_VECTOR (31 downto 0);
    signal i_V_fu_608_p2 : STD_LOGIC_VECTOR (31 downto 0);
    signal icmp_ln1073_fu_364_p0 : STD_LOGIC_VECTOR (31 downto 0);
    signal sext_ln232_fu_369_p0 : STD_LOGIC_VECTOR (31 downto 0);
    signal sext_ln232_fu_369_p1 : STD_LOGIC_VECTOR (33 downto 0);
    signal ret_V_fu_373_p2 : STD_LOGIC_VECTOR (33 downto 0);
    signal shl_ln_fu_383_p3 : STD_LOGIC_VECTOR (37 downto 0);
    signal sext_ln357_2_fu_391_p1 : STD_LOGIC_VECTOR (63 downto 0);
    signal ret_V_1_fu_378_p2 : STD_LOGIC_VECTOR (33 downto 0);
    signal shl_ln357_1_fu_400_p3 : STD_LOGIC_VECTOR (37 downto 0);
    signal sext_ln357_3_fu_408_p1 : STD_LOGIC_VECTOR (63 downto 0);
    signal ret_V_2_fu_417_p2 : STD_LOGIC_VECTOR (33 downto 0);
    signal shl_ln1_fu_422_p3 : STD_LOGIC_VECTOR (37 downto 0);
    signal sext_ln414_1_fu_430_p1 : STD_LOGIC_VECTOR (63 downto 0);
    signal add_ln357_fu_395_p2 : STD_LOGIC_VECTOR (63 downto 0);
    signal add_ln357_1_fu_412_p2 : STD_LOGIC_VECTOR (63 downto 0);
    signal add_ln414_fu_434_p2 : STD_LOGIC_VECTOR (63 downto 0);
    signal ap_block_pp0_stage26 : BOOLEAN;
    signal tmp_9_fu_525_p3 : STD_LOGIC_VECTOR (63 downto 0);
    signal ap_block_pp0_stage42 : BOOLEAN;
    signal tmp_12_fu_542_p4 : STD_LOGIC_VECTOR (95 downto 0);
    signal sub_ln414_3_fu_558_p2 : STD_LOGIC_VECTOR (31 downto 0);
    signal ap_block_pp0_stage59 : BOOLEAN;
    signal tmp_fu_579_p3 : STD_LOGIC_VECTOR (63 downto 0);
    signal ap_block_pp0_stage75 : BOOLEAN;
    signal tmp_4_fu_596_p4 : STD_LOGIC_VECTOR (95 downto 0);
    signal add_ln414_4_fu_618_p2 : STD_LOGIC_VECTOR (31 downto 0);
    signal ap_CS_fsm_state100 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_state100 : signal is "none";
    signal ap_NS_fsm : STD_LOGIC_VECTOR (84 downto 0);
    signal ap_ST_fsm_state1_blk : STD_LOGIC;
    signal ap_ST_fsm_state100_blk : STD_LOGIC;
    signal ap_block_pp0_stage1_subdone : BOOLEAN;
    signal ap_block_pp0_stage2_subdone : BOOLEAN;
    signal ap_block_pp0_stage3_subdone : BOOLEAN;
    signal ap_block_state6_pp0_stage4_iter0 : BOOLEAN;
    signal ap_block_state89_pp0_stage4_iter1 : BOOLEAN;
    signal ap_block_pp0_stage4_subdone : BOOLEAN;
    signal ap_block_pp0_stage4_11001 : BOOLEAN;
    signal ap_block_state7_pp0_stage5_iter0 : BOOLEAN;
    signal ap_block_state90_pp0_stage5_iter1 : BOOLEAN;
    signal ap_block_pp0_stage5_subdone : BOOLEAN;
    signal ap_block_pp0_stage5_11001 : BOOLEAN;
    signal ap_block_pp0_stage6_subdone : BOOLEAN;
    signal ap_block_pp0_stage7_subdone : BOOLEAN;
    signal ap_block_pp0_stage8_subdone : BOOLEAN;
    signal ap_block_pp0_stage9_subdone : BOOLEAN;
    signal ap_block_pp0_stage10_subdone : BOOLEAN;
    signal ap_block_pp0_stage11_subdone : BOOLEAN;
    signal ap_block_state14_pp0_stage12_iter0 : BOOLEAN;
    signal ap_block_state97_pp0_stage12_iter1 : BOOLEAN;
    signal ap_block_pp0_stage12_subdone : BOOLEAN;
    signal ap_block_pp0_stage12_11001 : BOOLEAN;
    signal ap_block_state15_pp0_stage13_iter0 : BOOLEAN;
    signal ap_block_state98_pp0_stage13_iter1 : BOOLEAN;
    signal ap_block_pp0_stage13_subdone : BOOLEAN;
    signal ap_block_pp0_stage13_11001 : BOOLEAN;
    signal ap_block_state17_pp0_stage15_iter0 : BOOLEAN;
    signal ap_block_pp0_stage15_subdone : BOOLEAN;
    signal ap_block_pp0_stage15_11001 : BOOLEAN;
    signal ap_block_pp0_stage16_subdone : BOOLEAN;
    signal ap_block_pp0_stage17_subdone : BOOLEAN;
    signal ap_block_pp0_stage18_subdone : BOOLEAN;
    signal ap_block_state21_pp0_stage19_iter0 : BOOLEAN;
    signal ap_block_pp0_stage19_subdone : BOOLEAN;
    signal ap_block_pp0_stage19_11001 : BOOLEAN;
    signal ap_block_state22_pp0_stage20_iter0 : BOOLEAN;
    signal ap_block_pp0_stage20_subdone : BOOLEAN;
    signal ap_block_pp0_stage20_11001 : BOOLEAN;
    signal ap_block_state23_pp0_stage21_iter0 : BOOLEAN;
    signal ap_block_pp0_stage21_subdone : BOOLEAN;
    signal ap_block_pp0_stage21_11001 : BOOLEAN;
    signal ap_block_state24_pp0_stage22_iter0 : BOOLEAN;
    signal ap_block_pp0_stage22_subdone : BOOLEAN;
    signal ap_block_pp0_stage22_11001 : BOOLEAN;
    signal ap_block_state25_pp0_stage23_iter0 : BOOLEAN;
    signal ap_block_pp0_stage23_subdone : BOOLEAN;
    signal ap_block_pp0_stage23_11001 : BOOLEAN;
    signal ap_block_pp0_stage24_subdone : BOOLEAN;
    signal ap_block_pp0_stage25_subdone : BOOLEAN;
    signal ap_block_pp0_stage26_subdone : BOOLEAN;
    signal ap_block_pp0_stage27_subdone : BOOLEAN;
    signal ap_block_state30_pp0_stage28_iter0 : BOOLEAN;
    signal ap_block_pp0_stage28_subdone : BOOLEAN;
    signal ap_block_pp0_stage28_11001 : BOOLEAN;
    signal ap_block_state31_pp0_stage29_iter0 : BOOLEAN;
    signal ap_block_pp0_stage29_subdone : BOOLEAN;
    signal ap_block_pp0_stage29_11001 : BOOLEAN;
    signal ap_block_state32_pp0_stage30_iter0 : BOOLEAN;
    signal ap_block_pp0_stage30_subdone : BOOLEAN;
    signal ap_block_pp0_stage30_11001 : BOOLEAN;
    signal ap_block_state33_pp0_stage31_iter0 : BOOLEAN;
    signal ap_block_pp0_stage31_subdone : BOOLEAN;
    signal ap_block_pp0_stage31_11001 : BOOLEAN;
    signal ap_block_pp0_stage32_subdone : BOOLEAN;
    signal ap_block_pp0_stage33_subdone : BOOLEAN;
    signal ap_block_pp0_stage34_subdone : BOOLEAN;
    signal ap_block_state37_pp0_stage35_iter0 : BOOLEAN;
    signal ap_block_pp0_stage35_subdone : BOOLEAN;
    signal ap_block_pp0_stage35_11001 : BOOLEAN;
    signal ap_block_state38_pp0_stage36_iter0 : BOOLEAN;
    signal ap_block_pp0_stage36_subdone : BOOLEAN;
    signal ap_block_pp0_stage36_11001 : BOOLEAN;
    signal ap_block_state39_pp0_stage37_iter0 : BOOLEAN;
    signal ap_block_pp0_stage37_subdone : BOOLEAN;
    signal ap_block_pp0_stage37_11001 : BOOLEAN;
    signal ap_block_state40_pp0_stage38_iter0 : BOOLEAN;
    signal ap_block_pp0_stage38_subdone : BOOLEAN;
    signal ap_block_pp0_stage38_11001 : BOOLEAN;
    signal ap_block_state41_pp0_stage39_iter0 : BOOLEAN;
    signal ap_block_pp0_stage39_subdone : BOOLEAN;
    signal ap_block_pp0_stage39_11001 : BOOLEAN;
    signal ap_block_pp0_stage40_subdone : BOOLEAN;
    signal ap_block_pp0_stage41_subdone : BOOLEAN;
    signal ap_block_pp0_stage42_subdone : BOOLEAN;
    signal ap_block_pp0_stage43_subdone : BOOLEAN;
    signal ap_block_pp0_stage44_subdone : BOOLEAN;
    signal ap_block_state47_pp0_stage45_iter0 : BOOLEAN;
    signal ap_block_pp0_stage45_subdone : BOOLEAN;
    signal ap_block_pp0_stage45_11001 : BOOLEAN;
    signal ap_block_state48_pp0_stage46_iter0 : BOOLEAN;
    signal ap_block_pp0_stage46_subdone : BOOLEAN;
    signal ap_block_pp0_stage46_11001 : BOOLEAN;
    signal ap_block_state49_pp0_stage47_iter0 : BOOLEAN;
    signal ap_block_pp0_stage47_subdone : BOOLEAN;
    signal ap_block_pp0_stage47_11001 : BOOLEAN;
    signal ap_block_pp0_stage48_subdone : BOOLEAN;
    signal ap_block_pp0_stage49_subdone : BOOLEAN;
    signal ap_block_pp0_stage50_subdone : BOOLEAN;
    signal ap_block_pp0_stage51_subdone : BOOLEAN;
    signal ap_block_state54_pp0_stage52_iter0 : BOOLEAN;
    signal ap_block_pp0_stage52_subdone : BOOLEAN;
    signal ap_block_pp0_stage52_11001 : BOOLEAN;
    signal ap_block_state55_pp0_stage53_iter0 : BOOLEAN;
    signal ap_block_pp0_stage53_subdone : BOOLEAN;
    signal ap_block_pp0_stage53_11001 : BOOLEAN;
    signal ap_block_state56_pp0_stage54_iter0 : BOOLEAN;
    signal ap_block_pp0_stage54_subdone : BOOLEAN;
    signal ap_block_pp0_stage54_11001 : BOOLEAN;
    signal ap_block_state57_pp0_stage55_iter0 : BOOLEAN;
    signal ap_block_pp0_stage55_subdone : BOOLEAN;
    signal ap_block_pp0_stage55_11001 : BOOLEAN;
    signal ap_block_pp0_stage56_subdone : BOOLEAN;
    signal ap_block_pp0_stage57_subdone : BOOLEAN;
    signal ap_block_pp0_stage58_subdone : BOOLEAN;
    signal ap_block_pp0_stage59_subdone : BOOLEAN;
    signal ap_block_pp0_stage60_subdone : BOOLEAN;
    signal ap_block_state63_pp0_stage61_iter0 : BOOLEAN;
    signal ap_block_pp0_stage61_subdone : BOOLEAN;
    signal ap_block_pp0_stage61_11001 : BOOLEAN;
    signal ap_block_state64_pp0_stage62_iter0 : BOOLEAN;
    signal ap_block_pp0_stage62_subdone : BOOLEAN;
    signal ap_block_pp0_stage62_11001 : BOOLEAN;
    signal ap_block_state65_pp0_stage63_iter0 : BOOLEAN;
    signal ap_block_pp0_stage63_subdone : BOOLEAN;
    signal ap_block_pp0_stage63_11001 : BOOLEAN;
    signal ap_block_state66_pp0_stage64_iter0 : BOOLEAN;
    signal ap_block_pp0_stage64_subdone : BOOLEAN;
    signal ap_block_pp0_stage64_11001 : BOOLEAN;
    signal ap_block_pp0_stage65_subdone : BOOLEAN;
    signal ap_block_pp0_stage66_subdone : BOOLEAN;
    signal ap_block_pp0_stage67_subdone : BOOLEAN;
    signal ap_block_state70_pp0_stage68_iter0 : BOOLEAN;
    signal ap_block_pp0_stage68_subdone : BOOLEAN;
    signal ap_block_pp0_stage68_11001 : BOOLEAN;
    signal ap_block_state71_pp0_stage69_iter0 : BOOLEAN;
    signal ap_block_pp0_stage69_subdone : BOOLEAN;
    signal ap_block_pp0_stage69_11001 : BOOLEAN;
    signal ap_block_state72_pp0_stage70_iter0 : BOOLEAN;
    signal ap_block_pp0_stage70_subdone : BOOLEAN;
    signal ap_block_pp0_stage70_11001 : BOOLEAN;
    signal ap_block_state73_pp0_stage71_iter0 : BOOLEAN;
    signal ap_block_pp0_stage71_subdone : BOOLEAN;
    signal ap_block_pp0_stage71_11001 : BOOLEAN;
    signal ap_block_state74_pp0_stage72_iter0 : BOOLEAN;
    signal ap_block_pp0_stage72_subdone : BOOLEAN;
    signal ap_block_pp0_stage72_11001 : BOOLEAN;
    signal ap_block_pp0_stage73_subdone : BOOLEAN;
    signal ap_block_pp0_stage74_subdone : BOOLEAN;
    signal ap_block_pp0_stage75_subdone : BOOLEAN;
    signal ap_block_pp0_stage76_subdone : BOOLEAN;
    signal ap_block_state79_pp0_stage77_iter0 : BOOLEAN;
    signal ap_block_pp0_stage77_subdone : BOOLEAN;
    signal ap_block_pp0_stage77_11001 : BOOLEAN;
    signal ap_block_state80_pp0_stage78_iter0 : BOOLEAN;
    signal ap_block_pp0_stage78_subdone : BOOLEAN;
    signal ap_block_pp0_stage78_11001 : BOOLEAN;
    signal ap_block_state81_pp0_stage79_iter0 : BOOLEAN;
    signal ap_block_pp0_stage79_subdone : BOOLEAN;
    signal ap_block_pp0_stage79_11001 : BOOLEAN;
    signal ap_block_state82_pp0_stage80_iter0 : BOOLEAN;
    signal ap_block_pp0_stage80_subdone : BOOLEAN;
    signal ap_block_pp0_stage80_11001 : BOOLEAN;
    signal ap_block_pp0_stage81_subdone : BOOLEAN;
    signal ap_idle_pp0 : STD_LOGIC;
    signal ap_enable_pp0 : STD_LOGIC;
    signal ap_ce_reg : STD_LOGIC;

    component add_sub_mm_control_s_axi IS
    generic (
        C_S_AXI_ADDR_WIDTH : INTEGER;
        C_S_AXI_DATA_WIDTH : INTEGER );
    port (
        AWVALID : IN STD_LOGIC;
        AWREADY : OUT STD_LOGIC;
        AWADDR : IN STD_LOGIC_VECTOR (C_S_AXI_ADDR_WIDTH-1 downto 0);
        WVALID : IN STD_LOGIC;
        WREADY : OUT STD_LOGIC;
        WDATA : IN STD_LOGIC_VECTOR (C_S_AXI_DATA_WIDTH-1 downto 0);
        WSTRB : IN STD_LOGIC_VECTOR (C_S_AXI_DATA_WIDTH/8-1 downto 0);
        ARVALID : IN STD_LOGIC;
        ARREADY : OUT STD_LOGIC;
        ARADDR : IN STD_LOGIC_VECTOR (C_S_AXI_ADDR_WIDTH-1 downto 0);
        RVALID : OUT STD_LOGIC;
        RREADY : IN STD_LOGIC;
        RDATA : OUT STD_LOGIC_VECTOR (C_S_AXI_DATA_WIDTH-1 downto 0);
        RRESP : OUT STD_LOGIC_VECTOR (1 downto 0);
        BVALID : OUT STD_LOGIC;
        BREADY : IN STD_LOGIC;
        BRESP : OUT STD_LOGIC_VECTOR (1 downto 0);
        ACLK : IN STD_LOGIC;
        ARESET : IN STD_LOGIC;
        ACLK_EN : IN STD_LOGIC;
        arg1 : OUT STD_LOGIC_VECTOR (63 downto 0);
        arg2 : OUT STD_LOGIC_VECTOR (63 downto 0);
        mem : OUT STD_LOGIC_VECTOR (63 downto 0);
        src_addr1 : OUT STD_LOGIC_VECTOR (31 downto 0);
        src_addr2 : OUT STD_LOGIC_VECTOR (31 downto 0);
        dst_addr : OUT STD_LOGIC_VECTOR (31 downto 0);
        size : OUT STD_LOGIC_VECTOR (31 downto 0);
        op : OUT STD_LOGIC_VECTOR (0 downto 0);
        ap_start : OUT STD_LOGIC;
        interrupt : OUT STD_LOGIC;
        ap_ready : IN STD_LOGIC;
        ap_done : IN STD_LOGIC;
        ap_idle : IN STD_LOGIC );
    end component;


    component add_sub_mm_gmem_m_axi IS
    generic (
        CONSERVATIVE : INTEGER;
        USER_MAXREQS : INTEGER;
        NUM_READ_OUTSTANDING : INTEGER;
        NUM_WRITE_OUTSTANDING : INTEGER;
        MAX_READ_BURST_LENGTH : INTEGER;
        MAX_WRITE_BURST_LENGTH : INTEGER;
        USER_RFIFONUM_WIDTH : INTEGER;
        C_M_AXI_ID_WIDTH : INTEGER;
        C_M_AXI_ADDR_WIDTH : INTEGER;
        C_M_AXI_DATA_WIDTH : INTEGER;
        C_M_AXI_AWUSER_WIDTH : INTEGER;
        C_M_AXI_ARUSER_WIDTH : INTEGER;
        C_M_AXI_WUSER_WIDTH : INTEGER;
        C_M_AXI_RUSER_WIDTH : INTEGER;
        C_M_AXI_BUSER_WIDTH : INTEGER;
        C_USER_VALUE : INTEGER;
        C_PROT_VALUE : INTEGER;
        C_CACHE_VALUE : INTEGER;
        USER_DW : INTEGER;
        USER_AW : INTEGER );
    port (
        AWVALID : OUT STD_LOGIC;
        AWREADY : IN STD_LOGIC;
        AWADDR : OUT STD_LOGIC_VECTOR (C_M_AXI_ADDR_WIDTH-1 downto 0);
        AWID : OUT STD_LOGIC_VECTOR (C_M_AXI_ID_WIDTH-1 downto 0);
        AWLEN : OUT STD_LOGIC_VECTOR (7 downto 0);
        AWSIZE : OUT STD_LOGIC_VECTOR (2 downto 0);
        AWBURST : OUT STD_LOGIC_VECTOR (1 downto 0);
        AWLOCK : OUT STD_LOGIC_VECTOR (1 downto 0);
        AWCACHE : OUT STD_LOGIC_VECTOR (3 downto 0);
        AWPROT : OUT STD_LOGIC_VECTOR (2 downto 0);
        AWQOS : OUT STD_LOGIC_VECTOR (3 downto 0);
        AWREGION : OUT STD_LOGIC_VECTOR (3 downto 0);
        AWUSER : OUT STD_LOGIC_VECTOR (C_M_AXI_AWUSER_WIDTH-1 downto 0);
        WVALID : OUT STD_LOGIC;
        WREADY : IN STD_LOGIC;
        WDATA : OUT STD_LOGIC_VECTOR (C_M_AXI_DATA_WIDTH-1 downto 0);
        WSTRB : OUT STD_LOGIC_VECTOR (C_M_AXI_DATA_WIDTH/8-1 downto 0);
        WLAST : OUT STD_LOGIC;
        WID : OUT STD_LOGIC_VECTOR (C_M_AXI_ID_WIDTH-1 downto 0);
        WUSER : OUT STD_LOGIC_VECTOR (C_M_AXI_WUSER_WIDTH-1 downto 0);
        ARVALID : OUT STD_LOGIC;
        ARREADY : IN STD_LOGIC;
        ARADDR : OUT STD_LOGIC_VECTOR (C_M_AXI_ADDR_WIDTH-1 downto 0);
        ARID : OUT STD_LOGIC_VECTOR (C_M_AXI_ID_WIDTH-1 downto 0);
        ARLEN : OUT STD_LOGIC_VECTOR (7 downto 0);
        ARSIZE : OUT STD_LOGIC_VECTOR (2 downto 0);
        ARBURST : OUT STD_LOGIC_VECTOR (1 downto 0);
        ARLOCK : OUT STD_LOGIC_VECTOR (1 downto 0);
        ARCACHE : OUT STD_LOGIC_VECTOR (3 downto 0);
        ARPROT : OUT STD_LOGIC_VECTOR (2 downto 0);
        ARQOS : OUT STD_LOGIC_VECTOR (3 downto 0);
        ARREGION : OUT STD_LOGIC_VECTOR (3 downto 0);
        ARUSER : OUT STD_LOGIC_VECTOR (C_M_AXI_ARUSER_WIDTH-1 downto 0);
        RVALID : IN STD_LOGIC;
        RREADY : OUT STD_LOGIC;
        RDATA : IN STD_LOGIC_VECTOR (C_M_AXI_DATA_WIDTH-1 downto 0);
        RLAST : IN STD_LOGIC;
        RID : IN STD_LOGIC_VECTOR (C_M_AXI_ID_WIDTH-1 downto 0);
        RUSER : IN STD_LOGIC_VECTOR (C_M_AXI_RUSER_WIDTH-1 downto 0);
        RRESP : IN STD_LOGIC_VECTOR (1 downto 0);
        BVALID : IN STD_LOGIC;
        BREADY : OUT STD_LOGIC;
        BRESP : IN STD_LOGIC_VECTOR (1 downto 0);
        BID : IN STD_LOGIC_VECTOR (C_M_AXI_ID_WIDTH-1 downto 0);
        BUSER : IN STD_LOGIC_VECTOR (C_M_AXI_BUSER_WIDTH-1 downto 0);
        ACLK : IN STD_LOGIC;
        ARESET : IN STD_LOGIC;
        ACLK_EN : IN STD_LOGIC;
        I_ARVALID : IN STD_LOGIC;
        I_ARREADY : OUT STD_LOGIC;
        I_ARADDR : IN STD_LOGIC_VECTOR (63 downto 0);
        I_ARLEN : IN STD_LOGIC_VECTOR (31 downto 0);
        I_RVALID : OUT STD_LOGIC;
        I_RREADY : IN STD_LOGIC;
        I_RDATA : OUT STD_LOGIC_VECTOR (127 downto 0);
        I_RFIFONUM : OUT STD_LOGIC_VECTOR (8 downto 0);
        I_AWVALID : IN STD_LOGIC;
        I_AWREADY : OUT STD_LOGIC;
        I_AWADDR : IN STD_LOGIC_VECTOR (63 downto 0);
        I_AWLEN : IN STD_LOGIC_VECTOR (31 downto 0);
        I_WVALID : IN STD_LOGIC;
        I_WREADY : OUT STD_LOGIC;
        I_WDATA : IN STD_LOGIC_VECTOR (127 downto 0);
        I_WSTRB : IN STD_LOGIC_VECTOR (15 downto 0);
        I_BVALID : OUT STD_LOGIC;
        I_BREADY : IN STD_LOGIC );
    end component;



begin
    control_s_axi_U : component add_sub_mm_control_s_axi
    generic map (
        C_S_AXI_ADDR_WIDTH => C_S_AXI_CONTROL_ADDR_WIDTH,
        C_S_AXI_DATA_WIDTH => C_S_AXI_CONTROL_DATA_WIDTH)
    port map (
        AWVALID => s_axi_control_AWVALID,
        AWREADY => s_axi_control_AWREADY,
        AWADDR => s_axi_control_AWADDR,
        WVALID => s_axi_control_WVALID,
        WREADY => s_axi_control_WREADY,
        WDATA => s_axi_control_WDATA,
        WSTRB => s_axi_control_WSTRB,
        ARVALID => s_axi_control_ARVALID,
        ARREADY => s_axi_control_ARREADY,
        ARADDR => s_axi_control_ARADDR,
        RVALID => s_axi_control_RVALID,
        RREADY => s_axi_control_RREADY,
        RDATA => s_axi_control_RDATA,
        RRESP => s_axi_control_RRESP,
        BVALID => s_axi_control_BVALID,
        BREADY => s_axi_control_BREADY,
        BRESP => s_axi_control_BRESP,
        ACLK => ap_clk,
        ARESET => ap_rst_n_inv,
        ACLK_EN => ap_const_logic_1,
        arg1 => arg1,
        arg2 => arg2,
        mem => mem,
        src_addr1 => src_addr1,
        src_addr2 => src_addr2,
        dst_addr => dst_addr,
        size => size,
        op => op,
        ap_start => ap_start,
        interrupt => interrupt,
        ap_ready => ap_ready,
        ap_done => ap_done,
        ap_idle => ap_idle);

    gmem_m_axi_U : component add_sub_mm_gmem_m_axi
    generic map (
        CONSERVATIVE => 1,
        USER_MAXREQS => 5,
        NUM_READ_OUTSTANDING => 16,
        NUM_WRITE_OUTSTANDING => 16,
        MAX_READ_BURST_LENGTH => 16,
        MAX_WRITE_BURST_LENGTH => 16,
        USER_RFIFONUM_WIDTH => 9,
        C_M_AXI_ID_WIDTH => C_M_AXI_GMEM_ID_WIDTH,
        C_M_AXI_ADDR_WIDTH => C_M_AXI_GMEM_ADDR_WIDTH,
        C_M_AXI_DATA_WIDTH => C_M_AXI_GMEM_DATA_WIDTH,
        C_M_AXI_AWUSER_WIDTH => C_M_AXI_GMEM_AWUSER_WIDTH,
        C_M_AXI_ARUSER_WIDTH => C_M_AXI_GMEM_ARUSER_WIDTH,
        C_M_AXI_WUSER_WIDTH => C_M_AXI_GMEM_WUSER_WIDTH,
        C_M_AXI_RUSER_WIDTH => C_M_AXI_GMEM_RUSER_WIDTH,
        C_M_AXI_BUSER_WIDTH => C_M_AXI_GMEM_BUSER_WIDTH,
        C_USER_VALUE => C_M_AXI_GMEM_USER_VALUE,
        C_PROT_VALUE => C_M_AXI_GMEM_PROT_VALUE,
        C_CACHE_VALUE => C_M_AXI_GMEM_CACHE_VALUE,
        USER_DW => 128,
        USER_AW => 64)
    port map (
        AWVALID => m_axi_gmem_AWVALID,
        AWREADY => m_axi_gmem_AWREADY,
        AWADDR => m_axi_gmem_AWADDR,
        AWID => m_axi_gmem_AWID,
        AWLEN => m_axi_gmem_AWLEN,
        AWSIZE => m_axi_gmem_AWSIZE,
        AWBURST => m_axi_gmem_AWBURST,
        AWLOCK => m_axi_gmem_AWLOCK,
        AWCACHE => m_axi_gmem_AWCACHE,
        AWPROT => m_axi_gmem_AWPROT,
        AWQOS => m_axi_gmem_AWQOS,
        AWREGION => m_axi_gmem_AWREGION,
        AWUSER => m_axi_gmem_AWUSER,
        WVALID => m_axi_gmem_WVALID,
        WREADY => m_axi_gmem_WREADY,
        WDATA => m_axi_gmem_WDATA,
        WSTRB => m_axi_gmem_WSTRB,
        WLAST => m_axi_gmem_WLAST,
        WID => m_axi_gmem_WID,
        WUSER => m_axi_gmem_WUSER,
        ARVALID => m_axi_gmem_ARVALID,
        ARREADY => m_axi_gmem_ARREADY,
        ARADDR => m_axi_gmem_ARADDR,
        ARID => m_axi_gmem_ARID,
        ARLEN => m_axi_gmem_ARLEN,
        ARSIZE => m_axi_gmem_ARSIZE,
        ARBURST => m_axi_gmem_ARBURST,
        ARLOCK => m_axi_gmem_ARLOCK,
        ARCACHE => m_axi_gmem_ARCACHE,
        ARPROT => m_axi_gmem_ARPROT,
        ARQOS => m_axi_gmem_ARQOS,
        ARREGION => m_axi_gmem_ARREGION,
        ARUSER => m_axi_gmem_ARUSER,
        RVALID => m_axi_gmem_RVALID,
        RREADY => m_axi_gmem_RREADY,
        RDATA => m_axi_gmem_RDATA,
        RLAST => m_axi_gmem_RLAST,
        RID => m_axi_gmem_RID,
        RUSER => m_axi_gmem_RUSER,
        RRESP => m_axi_gmem_RRESP,
        BVALID => m_axi_gmem_BVALID,
        BREADY => m_axi_gmem_BREADY,
        BRESP => m_axi_gmem_BRESP,
        BID => m_axi_gmem_BID,
        BUSER => m_axi_gmem_BUSER,
        ACLK => ap_clk,
        ARESET => ap_rst_n_inv,
        ACLK_EN => ap_const_logic_1,
        I_ARVALID => gmem_ARVALID,
        I_ARREADY => gmem_ARREADY,
        I_ARADDR => gmem_ARADDR,
        I_ARLEN => ap_const_lv32_1,
        I_RVALID => gmem_RVALID,
        I_RREADY => gmem_RREADY,
        I_RDATA => gmem_RDATA,
        I_RFIFONUM => gmem_RFIFONUM,
        I_AWVALID => gmem_AWVALID,
        I_AWREADY => gmem_AWREADY,
        I_AWADDR => gmem_AWADDR,
        I_AWLEN => ap_const_lv32_1,
        I_WVALID => gmem_WVALID,
        I_WREADY => gmem_WREADY,
        I_WDATA => gmem_WDATA,
        I_WSTRB => gmem_WSTRB,
        I_BVALID => gmem_BVALID,
        I_BREADY => gmem_BREADY);





    ap_CS_fsm_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_CS_fsm <= ap_ST_fsm_state1;
            else
                ap_CS_fsm <= ap_NS_fsm;
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter0_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter0 <= ap_const_logic_0;
            else
                if (((ap_const_logic_1 = ap_CS_fsm_pp0_stage0) and (ap_const_logic_1 = ap_condition_pp0_exit_iter0_state2) and (ap_const_boolean_0 = ap_block_pp0_stage0_subdone))) then 
                    ap_enable_reg_pp0_iter0 <= ap_const_logic_0;
                elsif (((ap_start = ap_const_logic_1) and (ap_const_logic_1 = ap_CS_fsm_state1))) then 
                    ap_enable_reg_pp0_iter0 <= ap_const_logic_1;
                end if; 
            end if;
        end if;
    end process;


    ap_enable_reg_pp0_iter1_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst_n_inv = '1') then
                ap_enable_reg_pp0_iter1 <= ap_const_logic_0;
            else
                if ((((ap_const_logic_1 = ap_CS_fsm_pp0_stage14) and (ap_const_boolean_0 = ap_block_pp0_stage14_subdone) and (ap_enable_reg_pp0_iter0 = ap_const_logic_0)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage82) and (ap_const_boolean_0 = ap_block_pp0_stage82_subdone)))) then 
                    ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
                elsif (((ap_start = ap_const_logic_1) and (ap_const_logic_1 = ap_CS_fsm_state1))) then 
                    ap_enable_reg_pp0_iter1 <= ap_const_logic_0;
                end if; 
            end if;
        end if;
    end process;


    ap_phi_reg_pp0_iter1_storemerge_reg_250_assign_proc : process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((icmp_ln1073_reg_676_pp0_iter1_reg = ap_const_lv1_1) and (ap_enable_reg_pp0_iter1 = ap_const_logic_1) and (op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage8) and (ap_const_boolean_0 = ap_block_pp0_stage8_11001))) then 
                ap_phi_reg_pp0_iter1_storemerge_reg_250 <= p_Result_s_fu_624_p5;
            elsif (((ap_const_logic_1 = ap_CS_fsm_pp0_stage82) and (ap_const_boolean_0 = ap_block_pp0_stage82_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1))) then 
                ap_phi_reg_pp0_iter1_storemerge_reg_250 <= ap_phi_reg_pp0_iter0_storemerge_reg_250;
            end if; 
        end if;
    end process;

    rhs_V_fu_122_assign_proc : process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_start = ap_const_logic_1) and (ap_const_logic_1 = ap_CS_fsm_state1))) then 
                rhs_V_fu_122 <= ap_const_lv32_0;
            elsif (((ap_const_logic_1 = ap_CS_fsm_pp0_stage82) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage82_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1))) then 
                rhs_V_fu_122 <= i_V_fu_608_p2;
            end if; 
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage10) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage10_11001))) then
                add_ln414_1_reg_739 <= add_ln414_1_fu_511_p2;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage59) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage59_11001))) then
                add_ln414_2_reg_765 <= add_ln414_2_fu_573_p2;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage75) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage75_11001))) then
                add_ln414_3_reg_772 <= add_ln414_3_fu_590_p2;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage58) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage58_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1))) then
                ap_phi_reg_pp0_iter0_storemerge_reg_250 <= p_Result_4_fu_564_p5;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_const_logic_1 = ap_CS_fsm_pp0_stage2) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage2_11001))) then
                gmem_addr_1_reg_713 <= sext_ln357_1_fu_489_p1;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_const_logic_1 = ap_CS_fsm_pp0_stage1) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage1_11001))) then
                gmem_addr_2_reg_701 <= sext_ln414_fu_479_p1;
                gmem_addr_reg_695 <= sext_ln357_fu_469_p1;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_const_logic_1 = ap_CS_fsm_pp0_stage0) and (ap_const_boolean_0 = ap_block_pp0_stage0_11001))) then
                i_V_2_reg_671 <= rhs_V_fu_122;
                icmp_ln1073_reg_676 <= icmp_ln1073_fu_364_p2;
                icmp_ln1073_reg_676_pp0_iter1_reg <= icmp_ln1073_reg_676;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if ((ap_const_logic_1 = ap_CS_fsm_state1)) then
                    lhs_5_reg_661(31 downto 0) <= lhs_5_fu_348_p1(31 downto 0);
                    lhs_6_reg_666(31 downto 0) <= lhs_6_fu_352_p1(31 downto 0);
                    lhs_reg_656(31 downto 0) <= lhs_fu_344_p1(31 downto 0);
                mem_read_reg_649 <= mem;
                op_read_reg_640 <= op;
                size_read_reg_644 <= size;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if ((((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage24) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage24_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage57) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage57_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)))) then
                reg_320 <= gmem_RDATA(63 downto 32);
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if ((((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage25) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage25_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage58) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage58_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)))) then
                reg_324 <= gmem_RDATA(63 downto 32);
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if ((((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage40) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage40_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage73) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage73_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)))) then
                reg_328 <= gmem_RDATA(95 downto 64);
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if ((((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage41) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage41_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage74) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage74_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)))) then
                reg_332 <= gmem_RDATA(95 downto 64);
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if ((((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage56) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage56_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((icmp_ln1073_reg_676_pp0_iter1_reg = ap_const_lv1_1) and (ap_enable_reg_pp0_iter1 = ap_const_logic_1) and (op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage6) and (ap_const_boolean_0 = ap_block_pp0_stage6_11001)))) then
                reg_336 <= gmem_RDATA(127 downto 96);
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if ((((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage57) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage57_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((icmp_ln1073_reg_676_pp0_iter1_reg = ap_const_lv1_1) and (ap_enable_reg_pp0_iter1 = ap_const_logic_1) and (op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage7) and (ap_const_boolean_0 = ap_block_pp0_stage7_11001)))) then
                reg_340 <= gmem_RDATA(127 downto 96);
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage26) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage26_11001))) then
                sub_ln414_1_reg_747 <= sub_ln414_1_fu_519_p2;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage42) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage42_11001))) then
                sub_ln414_2_reg_754 <= sub_ln414_2_fu_536_p2;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage10) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage10_11001))) then
                sub_ln414_reg_731 <= sub_ln414_fu_507_p2;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((icmp_ln1073_fu_364_p2 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0) and (ap_const_boolean_0 = ap_block_pp0_stage0_11001))) then
                trunc_ln1_reg_690 <= add_ln414_fu_434_p2(63 downto 4);
                trunc_ln357_1_reg_685 <= add_ln357_1_fu_412_p2(63 downto 4);
                trunc_ln_reg_680 <= add_ln357_fu_395_p2(63 downto 4);
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_const_logic_1 = ap_CS_fsm_pp0_stage9) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage9_11001))) then
                trunc_ln357_2_reg_725 <= trunc_ln357_2_fu_503_p1;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_const_logic_1 = ap_CS_fsm_pp0_stage8) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage8_11001))) then
                trunc_ln357_reg_719 <= trunc_ln357_fu_499_p1;
            end if;
        end if;
    end process;
    lhs_reg_656(33 downto 32) <= "00";
    lhs_5_reg_661(33 downto 32) <= "00";
    lhs_6_reg_666(33 downto 32) <= "00";

    ap_NS_fsm_assign_proc : process (ap_start, ap_CS_fsm, ap_CS_fsm_state1, ap_enable_reg_pp0_iter0, ap_enable_reg_pp0_iter1, ap_CS_fsm_pp0_stage14, icmp_ln1073_fu_364_p2, ap_block_pp0_stage0_subdone, ap_block_pp0_stage82_subdone, ap_block_pp0_stage14_subdone, ap_block_pp0_stage1_subdone, ap_block_pp0_stage2_subdone, ap_block_pp0_stage3_subdone, ap_block_pp0_stage4_subdone, ap_block_pp0_stage5_subdone, ap_block_pp0_stage6_subdone, ap_block_pp0_stage7_subdone, ap_block_pp0_stage8_subdone, ap_block_pp0_stage9_subdone, ap_block_pp0_stage10_subdone, ap_block_pp0_stage11_subdone, ap_block_pp0_stage12_subdone, ap_block_pp0_stage13_subdone, ap_block_pp0_stage15_subdone, ap_block_pp0_stage16_subdone, ap_block_pp0_stage17_subdone, ap_block_pp0_stage18_subdone, ap_block_pp0_stage19_subdone, ap_block_pp0_stage20_subdone, ap_block_pp0_stage21_subdone, ap_block_pp0_stage22_subdone, ap_block_pp0_stage23_subdone, ap_block_pp0_stage24_subdone, ap_block_pp0_stage25_subdone, ap_block_pp0_stage26_subdone, ap_block_pp0_stage27_subdone, ap_block_pp0_stage28_subdone, ap_block_pp0_stage29_subdone, ap_block_pp0_stage30_subdone, ap_block_pp0_stage31_subdone, ap_block_pp0_stage32_subdone, ap_block_pp0_stage33_subdone, ap_block_pp0_stage34_subdone, ap_block_pp0_stage35_subdone, ap_block_pp0_stage36_subdone, ap_block_pp0_stage37_subdone, ap_block_pp0_stage38_subdone, ap_block_pp0_stage39_subdone, ap_block_pp0_stage40_subdone, ap_block_pp0_stage41_subdone, ap_block_pp0_stage42_subdone, ap_block_pp0_stage43_subdone, ap_block_pp0_stage44_subdone, ap_block_pp0_stage45_subdone, ap_block_pp0_stage46_subdone, ap_block_pp0_stage47_subdone, ap_block_pp0_stage48_subdone, ap_block_pp0_stage49_subdone, ap_block_pp0_stage50_subdone, ap_block_pp0_stage51_subdone, ap_block_pp0_stage52_subdone, ap_block_pp0_stage53_subdone, ap_block_pp0_stage54_subdone, ap_block_pp0_stage55_subdone, ap_block_pp0_stage56_subdone, ap_block_pp0_stage57_subdone, ap_block_pp0_stage58_subdone, ap_block_pp0_stage59_subdone, ap_block_pp0_stage60_subdone, ap_block_pp0_stage61_subdone, ap_block_pp0_stage62_subdone, ap_block_pp0_stage63_subdone, ap_block_pp0_stage64_subdone, ap_block_pp0_stage65_subdone, ap_block_pp0_stage66_subdone, ap_block_pp0_stage67_subdone, ap_block_pp0_stage68_subdone, ap_block_pp0_stage69_subdone, ap_block_pp0_stage70_subdone, ap_block_pp0_stage71_subdone, ap_block_pp0_stage72_subdone, ap_block_pp0_stage73_subdone, ap_block_pp0_stage74_subdone, ap_block_pp0_stage75_subdone, ap_block_pp0_stage76_subdone, ap_block_pp0_stage77_subdone, ap_block_pp0_stage78_subdone, ap_block_pp0_stage79_subdone, ap_block_pp0_stage80_subdone, ap_block_pp0_stage81_subdone)
    begin
        case ap_CS_fsm is
            when ap_ST_fsm_state1 => 
                if (((ap_start = ap_const_logic_1) and (ap_const_logic_1 = ap_CS_fsm_state1))) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage0;
                else
                    ap_NS_fsm <= ap_ST_fsm_state1;
                end if;
            when ap_ST_fsm_pp0_stage0 => 
                if ((not(((icmp_ln1073_fu_364_p2 = ap_const_lv1_0) and (ap_enable_reg_pp0_iter1 = ap_const_logic_0) and (ap_const_boolean_0 = ap_block_pp0_stage0_subdone) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1))) and (ap_const_boolean_0 = ap_block_pp0_stage0_subdone))) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage1;
                elsif (((icmp_ln1073_fu_364_p2 = ap_const_lv1_0) and (ap_enable_reg_pp0_iter1 = ap_const_logic_0) and (ap_const_boolean_0 = ap_block_pp0_stage0_subdone) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1))) then
                    ap_NS_fsm <= ap_ST_fsm_state100;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage0;
                end if;
            when ap_ST_fsm_pp0_stage1 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage1_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage2;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage1;
                end if;
            when ap_ST_fsm_pp0_stage2 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage2_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage3;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage2;
                end if;
            when ap_ST_fsm_pp0_stage3 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage3_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage4;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage3;
                end if;
            when ap_ST_fsm_pp0_stage4 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage4_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage5;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage4;
                end if;
            when ap_ST_fsm_pp0_stage5 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage5_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage6;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage5;
                end if;
            when ap_ST_fsm_pp0_stage6 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage6_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage7;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage6;
                end if;
            when ap_ST_fsm_pp0_stage7 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage7_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage8;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage7;
                end if;
            when ap_ST_fsm_pp0_stage8 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage8_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage9;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage8;
                end if;
            when ap_ST_fsm_pp0_stage9 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage9_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage10;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage9;
                end if;
            when ap_ST_fsm_pp0_stage10 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage10_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage11;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage10;
                end if;
            when ap_ST_fsm_pp0_stage11 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage11_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage12;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage11;
                end if;
            when ap_ST_fsm_pp0_stage12 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage12_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage13;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage12;
                end if;
            when ap_ST_fsm_pp0_stage13 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage13_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage14;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage13;
                end if;
            when ap_ST_fsm_pp0_stage14 => 
                if ((not(((ap_enable_reg_pp0_iter1 = ap_const_logic_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage14) and (ap_const_boolean_0 = ap_block_pp0_stage14_subdone) and (ap_enable_reg_pp0_iter0 = ap_const_logic_0))) and (ap_const_boolean_0 = ap_block_pp0_stage14_subdone))) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage15;
                elsif (((ap_enable_reg_pp0_iter1 = ap_const_logic_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage14) and (ap_const_boolean_0 = ap_block_pp0_stage14_subdone) and (ap_enable_reg_pp0_iter0 = ap_const_logic_0))) then
                    ap_NS_fsm <= ap_ST_fsm_state100;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage14;
                end if;
            when ap_ST_fsm_pp0_stage15 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage15_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage16;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage15;
                end if;
            when ap_ST_fsm_pp0_stage16 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage16_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage17;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage16;
                end if;
            when ap_ST_fsm_pp0_stage17 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage17_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage18;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage17;
                end if;
            when ap_ST_fsm_pp0_stage18 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage18_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage19;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage18;
                end if;
            when ap_ST_fsm_pp0_stage19 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage19_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage20;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage19;
                end if;
            when ap_ST_fsm_pp0_stage20 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage20_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage21;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage20;
                end if;
            when ap_ST_fsm_pp0_stage21 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage21_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage22;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage21;
                end if;
            when ap_ST_fsm_pp0_stage22 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage22_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage23;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage22;
                end if;
            when ap_ST_fsm_pp0_stage23 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage23_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage24;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage23;
                end if;
            when ap_ST_fsm_pp0_stage24 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage24_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage25;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage24;
                end if;
            when ap_ST_fsm_pp0_stage25 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage25_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage26;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage25;
                end if;
            when ap_ST_fsm_pp0_stage26 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage26_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage27;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage26;
                end if;
            when ap_ST_fsm_pp0_stage27 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage27_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage28;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage27;
                end if;
            when ap_ST_fsm_pp0_stage28 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage28_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage29;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage28;
                end if;
            when ap_ST_fsm_pp0_stage29 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage29_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage30;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage29;
                end if;
            when ap_ST_fsm_pp0_stage30 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage30_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage31;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage30;
                end if;
            when ap_ST_fsm_pp0_stage31 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage31_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage32;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage31;
                end if;
            when ap_ST_fsm_pp0_stage32 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage32_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage33;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage32;
                end if;
            when ap_ST_fsm_pp0_stage33 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage33_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage34;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage33;
                end if;
            when ap_ST_fsm_pp0_stage34 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage34_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage35;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage34;
                end if;
            when ap_ST_fsm_pp0_stage35 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage35_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage36;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage35;
                end if;
            when ap_ST_fsm_pp0_stage36 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage36_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage37;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage36;
                end if;
            when ap_ST_fsm_pp0_stage37 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage37_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage38;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage37;
                end if;
            when ap_ST_fsm_pp0_stage38 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage38_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage39;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage38;
                end if;
            when ap_ST_fsm_pp0_stage39 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage39_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage40;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage39;
                end if;
            when ap_ST_fsm_pp0_stage40 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage40_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage41;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage40;
                end if;
            when ap_ST_fsm_pp0_stage41 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage41_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage42;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage41;
                end if;
            when ap_ST_fsm_pp0_stage42 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage42_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage43;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage42;
                end if;
            when ap_ST_fsm_pp0_stage43 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage43_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage44;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage43;
                end if;
            when ap_ST_fsm_pp0_stage44 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage44_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage45;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage44;
                end if;
            when ap_ST_fsm_pp0_stage45 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage45_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage46;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage45;
                end if;
            when ap_ST_fsm_pp0_stage46 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage46_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage47;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage46;
                end if;
            when ap_ST_fsm_pp0_stage47 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage47_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage48;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage47;
                end if;
            when ap_ST_fsm_pp0_stage48 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage48_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage49;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage48;
                end if;
            when ap_ST_fsm_pp0_stage49 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage49_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage50;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage49;
                end if;
            when ap_ST_fsm_pp0_stage50 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage50_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage51;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage50;
                end if;
            when ap_ST_fsm_pp0_stage51 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage51_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage52;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage51;
                end if;
            when ap_ST_fsm_pp0_stage52 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage52_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage53;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage52;
                end if;
            when ap_ST_fsm_pp0_stage53 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage53_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage54;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage53;
                end if;
            when ap_ST_fsm_pp0_stage54 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage54_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage55;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage54;
                end if;
            when ap_ST_fsm_pp0_stage55 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage55_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage56;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage55;
                end if;
            when ap_ST_fsm_pp0_stage56 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage56_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage57;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage56;
                end if;
            when ap_ST_fsm_pp0_stage57 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage57_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage58;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage57;
                end if;
            when ap_ST_fsm_pp0_stage58 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage58_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage59;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage58;
                end if;
            when ap_ST_fsm_pp0_stage59 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage59_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage60;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage59;
                end if;
            when ap_ST_fsm_pp0_stage60 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage60_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage61;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage60;
                end if;
            when ap_ST_fsm_pp0_stage61 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage61_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage62;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage61;
                end if;
            when ap_ST_fsm_pp0_stage62 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage62_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage63;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage62;
                end if;
            when ap_ST_fsm_pp0_stage63 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage63_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage64;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage63;
                end if;
            when ap_ST_fsm_pp0_stage64 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage64_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage65;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage64;
                end if;
            when ap_ST_fsm_pp0_stage65 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage65_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage66;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage65;
                end if;
            when ap_ST_fsm_pp0_stage66 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage66_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage67;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage66;
                end if;
            when ap_ST_fsm_pp0_stage67 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage67_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage68;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage67;
                end if;
            when ap_ST_fsm_pp0_stage68 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage68_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage69;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage68;
                end if;
            when ap_ST_fsm_pp0_stage69 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage69_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage70;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage69;
                end if;
            when ap_ST_fsm_pp0_stage70 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage70_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage71;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage70;
                end if;
            when ap_ST_fsm_pp0_stage71 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage71_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage72;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage71;
                end if;
            when ap_ST_fsm_pp0_stage72 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage72_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage73;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage72;
                end if;
            when ap_ST_fsm_pp0_stage73 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage73_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage74;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage73;
                end if;
            when ap_ST_fsm_pp0_stage74 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage74_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage75;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage74;
                end if;
            when ap_ST_fsm_pp0_stage75 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage75_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage76;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage75;
                end if;
            when ap_ST_fsm_pp0_stage76 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage76_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage77;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage76;
                end if;
            when ap_ST_fsm_pp0_stage77 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage77_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage78;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage77;
                end if;
            when ap_ST_fsm_pp0_stage78 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage78_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage79;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage78;
                end if;
            when ap_ST_fsm_pp0_stage79 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage79_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage80;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage79;
                end if;
            when ap_ST_fsm_pp0_stage80 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage80_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage81;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage80;
                end if;
            when ap_ST_fsm_pp0_stage81 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage81_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage82;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage81;
                end if;
            when ap_ST_fsm_pp0_stage82 => 
                if ((ap_const_boolean_0 = ap_block_pp0_stage82_subdone)) then
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage0;
                else
                    ap_NS_fsm <= ap_ST_fsm_pp0_stage82;
                end if;
            when ap_ST_fsm_state100 => 
                ap_NS_fsm <= ap_ST_fsm_state1;
            when others =>  
                ap_NS_fsm <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
        end case;
    end process;
    add_ln357_1_fu_412_p2 <= std_logic_vector(signed(sext_ln357_3_fu_408_p1) + signed(mem_read_reg_649));
    add_ln357_fu_395_p2 <= std_logic_vector(signed(sext_ln357_2_fu_391_p1) + signed(mem_read_reg_649));
    add_ln414_1_fu_511_p2 <= std_logic_vector(unsigned(trunc_ln357_2_reg_725) + unsigned(trunc_ln357_reg_719));
    add_ln414_2_fu_573_p2 <= std_logic_vector(unsigned(reg_324) + unsigned(reg_320));
    add_ln414_3_fu_590_p2 <= std_logic_vector(unsigned(reg_332) + unsigned(reg_328));
    add_ln414_4_fu_618_p2 <= std_logic_vector(unsigned(reg_340) + unsigned(reg_336));
    add_ln414_fu_434_p2 <= std_logic_vector(signed(sext_ln414_1_fu_430_p1) + signed(mem_read_reg_649));
    ap_CS_fsm_pp0_stage0 <= ap_CS_fsm(1);
    ap_CS_fsm_pp0_stage1 <= ap_CS_fsm(2);
    ap_CS_fsm_pp0_stage10 <= ap_CS_fsm(11);
    ap_CS_fsm_pp0_stage11 <= ap_CS_fsm(12);
    ap_CS_fsm_pp0_stage14 <= ap_CS_fsm(15);
    ap_CS_fsm_pp0_stage16 <= ap_CS_fsm(17);
    ap_CS_fsm_pp0_stage17 <= ap_CS_fsm(18);
    ap_CS_fsm_pp0_stage18 <= ap_CS_fsm(19);
    ap_CS_fsm_pp0_stage2 <= ap_CS_fsm(3);
    ap_CS_fsm_pp0_stage24 <= ap_CS_fsm(25);
    ap_CS_fsm_pp0_stage25 <= ap_CS_fsm(26);
    ap_CS_fsm_pp0_stage26 <= ap_CS_fsm(27);
    ap_CS_fsm_pp0_stage27 <= ap_CS_fsm(28);
    ap_CS_fsm_pp0_stage3 <= ap_CS_fsm(4);
    ap_CS_fsm_pp0_stage32 <= ap_CS_fsm(33);
    ap_CS_fsm_pp0_stage33 <= ap_CS_fsm(34);
    ap_CS_fsm_pp0_stage34 <= ap_CS_fsm(35);
    ap_CS_fsm_pp0_stage40 <= ap_CS_fsm(41);
    ap_CS_fsm_pp0_stage41 <= ap_CS_fsm(42);
    ap_CS_fsm_pp0_stage42 <= ap_CS_fsm(43);
    ap_CS_fsm_pp0_stage43 <= ap_CS_fsm(44);
    ap_CS_fsm_pp0_stage44 <= ap_CS_fsm(45);
    ap_CS_fsm_pp0_stage48 <= ap_CS_fsm(49);
    ap_CS_fsm_pp0_stage49 <= ap_CS_fsm(50);
    ap_CS_fsm_pp0_stage50 <= ap_CS_fsm(51);
    ap_CS_fsm_pp0_stage51 <= ap_CS_fsm(52);
    ap_CS_fsm_pp0_stage56 <= ap_CS_fsm(57);
    ap_CS_fsm_pp0_stage57 <= ap_CS_fsm(58);
    ap_CS_fsm_pp0_stage58 <= ap_CS_fsm(59);
    ap_CS_fsm_pp0_stage59 <= ap_CS_fsm(60);
    ap_CS_fsm_pp0_stage6 <= ap_CS_fsm(7);
    ap_CS_fsm_pp0_stage60 <= ap_CS_fsm(61);
    ap_CS_fsm_pp0_stage65 <= ap_CS_fsm(66);
    ap_CS_fsm_pp0_stage66 <= ap_CS_fsm(67);
    ap_CS_fsm_pp0_stage67 <= ap_CS_fsm(68);
    ap_CS_fsm_pp0_stage7 <= ap_CS_fsm(8);
    ap_CS_fsm_pp0_stage73 <= ap_CS_fsm(74);
    ap_CS_fsm_pp0_stage74 <= ap_CS_fsm(75);
    ap_CS_fsm_pp0_stage75 <= ap_CS_fsm(76);
    ap_CS_fsm_pp0_stage76 <= ap_CS_fsm(77);
    ap_CS_fsm_pp0_stage8 <= ap_CS_fsm(9);
    ap_CS_fsm_pp0_stage81 <= ap_CS_fsm(82);
    ap_CS_fsm_pp0_stage82 <= ap_CS_fsm(83);
    ap_CS_fsm_pp0_stage9 <= ap_CS_fsm(10);
    ap_CS_fsm_state1 <= ap_CS_fsm(0);
    ap_CS_fsm_state100 <= ap_CS_fsm(84);
    ap_ST_fsm_state100_blk <= ap_const_logic_0;

    ap_ST_fsm_state1_blk_assign_proc : process(ap_start)
    begin
        if ((ap_start = ap_const_logic_0)) then 
            ap_ST_fsm_state1_blk <= ap_const_logic_1;
        else 
            ap_ST_fsm_state1_blk <= ap_const_logic_0;
        end if; 
    end process;

        ap_block_pp0_stage0 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage0_11001_assign_proc : process(ap_enable_reg_pp0_iter1, ap_block_state85_io)
    begin
                ap_block_pp0_stage0_11001 <= ((ap_enable_reg_pp0_iter1 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state85_io));
    end process;


    ap_block_pp0_stage0_subdone_assign_proc : process(ap_enable_reg_pp0_iter1, ap_block_state85_io)
    begin
                ap_block_pp0_stage0_subdone <= ((ap_enable_reg_pp0_iter1 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state85_io));
    end process;

        ap_block_pp0_stage1 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage10 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage10_11001_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state12_io)
    begin
                ap_block_pp0_stage10_11001 <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state12_io));
    end process;


    ap_block_pp0_stage10_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state12_io)
    begin
                ap_block_pp0_stage10_subdone <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state12_io));
    end process;

        ap_block_pp0_stage11 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage11_01001 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage11_11001_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state13_io)
    begin
                ap_block_pp0_stage11_11001 <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state13_io));
    end process;


    ap_block_pp0_stage11_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state13_io)
    begin
                ap_block_pp0_stage11_subdone <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state13_io));
    end process;

        ap_block_pp0_stage12_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage12_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage13_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage13_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage14 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage14_11001_assign_proc : process(ap_enable_reg_pp0_iter1, gmem_BVALID)
    begin
                ap_block_pp0_stage14_11001 <= ((gmem_BVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter1 = ap_const_logic_1));
    end process;


    ap_block_pp0_stage14_subdone_assign_proc : process(ap_enable_reg_pp0_iter1, gmem_BVALID)
    begin
                ap_block_pp0_stage14_subdone <= ((gmem_BVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter1 = ap_const_logic_1));
    end process;

        ap_block_pp0_stage15_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage15_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage16 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage16_11001_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_BVALID, ap_predicate_op199_writeresp_state18)
    begin
                ap_block_pp0_stage16_11001 <= ((gmem_BVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op199_writeresp_state18 = ap_const_boolean_1));
    end process;


    ap_block_pp0_stage16_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_BVALID, ap_predicate_op199_writeresp_state18)
    begin
                ap_block_pp0_stage16_subdone <= ((gmem_BVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op199_writeresp_state18 = ap_const_boolean_1));
    end process;

        ap_block_pp0_stage17 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage17_11001_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state19_io)
    begin
                ap_block_pp0_stage17_11001 <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state19_io));
    end process;


    ap_block_pp0_stage17_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state19_io)
    begin
                ap_block_pp0_stage17_subdone <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state19_io));
    end process;

        ap_block_pp0_stage18 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage18_11001_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state20_io)
    begin
                ap_block_pp0_stage18_11001 <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state20_io));
    end process;


    ap_block_pp0_stage18_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state20_io)
    begin
                ap_block_pp0_stage18_subdone <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state20_io));
    end process;

        ap_block_pp0_stage19_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage19_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage1_11001_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state3_io)
    begin
                ap_block_pp0_stage1_11001 <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state3_io));
    end process;


    ap_block_pp0_stage1_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state3_io)
    begin
                ap_block_pp0_stage1_subdone <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state3_io));
    end process;

        ap_block_pp0_stage2 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage20_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage20_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage21_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage21_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage22_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage22_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage23_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage23_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage24 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage24_11001_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_RVALID, ap_predicate_op213_read_state26)
    begin
                ap_block_pp0_stage24_11001 <= ((ap_predicate_op213_read_state26 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1));
    end process;


    ap_block_pp0_stage24_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_RVALID, ap_predicate_op213_read_state26)
    begin
                ap_block_pp0_stage24_subdone <= ((ap_predicate_op213_read_state26 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1));
    end process;

        ap_block_pp0_stage25 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage25_11001_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_RVALID, ap_predicate_op216_read_state27)
    begin
                ap_block_pp0_stage25_11001 <= ((ap_predicate_op216_read_state27 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1));
    end process;


    ap_block_pp0_stage25_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_RVALID, ap_predicate_op216_read_state27)
    begin
                ap_block_pp0_stage25_subdone <= ((ap_predicate_op216_read_state27 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1));
    end process;

        ap_block_pp0_stage26 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage26_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage26_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage27 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage27_01001 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage27_11001_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state29_io)
    begin
                ap_block_pp0_stage27_11001 <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state29_io));
    end process;


    ap_block_pp0_stage27_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state29_io)
    begin
                ap_block_pp0_stage27_subdone <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state29_io));
    end process;

        ap_block_pp0_stage28_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage28_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage29_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage29_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage2_11001_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state4_io)
    begin
                ap_block_pp0_stage2_11001 <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state4_io));
    end process;


    ap_block_pp0_stage2_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state4_io)
    begin
                ap_block_pp0_stage2_subdone <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state4_io));
    end process;

        ap_block_pp0_stage3 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage30_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage30_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage31_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage31_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage32 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage32_11001_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_BVALID, ap_predicate_op226_writeresp_state34)
    begin
                ap_block_pp0_stage32_11001 <= ((gmem_BVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op226_writeresp_state34 = ap_const_boolean_1));
    end process;


    ap_block_pp0_stage32_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_BVALID, ap_predicate_op226_writeresp_state34)
    begin
                ap_block_pp0_stage32_subdone <= ((gmem_BVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op226_writeresp_state34 = ap_const_boolean_1));
    end process;

        ap_block_pp0_stage33 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage33_11001_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state35_io)
    begin
                ap_block_pp0_stage33_11001 <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state35_io));
    end process;


    ap_block_pp0_stage33_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state35_io)
    begin
                ap_block_pp0_stage33_subdone <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state35_io));
    end process;

        ap_block_pp0_stage34 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage34_11001_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state36_io)
    begin
                ap_block_pp0_stage34_11001 <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state36_io));
    end process;


    ap_block_pp0_stage34_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state36_io)
    begin
                ap_block_pp0_stage34_subdone <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state36_io));
    end process;

        ap_block_pp0_stage35_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage35_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage36_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage36_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage37_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage37_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage38_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage38_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage39_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage39_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage3_11001_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state5_io)
    begin
                ap_block_pp0_stage3_11001 <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state5_io));
    end process;


    ap_block_pp0_stage3_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state5_io)
    begin
                ap_block_pp0_stage3_subdone <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state5_io));
    end process;

        ap_block_pp0_stage40 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage40_11001_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_RVALID, ap_predicate_op240_read_state42)
    begin
                ap_block_pp0_stage40_11001 <= ((ap_predicate_op240_read_state42 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1));
    end process;


    ap_block_pp0_stage40_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_RVALID, ap_predicate_op240_read_state42)
    begin
                ap_block_pp0_stage40_subdone <= ((ap_predicate_op240_read_state42 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1));
    end process;

        ap_block_pp0_stage41 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage41_11001_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_RVALID, ap_predicate_op243_read_state43)
    begin
                ap_block_pp0_stage41_11001 <= ((ap_predicate_op243_read_state43 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1));
    end process;


    ap_block_pp0_stage41_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_RVALID, ap_predicate_op243_read_state43)
    begin
                ap_block_pp0_stage41_subdone <= ((ap_predicate_op243_read_state43 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1));
    end process;

        ap_block_pp0_stage42 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage42_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage42_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage43 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage43_01001 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage43_11001_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state45_io)
    begin
                ap_block_pp0_stage43_11001 <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state45_io));
    end process;


    ap_block_pp0_stage43_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state45_io)
    begin
                ap_block_pp0_stage43_subdone <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state45_io));
    end process;

        ap_block_pp0_stage44 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage44_01001 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage44_11001_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state46_io)
    begin
                ap_block_pp0_stage44_11001 <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state46_io));
    end process;


    ap_block_pp0_stage44_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state46_io)
    begin
                ap_block_pp0_stage44_subdone <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state46_io));
    end process;

        ap_block_pp0_stage45_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage45_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage46_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage46_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage47_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage47_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage48 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage48_11001_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_BVALID, ap_predicate_op258_writeresp_state50)
    begin
                ap_block_pp0_stage48_11001 <= ((gmem_BVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op258_writeresp_state50 = ap_const_boolean_1));
    end process;


    ap_block_pp0_stage48_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_BVALID, ap_predicate_op258_writeresp_state50)
    begin
                ap_block_pp0_stage48_subdone <= ((gmem_BVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op258_writeresp_state50 = ap_const_boolean_1));
    end process;

        ap_block_pp0_stage49 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage49_11001_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_BVALID, ap_predicate_op261_writeresp_state51, ap_block_state51_io)
    begin
                ap_block_pp0_stage49_11001 <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and ((ap_const_boolean_1 = ap_block_state51_io) or ((gmem_BVALID = ap_const_logic_0) and (ap_predicate_op261_writeresp_state51 = ap_const_boolean_1))));
    end process;


    ap_block_pp0_stage49_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_BVALID, ap_predicate_op261_writeresp_state51, ap_block_state51_io)
    begin
                ap_block_pp0_stage49_subdone <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and ((ap_const_boolean_1 = ap_block_state51_io) or ((gmem_BVALID = ap_const_logic_0) and (ap_predicate_op261_writeresp_state51 = ap_const_boolean_1))));
    end process;

        ap_block_pp0_stage4_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage4_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage50 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage50_11001_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state52_io)
    begin
                ap_block_pp0_stage50_11001 <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state52_io));
    end process;


    ap_block_pp0_stage50_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state52_io)
    begin
                ap_block_pp0_stage50_subdone <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state52_io));
    end process;

        ap_block_pp0_stage51 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage51_11001_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state53_io)
    begin
                ap_block_pp0_stage51_11001 <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state53_io));
    end process;


    ap_block_pp0_stage51_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state53_io)
    begin
                ap_block_pp0_stage51_subdone <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state53_io));
    end process;

        ap_block_pp0_stage52_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage52_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage53_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage53_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage54_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage54_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage55_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage55_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage56 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage56_11001_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_RVALID, ap_predicate_op285_read_state58)
    begin
                ap_block_pp0_stage56_11001 <= ((ap_predicate_op285_read_state58 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1));
    end process;


    ap_block_pp0_stage56_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_RVALID, ap_predicate_op285_read_state58)
    begin
                ap_block_pp0_stage56_subdone <= ((ap_predicate_op285_read_state58 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1));
    end process;

        ap_block_pp0_stage57 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage57_11001_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_RVALID, ap_predicate_op290_read_state59, ap_predicate_op292_read_state59)
    begin
                ap_block_pp0_stage57_11001 <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (((ap_predicate_op292_read_state59 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0)) or ((ap_predicate_op290_read_state59 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0))));
    end process;


    ap_block_pp0_stage57_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_RVALID, ap_predicate_op290_read_state59, ap_predicate_op292_read_state59)
    begin
                ap_block_pp0_stage57_subdone <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (((ap_predicate_op292_read_state59 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0)) or ((ap_predicate_op290_read_state59 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0))));
    end process;

        ap_block_pp0_stage58 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage58_11001_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_RVALID, ap_predicate_op298_read_state60)
    begin
                ap_block_pp0_stage58_11001 <= ((ap_predicate_op298_read_state60 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1));
    end process;


    ap_block_pp0_stage58_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_RVALID, ap_predicate_op298_read_state60)
    begin
                ap_block_pp0_stage58_subdone <= ((ap_predicate_op298_read_state60 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1));
    end process;

        ap_block_pp0_stage59 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage59_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage59_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage5_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage5_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage6 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage60 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage60_01001 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage60_11001_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state62_io)
    begin
                ap_block_pp0_stage60_11001 <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state62_io));
    end process;


    ap_block_pp0_stage60_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state62_io)
    begin
                ap_block_pp0_stage60_subdone <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state62_io));
    end process;

        ap_block_pp0_stage61_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage61_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage62_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage62_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage63_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage63_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage64_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage64_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage65 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage65_11001_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_BVALID, ap_predicate_op308_writeresp_state67)
    begin
                ap_block_pp0_stage65_11001 <= ((gmem_BVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op308_writeresp_state67 = ap_const_boolean_1));
    end process;


    ap_block_pp0_stage65_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_BVALID, ap_predicate_op308_writeresp_state67)
    begin
                ap_block_pp0_stage65_subdone <= ((gmem_BVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op308_writeresp_state67 = ap_const_boolean_1));
    end process;

        ap_block_pp0_stage66 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage66_11001_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state68_io)
    begin
                ap_block_pp0_stage66_11001 <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state68_io));
    end process;


    ap_block_pp0_stage66_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state68_io)
    begin
                ap_block_pp0_stage66_subdone <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state68_io));
    end process;

        ap_block_pp0_stage67 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage67_11001_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state69_io)
    begin
                ap_block_pp0_stage67_11001 <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state69_io));
    end process;


    ap_block_pp0_stage67_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state69_io)
    begin
                ap_block_pp0_stage67_subdone <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state69_io));
    end process;

        ap_block_pp0_stage68_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage68_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage69_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage69_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage6_11001_assign_proc : process(ap_enable_reg_pp0_iter1, gmem_RVALID, ap_predicate_op351_read_state91)
    begin
                ap_block_pp0_stage6_11001 <= ((ap_predicate_op351_read_state91 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter1 = ap_const_logic_1));
    end process;


    ap_block_pp0_stage6_subdone_assign_proc : process(ap_enable_reg_pp0_iter1, gmem_RVALID, ap_predicate_op351_read_state91)
    begin
                ap_block_pp0_stage6_subdone <= ((ap_predicate_op351_read_state91 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter1 = ap_const_logic_1));
    end process;

        ap_block_pp0_stage7 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage70_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage70_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage71_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage71_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage72_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage72_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage73 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage73_11001_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_RVALID, ap_predicate_op322_read_state75)
    begin
                ap_block_pp0_stage73_11001 <= ((ap_predicate_op322_read_state75 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1));
    end process;


    ap_block_pp0_stage73_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_RVALID, ap_predicate_op322_read_state75)
    begin
                ap_block_pp0_stage73_subdone <= ((ap_predicate_op322_read_state75 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1));
    end process;

        ap_block_pp0_stage74 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage74_11001_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_RVALID, ap_predicate_op325_read_state76)
    begin
                ap_block_pp0_stage74_11001 <= ((ap_predicate_op325_read_state76 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1));
    end process;


    ap_block_pp0_stage74_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_RVALID, ap_predicate_op325_read_state76)
    begin
                ap_block_pp0_stage74_subdone <= ((ap_predicate_op325_read_state76 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1));
    end process;

        ap_block_pp0_stage75 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage75_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage75_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage76 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage76_01001 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage76_11001_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state78_io)
    begin
                ap_block_pp0_stage76_11001 <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state78_io));
    end process;


    ap_block_pp0_stage76_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state78_io)
    begin
                ap_block_pp0_stage76_subdone <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state78_io));
    end process;

        ap_block_pp0_stage77_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage77_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage78_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage78_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage79_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage79_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage7_11001_assign_proc : process(ap_enable_reg_pp0_iter1, gmem_RVALID, ap_predicate_op354_read_state92)
    begin
                ap_block_pp0_stage7_11001 <= ((ap_predicate_op354_read_state92 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter1 = ap_const_logic_1));
    end process;


    ap_block_pp0_stage7_subdone_assign_proc : process(ap_enable_reg_pp0_iter1, gmem_RVALID, ap_predicate_op354_read_state92)
    begin
                ap_block_pp0_stage7_subdone <= ((ap_predicate_op354_read_state92 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter1 = ap_const_logic_1));
    end process;

        ap_block_pp0_stage8 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage80_11001 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage80_subdone <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_pp0_stage81 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage81_11001_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_BVALID, ap_predicate_op335_writeresp_state83)
    begin
                ap_block_pp0_stage81_11001 <= ((gmem_BVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op335_writeresp_state83 = ap_const_boolean_1));
    end process;


    ap_block_pp0_stage81_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, gmem_BVALID, ap_predicate_op335_writeresp_state83)
    begin
                ap_block_pp0_stage81_subdone <= ((gmem_BVALID = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op335_writeresp_state83 = ap_const_boolean_1));
    end process;

        ap_block_pp0_stage82 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage82_11001_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state84_io)
    begin
                ap_block_pp0_stage82_11001 <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state84_io));
    end process;


    ap_block_pp0_stage82_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, ap_block_state84_io)
    begin
                ap_block_pp0_stage82_subdone <= ((ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_const_boolean_1 = ap_block_state84_io));
    end process;


    ap_block_pp0_stage8_11001_assign_proc : process(ap_enable_reg_pp0_iter0, icmp_ln1073_reg_676, gmem_RVALID)
    begin
                ap_block_pp0_stage8_11001 <= ((gmem_RVALID = ap_const_logic_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1));
    end process;


    ap_block_pp0_stage8_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, icmp_ln1073_reg_676, gmem_RVALID)
    begin
                ap_block_pp0_stage8_subdone <= ((gmem_RVALID = ap_const_logic_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1));
    end process;

        ap_block_pp0_stage9 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_pp0_stage9_01001_assign_proc : process(ap_enable_reg_pp0_iter0, icmp_ln1073_reg_676, gmem_RVALID)
    begin
                ap_block_pp0_stage9_01001 <= ((gmem_RVALID = ap_const_logic_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1));
    end process;


    ap_block_pp0_stage9_11001_assign_proc : process(ap_enable_reg_pp0_iter0, icmp_ln1073_reg_676, ap_enable_reg_pp0_iter1, gmem_WREADY, gmem_RVALID)
    begin
                ap_block_pp0_stage9_11001 <= (((gmem_WREADY = ap_const_logic_0) and (ap_enable_reg_pp0_iter1 = ap_const_logic_1)) or ((gmem_RVALID = ap_const_logic_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)));
    end process;


    ap_block_pp0_stage9_subdone_assign_proc : process(ap_enable_reg_pp0_iter0, icmp_ln1073_reg_676, ap_enable_reg_pp0_iter1, gmem_WREADY, gmem_RVALID)
    begin
                ap_block_pp0_stage9_subdone <= (((gmem_WREADY = ap_const_logic_0) and (ap_enable_reg_pp0_iter1 = ap_const_logic_1)) or ((gmem_RVALID = ap_const_logic_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)));
    end process;


    ap_block_state10_pp0_stage8_iter0_assign_proc : process(icmp_ln1073_reg_676, gmem_RVALID)
    begin
                ap_block_state10_pp0_stage8_iter0 <= ((gmem_RVALID = ap_const_logic_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_block_state11_pp0_stage9_iter0_assign_proc : process(icmp_ln1073_reg_676, gmem_RVALID)
    begin
                ap_block_state11_pp0_stage9_iter0 <= ((gmem_RVALID = ap_const_logic_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_block_state12_io_assign_proc : process(icmp_ln1073_reg_676, gmem_AWREADY)
    begin
                ap_block_state12_io <= ((gmem_AWREADY = ap_const_logic_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;

        ap_block_state12_pp0_stage10_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_state13_io_assign_proc : process(gmem_WREADY, ap_predicate_op194_write_state13)
    begin
                ap_block_state13_io <= ((gmem_WREADY = ap_const_logic_0) and (ap_predicate_op194_write_state13 = ap_const_boolean_1));
    end process;

        ap_block_state13_pp0_stage11_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state14_pp0_stage12_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state15_pp0_stage13_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state16_pp0_stage14_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state17_pp0_stage15_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_state18_pp0_stage16_iter0_assign_proc : process(gmem_BVALID, ap_predicate_op199_writeresp_state18)
    begin
                ap_block_state18_pp0_stage16_iter0 <= ((gmem_BVALID = ap_const_logic_0) and (ap_predicate_op199_writeresp_state18 = ap_const_boolean_1));
    end process;


    ap_block_state19_io_assign_proc : process(gmem_ARREADY, ap_predicate_op200_readreq_state19)
    begin
                ap_block_state19_io <= ((gmem_ARREADY = ap_const_logic_0) and (ap_predicate_op200_readreq_state19 = ap_const_boolean_1));
    end process;

        ap_block_state19_pp0_stage17_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_state20_io_assign_proc : process(gmem_ARREADY, ap_predicate_op202_readreq_state20)
    begin
                ap_block_state20_io <= ((gmem_ARREADY = ap_const_logic_0) and (ap_predicate_op202_readreq_state20 = ap_const_boolean_1));
    end process;

        ap_block_state20_pp0_stage18_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state21_pp0_stage19_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state22_pp0_stage20_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state23_pp0_stage21_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state24_pp0_stage22_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state25_pp0_stage23_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_state26_pp0_stage24_iter0_assign_proc : process(gmem_RVALID, ap_predicate_op213_read_state26)
    begin
                ap_block_state26_pp0_stage24_iter0 <= ((ap_predicate_op213_read_state26 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0));
    end process;


    ap_block_state27_pp0_stage25_iter0_assign_proc : process(gmem_RVALID, ap_predicate_op216_read_state27)
    begin
                ap_block_state27_pp0_stage25_iter0 <= ((ap_predicate_op216_read_state27 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0));
    end process;

        ap_block_state28_pp0_stage26_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_state29_io_assign_proc : process(gmem_WREADY, ap_predicate_op221_write_state29)
    begin
                ap_block_state29_io <= ((gmem_WREADY = ap_const_logic_0) and (ap_predicate_op221_write_state29 = ap_const_boolean_1));
    end process;

        ap_block_state29_pp0_stage27_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state2_pp0_stage0_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state30_pp0_stage28_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state31_pp0_stage29_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state32_pp0_stage30_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state33_pp0_stage31_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_state34_pp0_stage32_iter0_assign_proc : process(gmem_BVALID, ap_predicate_op226_writeresp_state34)
    begin
                ap_block_state34_pp0_stage32_iter0 <= ((gmem_BVALID = ap_const_logic_0) and (ap_predicate_op226_writeresp_state34 = ap_const_boolean_1));
    end process;


    ap_block_state35_io_assign_proc : process(gmem_ARREADY, ap_predicate_op227_readreq_state35)
    begin
                ap_block_state35_io <= ((gmem_ARREADY = ap_const_logic_0) and (ap_predicate_op227_readreq_state35 = ap_const_boolean_1));
    end process;

        ap_block_state35_pp0_stage33_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_state36_io_assign_proc : process(gmem_ARREADY, ap_predicate_op229_readreq_state36)
    begin
                ap_block_state36_io <= ((gmem_ARREADY = ap_const_logic_0) and (ap_predicate_op229_readreq_state36 = ap_const_boolean_1));
    end process;

        ap_block_state36_pp0_stage34_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state37_pp0_stage35_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state38_pp0_stage36_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state39_pp0_stage37_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_state3_io_assign_proc : process(icmp_ln1073_reg_676, gmem_AWREADY, gmem_ARREADY, ap_predicate_op164_writereq_state3, ap_predicate_op165_writereq_state3)
    begin
                ap_block_state3_io <= (((ap_predicate_op165_writereq_state3 = ap_const_boolean_1) and (gmem_AWREADY = ap_const_logic_0)) or ((ap_predicate_op164_writereq_state3 = ap_const_boolean_1) and (gmem_AWREADY = ap_const_logic_0)) or ((gmem_ARREADY = ap_const_logic_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1)));
    end process;

        ap_block_state3_pp0_stage1_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state40_pp0_stage38_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state41_pp0_stage39_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_state42_pp0_stage40_iter0_assign_proc : process(gmem_RVALID, ap_predicate_op240_read_state42)
    begin
                ap_block_state42_pp0_stage40_iter0 <= ((ap_predicate_op240_read_state42 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0));
    end process;


    ap_block_state43_pp0_stage41_iter0_assign_proc : process(gmem_RVALID, ap_predicate_op243_read_state43)
    begin
                ap_block_state43_pp0_stage41_iter0 <= ((ap_predicate_op243_read_state43 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0));
    end process;

        ap_block_state44_pp0_stage42_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_state45_io_assign_proc : process(gmem_WREADY, ap_predicate_op248_write_state45)
    begin
                ap_block_state45_io <= ((gmem_WREADY = ap_const_logic_0) and (ap_predicate_op248_write_state45 = ap_const_boolean_1));
    end process;

        ap_block_state45_pp0_stage43_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_state46_io_assign_proc : process(gmem_WREADY, ap_predicate_op251_write_state46)
    begin
                ap_block_state46_io <= ((gmem_WREADY = ap_const_logic_0) and (ap_predicate_op251_write_state46 = ap_const_boolean_1));
    end process;

        ap_block_state46_pp0_stage44_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state47_pp0_stage45_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state48_pp0_stage46_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state49_pp0_stage47_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_state4_io_assign_proc : process(icmp_ln1073_reg_676, gmem_AWREADY, gmem_ARREADY, ap_predicate_op170_writereq_state4, ap_predicate_op171_writereq_state4)
    begin
                ap_block_state4_io <= (((ap_predicate_op171_writereq_state4 = ap_const_boolean_1) and (gmem_AWREADY = ap_const_logic_0)) or ((ap_predicate_op170_writereq_state4 = ap_const_boolean_1) and (gmem_AWREADY = ap_const_logic_0)) or ((gmem_ARREADY = ap_const_logic_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1)));
    end process;

        ap_block_state4_pp0_stage2_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_state50_pp0_stage48_iter0_assign_proc : process(gmem_BVALID, ap_predicate_op258_writeresp_state50)
    begin
                ap_block_state50_pp0_stage48_iter0 <= ((gmem_BVALID = ap_const_logic_0) and (ap_predicate_op258_writeresp_state50 = ap_const_boolean_1));
    end process;


    ap_block_state51_io_assign_proc : process(gmem_ARREADY, ap_predicate_op260_readreq_state51)
    begin
                ap_block_state51_io <= ((gmem_ARREADY = ap_const_logic_0) and (ap_predicate_op260_readreq_state51 = ap_const_boolean_1));
    end process;


    ap_block_state51_pp0_stage49_iter0_assign_proc : process(gmem_BVALID, ap_predicate_op261_writeresp_state51)
    begin
                ap_block_state51_pp0_stage49_iter0 <= ((gmem_BVALID = ap_const_logic_0) and (ap_predicate_op261_writeresp_state51 = ap_const_boolean_1));
    end process;


    ap_block_state52_io_assign_proc : process(gmem_ARREADY, ap_predicate_op263_readreq_state52, ap_predicate_op264_readreq_state52)
    begin
                ap_block_state52_io <= (((gmem_ARREADY = ap_const_logic_0) and (ap_predicate_op264_readreq_state52 = ap_const_boolean_1)) or ((gmem_ARREADY = ap_const_logic_0) and (ap_predicate_op263_readreq_state52 = ap_const_boolean_1)));
    end process;

        ap_block_state52_pp0_stage50_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_state53_io_assign_proc : process(gmem_ARREADY, ap_predicate_op268_readreq_state53)
    begin
                ap_block_state53_io <= ((gmem_ARREADY = ap_const_logic_0) and (ap_predicate_op268_readreq_state53 = ap_const_boolean_1));
    end process;

        ap_block_state53_pp0_stage51_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state54_pp0_stage52_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state55_pp0_stage53_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state56_pp0_stage54_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state57_pp0_stage55_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_state58_pp0_stage56_iter0_assign_proc : process(gmem_RVALID, ap_predicate_op285_read_state58)
    begin
                ap_block_state58_pp0_stage56_iter0 <= ((ap_predicate_op285_read_state58 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0));
    end process;


    ap_block_state59_pp0_stage57_iter0_assign_proc : process(gmem_RVALID, ap_predicate_op290_read_state59, ap_predicate_op292_read_state59)
    begin
                ap_block_state59_pp0_stage57_iter0 <= (((ap_predicate_op292_read_state59 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0)) or ((ap_predicate_op290_read_state59 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0)));
    end process;


    ap_block_state5_io_assign_proc : process(gmem_AWREADY, ap_predicate_op174_writereq_state5, ap_predicate_op175_writereq_state5)
    begin
                ap_block_state5_io <= (((gmem_AWREADY = ap_const_logic_0) and (ap_predicate_op175_writereq_state5 = ap_const_boolean_1)) or ((gmem_AWREADY = ap_const_logic_0) and (ap_predicate_op174_writereq_state5 = ap_const_boolean_1)));
    end process;

        ap_block_state5_pp0_stage3_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_state60_pp0_stage58_iter0_assign_proc : process(gmem_RVALID, ap_predicate_op298_read_state60)
    begin
                ap_block_state60_pp0_stage58_iter0 <= ((ap_predicate_op298_read_state60 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0));
    end process;

        ap_block_state61_pp0_stage59_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_state62_io_assign_proc : process(gmem_WREADY, ap_predicate_op303_write_state62)
    begin
                ap_block_state62_io <= ((gmem_WREADY = ap_const_logic_0) and (ap_predicate_op303_write_state62 = ap_const_boolean_1));
    end process;

        ap_block_state62_pp0_stage60_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state63_pp0_stage61_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state64_pp0_stage62_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state65_pp0_stage63_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state66_pp0_stage64_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_state67_pp0_stage65_iter0_assign_proc : process(gmem_BVALID, ap_predicate_op308_writeresp_state67)
    begin
                ap_block_state67_pp0_stage65_iter0 <= ((gmem_BVALID = ap_const_logic_0) and (ap_predicate_op308_writeresp_state67 = ap_const_boolean_1));
    end process;


    ap_block_state68_io_assign_proc : process(gmem_ARREADY, ap_predicate_op309_readreq_state68)
    begin
                ap_block_state68_io <= ((gmem_ARREADY = ap_const_logic_0) and (ap_predicate_op309_readreq_state68 = ap_const_boolean_1));
    end process;

        ap_block_state68_pp0_stage66_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_state69_io_assign_proc : process(gmem_ARREADY, ap_predicate_op311_readreq_state69)
    begin
                ap_block_state69_io <= ((gmem_ARREADY = ap_const_logic_0) and (ap_predicate_op311_readreq_state69 = ap_const_boolean_1));
    end process;

        ap_block_state69_pp0_stage67_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state6_pp0_stage4_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state70_pp0_stage68_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state71_pp0_stage69_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state72_pp0_stage70_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state73_pp0_stage71_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state74_pp0_stage72_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_state75_pp0_stage73_iter0_assign_proc : process(gmem_RVALID, ap_predicate_op322_read_state75)
    begin
                ap_block_state75_pp0_stage73_iter0 <= ((ap_predicate_op322_read_state75 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0));
    end process;


    ap_block_state76_pp0_stage74_iter0_assign_proc : process(gmem_RVALID, ap_predicate_op325_read_state76)
    begin
                ap_block_state76_pp0_stage74_iter0 <= ((ap_predicate_op325_read_state76 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0));
    end process;

        ap_block_state77_pp0_stage75_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_state78_io_assign_proc : process(gmem_WREADY, ap_predicate_op330_write_state78)
    begin
                ap_block_state78_io <= ((gmem_WREADY = ap_const_logic_0) and (ap_predicate_op330_write_state78 = ap_const_boolean_1));
    end process;

        ap_block_state78_pp0_stage76_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state79_pp0_stage77_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state7_pp0_stage5_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state80_pp0_stage78_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state81_pp0_stage79_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state82_pp0_stage80_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_state83_pp0_stage81_iter0_assign_proc : process(gmem_BVALID, ap_predicate_op335_writeresp_state83)
    begin
                ap_block_state83_pp0_stage81_iter0 <= ((gmem_BVALID = ap_const_logic_0) and (ap_predicate_op335_writeresp_state83 = ap_const_boolean_1));
    end process;


    ap_block_state84_io_assign_proc : process(gmem_ARREADY, ap_predicate_op336_readreq_state84)
    begin
                ap_block_state84_io <= ((gmem_ARREADY = ap_const_logic_0) and (ap_predicate_op336_readreq_state84 = ap_const_boolean_1));
    end process;

        ap_block_state84_pp0_stage82_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_state85_io_assign_proc : process(gmem_ARREADY, ap_predicate_op340_readreq_state85)
    begin
                ap_block_state85_io <= ((ap_predicate_op340_readreq_state85 = ap_const_boolean_1) and (gmem_ARREADY = ap_const_logic_0));
    end process;

        ap_block_state85_pp0_stage0_iter1 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state86_pp0_stage1_iter1 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state87_pp0_stage2_iter1 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state88_pp0_stage3_iter1 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state89_pp0_stage4_iter1 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state8_pp0_stage6_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state90_pp0_stage5_iter1 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_state91_pp0_stage6_iter1_assign_proc : process(gmem_RVALID, ap_predicate_op351_read_state91)
    begin
                ap_block_state91_pp0_stage6_iter1 <= ((ap_predicate_op351_read_state91 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0));
    end process;


    ap_block_state92_pp0_stage7_iter1_assign_proc : process(gmem_RVALID, ap_predicate_op354_read_state92)
    begin
                ap_block_state92_pp0_stage7_iter1 <= ((ap_predicate_op354_read_state92 = ap_const_boolean_1) and (gmem_RVALID = ap_const_logic_0));
    end process;

        ap_block_state93_pp0_stage8_iter1 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state94_pp0_stage9_iter1 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state95_pp0_stage10_iter1 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state96_pp0_stage11_iter1 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state97_pp0_stage12_iter1 <= not((ap_const_boolean_1 = ap_const_boolean_1));
        ap_block_state98_pp0_stage13_iter1 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_block_state99_pp0_stage14_iter1_assign_proc : process(gmem_BVALID)
    begin
                ap_block_state99_pp0_stage14_iter1 <= (gmem_BVALID = ap_const_logic_0);
    end process;

        ap_block_state9_pp0_stage7_iter0 <= not((ap_const_boolean_1 = ap_const_boolean_1));

    ap_condition_pp0_exit_iter0_state2_assign_proc : process(icmp_ln1073_fu_364_p2)
    begin
        if ((icmp_ln1073_fu_364_p2 = ap_const_lv1_0)) then 
            ap_condition_pp0_exit_iter0_state2 <= ap_const_logic_1;
        else 
            ap_condition_pp0_exit_iter0_state2 <= ap_const_logic_0;
        end if; 
    end process;


    ap_done_assign_proc : process(ap_CS_fsm_state100)
    begin
        if ((ap_const_logic_1 = ap_CS_fsm_state100)) then 
            ap_done <= ap_const_logic_1;
        else 
            ap_done <= ap_const_logic_0;
        end if; 
    end process;

    ap_enable_pp0 <= (ap_idle_pp0 xor ap_const_logic_1);

    ap_idle_assign_proc : process(ap_start, ap_CS_fsm_state1)
    begin
        if (((ap_start = ap_const_logic_0) and (ap_const_logic_1 = ap_CS_fsm_state1))) then 
            ap_idle <= ap_const_logic_1;
        else 
            ap_idle <= ap_const_logic_0;
        end if; 
    end process;


    ap_idle_pp0_assign_proc : process(ap_enable_reg_pp0_iter0, ap_enable_reg_pp0_iter1)
    begin
        if (((ap_enable_reg_pp0_iter1 = ap_const_logic_0) and (ap_enable_reg_pp0_iter0 = ap_const_logic_0))) then 
            ap_idle_pp0 <= ap_const_logic_1;
        else 
            ap_idle_pp0 <= ap_const_logic_0;
        end if; 
    end process;


    ap_predicate_op164_writereq_state3_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op164_writereq_state3 <= ((op_read_reg_640 = ap_const_lv1_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op165_writereq_state3_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op165_writereq_state3 <= ((op_read_reg_640 = ap_const_lv1_1) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op170_writereq_state4_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op170_writereq_state4 <= ((op_read_reg_640 = ap_const_lv1_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op171_writereq_state4_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op171_writereq_state4 <= ((op_read_reg_640 = ap_const_lv1_1) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op174_writereq_state5_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op174_writereq_state5 <= ((op_read_reg_640 = ap_const_lv1_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op175_writereq_state5_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op175_writereq_state5 <= ((op_read_reg_640 = ap_const_lv1_1) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op194_write_state13_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op194_write_state13 <= ((op_read_reg_640 = ap_const_lv1_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op199_writeresp_state18_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op199_writeresp_state18 <= ((op_read_reg_640 = ap_const_lv1_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op200_readreq_state19_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op200_readreq_state19 <= ((op_read_reg_640 = ap_const_lv1_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op202_readreq_state20_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op202_readreq_state20 <= ((op_read_reg_640 = ap_const_lv1_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op213_read_state26_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op213_read_state26 <= ((op_read_reg_640 = ap_const_lv1_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op216_read_state27_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op216_read_state27 <= ((op_read_reg_640 = ap_const_lv1_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op221_write_state29_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op221_write_state29 <= ((op_read_reg_640 = ap_const_lv1_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op226_writeresp_state34_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op226_writeresp_state34 <= ((op_read_reg_640 = ap_const_lv1_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op227_readreq_state35_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op227_readreq_state35 <= ((op_read_reg_640 = ap_const_lv1_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op229_readreq_state36_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op229_readreq_state36 <= ((op_read_reg_640 = ap_const_lv1_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op240_read_state42_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op240_read_state42 <= ((op_read_reg_640 = ap_const_lv1_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op243_read_state43_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op243_read_state43 <= ((op_read_reg_640 = ap_const_lv1_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op248_write_state45_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op248_write_state45 <= ((op_read_reg_640 = ap_const_lv1_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op251_write_state46_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op251_write_state46 <= ((op_read_reg_640 = ap_const_lv1_1) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op258_writeresp_state50_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op258_writeresp_state50 <= ((op_read_reg_640 = ap_const_lv1_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op260_readreq_state51_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op260_readreq_state51 <= ((op_read_reg_640 = ap_const_lv1_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op261_writeresp_state51_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op261_writeresp_state51 <= ((op_read_reg_640 = ap_const_lv1_1) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op263_readreq_state52_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op263_readreq_state52 <= ((op_read_reg_640 = ap_const_lv1_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op264_readreq_state52_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op264_readreq_state52 <= ((op_read_reg_640 = ap_const_lv1_1) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op268_readreq_state53_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op268_readreq_state53 <= ((op_read_reg_640 = ap_const_lv1_1) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op285_read_state58_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op285_read_state58 <= ((op_read_reg_640 = ap_const_lv1_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op290_read_state59_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op290_read_state59 <= ((op_read_reg_640 = ap_const_lv1_0) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op292_read_state59_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op292_read_state59 <= ((op_read_reg_640 = ap_const_lv1_1) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op298_read_state60_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op298_read_state60 <= ((op_read_reg_640 = ap_const_lv1_1) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op303_write_state62_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op303_write_state62 <= ((op_read_reg_640 = ap_const_lv1_1) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op308_writeresp_state67_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op308_writeresp_state67 <= ((op_read_reg_640 = ap_const_lv1_1) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op309_readreq_state68_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op309_readreq_state68 <= ((op_read_reg_640 = ap_const_lv1_1) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op311_readreq_state69_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op311_readreq_state69 <= ((op_read_reg_640 = ap_const_lv1_1) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op322_read_state75_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op322_read_state75 <= ((op_read_reg_640 = ap_const_lv1_1) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op325_read_state76_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op325_read_state76 <= ((op_read_reg_640 = ap_const_lv1_1) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op330_write_state78_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op330_write_state78 <= ((op_read_reg_640 = ap_const_lv1_1) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op335_writeresp_state83_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op335_writeresp_state83 <= ((op_read_reg_640 = ap_const_lv1_1) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op336_readreq_state84_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op336_readreq_state84 <= ((op_read_reg_640 = ap_const_lv1_1) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op340_readreq_state85_assign_proc : process(icmp_ln1073_reg_676, op_read_reg_640)
    begin
                ap_predicate_op340_readreq_state85 <= ((op_read_reg_640 = ap_const_lv1_1) and (icmp_ln1073_reg_676 = ap_const_lv1_1));
    end process;


    ap_predicate_op351_read_state91_assign_proc : process(op_read_reg_640, icmp_ln1073_reg_676_pp0_iter1_reg)
    begin
                ap_predicate_op351_read_state91 <= ((icmp_ln1073_reg_676_pp0_iter1_reg = ap_const_lv1_1) and (op_read_reg_640 = ap_const_lv1_1));
    end process;


    ap_predicate_op354_read_state92_assign_proc : process(op_read_reg_640, icmp_ln1073_reg_676_pp0_iter1_reg)
    begin
                ap_predicate_op354_read_state92 <= ((icmp_ln1073_reg_676_pp0_iter1_reg = ap_const_lv1_1) and (op_read_reg_640 = ap_const_lv1_1));
    end process;


    ap_ready_assign_proc : process(ap_CS_fsm_state100)
    begin
        if ((ap_const_logic_1 = ap_CS_fsm_state100)) then 
            ap_ready <= ap_const_logic_1;
        else 
            ap_ready <= ap_const_logic_0;
        end if; 
    end process;


    ap_rst_n_inv_assign_proc : process(ap_rst_n)
    begin
                ap_rst_n_inv <= not(ap_rst_n);
    end process;


    gmem_ARADDR_assign_proc : process(ap_CS_fsm_pp0_stage1, ap_enable_reg_pp0_iter0, icmp_ln1073_reg_676, ap_CS_fsm_pp0_stage50, ap_CS_fsm_pp0_stage66, ap_CS_fsm_pp0_stage82, ap_enable_reg_pp0_iter1, ap_CS_fsm_pp0_stage17, ap_CS_fsm_pp0_stage33, ap_CS_fsm_pp0_stage49, ap_CS_fsm_pp0_stage2, ap_CS_fsm_pp0_stage51, ap_CS_fsm_pp0_stage67, ap_CS_fsm_pp0_stage0, ap_CS_fsm_pp0_stage18, ap_CS_fsm_pp0_stage34, ap_predicate_op340_readreq_state85, ap_block_pp0_stage0_11001, gmem_addr_reg_695, ap_block_pp0_stage1_11001, gmem_addr_1_reg_713, ap_block_pp0_stage2_11001, ap_predicate_op336_readreq_state84, ap_block_pp0_stage82_11001, sext_ln357_fu_469_p1, sext_ln357_1_fu_489_p1, ap_predicate_op200_readreq_state19, ap_block_pp0_stage17_11001, ap_predicate_op227_readreq_state35, ap_block_pp0_stage33_11001, ap_predicate_op260_readreq_state51, ap_block_pp0_stage49_11001, ap_predicate_op263_readreq_state52, ap_predicate_op264_readreq_state52, ap_block_pp0_stage50_11001, ap_predicate_op309_readreq_state68, ap_block_pp0_stage66_11001, ap_predicate_op202_readreq_state20, ap_block_pp0_stage18_11001, ap_predicate_op229_readreq_state36, ap_block_pp0_stage34_11001, ap_predicate_op268_readreq_state53, ap_block_pp0_stage51_11001, ap_predicate_op311_readreq_state69, ap_block_pp0_stage67_11001)
    begin
        if ((((ap_predicate_op340_readreq_state85 = ap_const_boolean_1) and (ap_enable_reg_pp0_iter1 = ap_const_logic_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0) and (ap_const_boolean_0 = ap_block_pp0_stage0_11001)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage34) and (ap_const_boolean_0 = ap_block_pp0_stage34_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op229_readreq_state36 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage18) and (ap_const_boolean_0 = ap_block_pp0_stage18_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op202_readreq_state20 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage67) and (ap_const_boolean_0 = ap_block_pp0_stage67_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op311_readreq_state69 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage51) and (ap_const_boolean_0 = ap_block_pp0_stage51_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op268_readreq_state53 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage50) and (ap_const_boolean_0 = ap_block_pp0_stage50_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op263_readreq_state52 = ap_const_boolean_1)))) then 
            gmem_ARADDR <= gmem_addr_1_reg_713;
        elsif (((ap_const_logic_1 = ap_CS_fsm_pp0_stage2) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage2_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1))) then 
            gmem_ARADDR <= sext_ln357_1_fu_489_p1;
        elsif ((((ap_const_logic_1 = ap_CS_fsm_pp0_stage49) and (ap_const_boolean_0 = ap_block_pp0_stage49_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op260_readreq_state51 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage33) and (ap_const_boolean_0 = ap_block_pp0_stage33_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op227_readreq_state35 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage17) and (ap_const_boolean_0 = ap_block_pp0_stage17_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op200_readreq_state19 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage82) and (ap_const_boolean_0 = ap_block_pp0_stage82_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op336_readreq_state84 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage66) and (ap_const_boolean_0 = ap_block_pp0_stage66_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op309_readreq_state68 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage50) and (ap_const_boolean_0 = ap_block_pp0_stage50_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op264_readreq_state52 = ap_const_boolean_1)))) then 
            gmem_ARADDR <= gmem_addr_reg_695;
        elsif (((ap_const_logic_1 = ap_CS_fsm_pp0_stage1) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage1_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1))) then 
            gmem_ARADDR <= sext_ln357_fu_469_p1;
        else 
            gmem_ARADDR <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
        end if; 
    end process;


    gmem_ARVALID_assign_proc : process(ap_CS_fsm_pp0_stage1, ap_enable_reg_pp0_iter0, icmp_ln1073_reg_676, ap_CS_fsm_pp0_stage50, ap_CS_fsm_pp0_stage66, ap_CS_fsm_pp0_stage82, ap_enable_reg_pp0_iter1, ap_CS_fsm_pp0_stage17, ap_CS_fsm_pp0_stage33, ap_CS_fsm_pp0_stage49, ap_CS_fsm_pp0_stage2, ap_CS_fsm_pp0_stage51, ap_CS_fsm_pp0_stage67, ap_CS_fsm_pp0_stage0, ap_CS_fsm_pp0_stage18, ap_CS_fsm_pp0_stage34, ap_predicate_op340_readreq_state85, ap_block_pp0_stage0_11001, ap_block_pp0_stage1_11001, ap_block_pp0_stage2_11001, ap_predicate_op336_readreq_state84, ap_block_pp0_stage82_11001, ap_predicate_op200_readreq_state19, ap_block_pp0_stage17_11001, ap_predicate_op227_readreq_state35, ap_block_pp0_stage33_11001, ap_predicate_op260_readreq_state51, ap_block_pp0_stage49_11001, ap_predicate_op263_readreq_state52, ap_predicate_op264_readreq_state52, ap_block_pp0_stage50_11001, ap_predicate_op309_readreq_state68, ap_block_pp0_stage66_11001, ap_predicate_op202_readreq_state20, ap_block_pp0_stage18_11001, ap_predicate_op229_readreq_state36, ap_block_pp0_stage34_11001, ap_predicate_op268_readreq_state53, ap_block_pp0_stage51_11001, ap_predicate_op311_readreq_state69, ap_block_pp0_stage67_11001)
    begin
        if ((((ap_predicate_op340_readreq_state85 = ap_const_boolean_1) and (ap_enable_reg_pp0_iter1 = ap_const_logic_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0) and (ap_const_boolean_0 = ap_block_pp0_stage0_11001)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage34) and (ap_const_boolean_0 = ap_block_pp0_stage34_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op229_readreq_state36 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage18) and (ap_const_boolean_0 = ap_block_pp0_stage18_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op202_readreq_state20 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage67) and (ap_const_boolean_0 = ap_block_pp0_stage67_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op311_readreq_state69 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage51) and (ap_const_boolean_0 = ap_block_pp0_stage51_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op268_readreq_state53 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage2) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage2_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage49) and (ap_const_boolean_0 = ap_block_pp0_stage49_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op260_readreq_state51 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage33) and (ap_const_boolean_0 = ap_block_pp0_stage33_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op227_readreq_state35 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage17) and (ap_const_boolean_0 = ap_block_pp0_stage17_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op200_readreq_state19 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage82) and (ap_const_boolean_0 = ap_block_pp0_stage82_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op336_readreq_state84 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage66) and (ap_const_boolean_0 = ap_block_pp0_stage66_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op309_readreq_state68 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage50) and (ap_const_boolean_0 = ap_block_pp0_stage50_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op264_readreq_state52 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage50) and (ap_const_boolean_0 = ap_block_pp0_stage50_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op263_readreq_state52 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage1) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage1_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)))) then 
            gmem_ARVALID <= ap_const_logic_1;
        else 
            gmem_ARVALID <= ap_const_logic_0;
        end if; 
    end process;


    gmem_AWADDR_assign_proc : process(ap_CS_fsm_pp0_stage1, ap_enable_reg_pp0_iter0, icmp_ln1073_reg_676, ap_CS_fsm_pp0_stage2, ap_CS_fsm_pp0_stage3, ap_CS_fsm_pp0_stage10, ap_predicate_op164_writereq_state3, ap_predicate_op165_writereq_state3, ap_block_pp0_stage1_11001, gmem_addr_2_reg_701, ap_predicate_op170_writereq_state4, ap_predicate_op171_writereq_state4, ap_block_pp0_stage2_11001, ap_block_pp0_stage10_11001, sext_ln414_fu_479_p1, ap_predicate_op174_writereq_state5, ap_predicate_op175_writereq_state5, ap_block_pp0_stage3_11001)
    begin
        if ((((ap_predicate_op171_writereq_state4 = ap_const_boolean_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage2) and (ap_const_boolean_0 = ap_block_pp0_stage2_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((ap_predicate_op170_writereq_state4 = ap_const_boolean_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage2) and (ap_const_boolean_0 = ap_block_pp0_stage2_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage10) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage10_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage3) and (ap_const_boolean_0 = ap_block_pp0_stage3_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op175_writereq_state5 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage3) and (ap_const_boolean_0 = ap_block_pp0_stage3_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op174_writereq_state5 = ap_const_boolean_1)))) then 
            gmem_AWADDR <= gmem_addr_2_reg_701;
        elsif ((((ap_predicate_op165_writereq_state3 = ap_const_boolean_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage1) and (ap_const_boolean_0 = ap_block_pp0_stage1_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((ap_predicate_op164_writereq_state3 = ap_const_boolean_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage1) and (ap_const_boolean_0 = ap_block_pp0_stage1_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)))) then 
            gmem_AWADDR <= sext_ln414_fu_479_p1;
        else 
            gmem_AWADDR <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
        end if; 
    end process;


    gmem_AWVALID_assign_proc : process(ap_CS_fsm_pp0_stage1, ap_enable_reg_pp0_iter0, icmp_ln1073_reg_676, ap_CS_fsm_pp0_stage2, ap_CS_fsm_pp0_stage3, ap_CS_fsm_pp0_stage10, ap_predicate_op164_writereq_state3, ap_predicate_op165_writereq_state3, ap_block_pp0_stage1_11001, ap_predicate_op170_writereq_state4, ap_predicate_op171_writereq_state4, ap_block_pp0_stage2_11001, ap_block_pp0_stage10_11001, ap_predicate_op174_writereq_state5, ap_predicate_op175_writereq_state5, ap_block_pp0_stage3_11001)
    begin
        if ((((ap_predicate_op171_writereq_state4 = ap_const_boolean_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage2) and (ap_const_boolean_0 = ap_block_pp0_stage2_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((ap_predicate_op170_writereq_state4 = ap_const_boolean_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage2) and (ap_const_boolean_0 = ap_block_pp0_stage2_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((ap_predicate_op165_writereq_state3 = ap_const_boolean_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage1) and (ap_const_boolean_0 = ap_block_pp0_stage1_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((ap_predicate_op164_writereq_state3 = ap_const_boolean_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage1) and (ap_const_boolean_0 = ap_block_pp0_stage1_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage10) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage10_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage3) and (ap_const_boolean_0 = ap_block_pp0_stage3_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op175_writereq_state5 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage3) and (ap_const_boolean_0 = ap_block_pp0_stage3_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op174_writereq_state5 = ap_const_boolean_1)))) then 
            gmem_AWVALID <= ap_const_logic_1;
        else 
            gmem_AWVALID <= ap_const_logic_0;
        end if; 
    end process;


    gmem_BREADY_assign_proc : process(ap_enable_reg_pp0_iter0, ap_enable_reg_pp0_iter1, ap_CS_fsm_pp0_stage49, ap_CS_fsm_pp0_stage65, ap_CS_fsm_pp0_stage81, ap_CS_fsm_pp0_stage16, ap_CS_fsm_pp0_stage32, ap_CS_fsm_pp0_stage48, ap_CS_fsm_pp0_stage14, ap_predicate_op261_writeresp_state51, ap_block_pp0_stage49_11001, ap_predicate_op199_writeresp_state18, ap_block_pp0_stage16_11001, ap_predicate_op226_writeresp_state34, ap_block_pp0_stage32_11001, ap_predicate_op258_writeresp_state50, ap_block_pp0_stage48_11001, ap_predicate_op308_writeresp_state67, ap_block_pp0_stage65_11001, ap_predicate_op335_writeresp_state83, ap_block_pp0_stage81_11001, ap_block_pp0_stage14_11001)
    begin
        if ((((ap_const_logic_1 = ap_CS_fsm_pp0_stage48) and (ap_const_boolean_0 = ap_block_pp0_stage48_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op258_writeresp_state50 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage32) and (ap_const_boolean_0 = ap_block_pp0_stage32_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op226_writeresp_state34 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage16) and (ap_const_boolean_0 = ap_block_pp0_stage16_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op199_writeresp_state18 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage81) and (ap_const_boolean_0 = ap_block_pp0_stage81_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op335_writeresp_state83 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage65) and (ap_const_boolean_0 = ap_block_pp0_stage65_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op308_writeresp_state67 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage49) and (ap_const_boolean_0 = ap_block_pp0_stage49_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op261_writeresp_state51 = ap_const_boolean_1)) or ((ap_enable_reg_pp0_iter1 = ap_const_logic_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage14) and (ap_const_boolean_0 = ap_block_pp0_stage14_11001)))) then 
            gmem_BREADY <= ap_const_logic_1;
        else 
            gmem_BREADY <= ap_const_logic_0;
        end if; 
    end process;


    gmem_RREADY_assign_proc : process(ap_enable_reg_pp0_iter0, icmp_ln1073_reg_676, ap_CS_fsm_pp0_stage8, ap_CS_fsm_pp0_stage57, ap_CS_fsm_pp0_stage73, ap_CS_fsm_pp0_stage6, ap_enable_reg_pp0_iter1, ap_CS_fsm_pp0_stage24, ap_CS_fsm_pp0_stage40, ap_CS_fsm_pp0_stage56, ap_CS_fsm_pp0_stage9, ap_CS_fsm_pp0_stage58, ap_CS_fsm_pp0_stage74, ap_CS_fsm_pp0_stage7, ap_CS_fsm_pp0_stage25, ap_CS_fsm_pp0_stage41, ap_predicate_op213_read_state26, ap_block_pp0_stage24_11001, ap_predicate_op290_read_state59, ap_predicate_op292_read_state59, ap_block_pp0_stage57_11001, ap_predicate_op216_read_state27, ap_block_pp0_stage25_11001, ap_predicate_op298_read_state60, ap_block_pp0_stage58_11001, ap_predicate_op240_read_state42, ap_block_pp0_stage40_11001, ap_predicate_op322_read_state75, ap_block_pp0_stage73_11001, ap_predicate_op243_read_state43, ap_block_pp0_stage41_11001, ap_predicate_op325_read_state76, ap_block_pp0_stage74_11001, ap_predicate_op285_read_state58, ap_block_pp0_stage56_11001, ap_predicate_op351_read_state91, ap_block_pp0_stage6_11001, ap_predicate_op354_read_state92, ap_block_pp0_stage7_11001, ap_block_pp0_stage8_11001, ap_block_pp0_stage9_11001)
    begin
        if ((((ap_predicate_op354_read_state92 = ap_const_boolean_1) and (ap_enable_reg_pp0_iter1 = ap_const_logic_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage7) and (ap_const_boolean_0 = ap_block_pp0_stage7_11001)) or ((ap_predicate_op351_read_state91 = ap_const_boolean_1) and (ap_enable_reg_pp0_iter1 = ap_const_logic_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage6) and (ap_const_boolean_0 = ap_block_pp0_stage6_11001)) or ((ap_predicate_op285_read_state58 = ap_const_boolean_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage56) and (ap_const_boolean_0 = ap_block_pp0_stage56_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((ap_predicate_op325_read_state76 = ap_const_boolean_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage74) and (ap_const_boolean_0 = ap_block_pp0_stage74_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((ap_predicate_op243_read_state43 = ap_const_boolean_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage41) and (ap_const_boolean_0 = ap_block_pp0_stage41_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((ap_predicate_op322_read_state75 = ap_const_boolean_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage73) and (ap_const_boolean_0 = ap_block_pp0_stage73_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((ap_predicate_op240_read_state42 = ap_const_boolean_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage40) and (ap_const_boolean_0 = ap_block_pp0_stage40_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((ap_predicate_op298_read_state60 = ap_const_boolean_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage58) and (ap_const_boolean_0 = ap_block_pp0_stage58_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((ap_predicate_op216_read_state27 = ap_const_boolean_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage25) and (ap_const_boolean_0 = ap_block_pp0_stage25_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((ap_predicate_op292_read_state59 = ap_const_boolean_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage57) and (ap_const_boolean_0 = ap_block_pp0_stage57_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((ap_predicate_op290_read_state59 = ap_const_boolean_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage57) and (ap_const_boolean_0 = ap_block_pp0_stage57_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((ap_predicate_op213_read_state26 = ap_const_boolean_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage24) and (ap_const_boolean_0 = ap_block_pp0_stage24_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage9) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage9_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage8) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage8_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)))) then 
            gmem_RREADY <= ap_const_logic_1;
        else 
            gmem_RREADY <= ap_const_logic_0;
        end if; 
    end process;


    gmem_WDATA_assign_proc : process(ap_enable_reg_pp0_iter0, ap_enable_reg_pp0_iter1, ap_CS_fsm_pp0_stage9, ap_CS_fsm_pp0_stage44, ap_CS_fsm_pp0_stage60, ap_CS_fsm_pp0_stage76, ap_CS_fsm_pp0_stage11, ap_CS_fsm_pp0_stage27, ap_CS_fsm_pp0_stage43, ap_phi_reg_pp0_iter1_storemerge_reg_250, ap_predicate_op194_write_state13, p_Result_11_fu_515_p1, ap_block_pp0_stage11_01001, ap_predicate_op221_write_state29, p_Result_12_fu_531_p1, ap_block_pp0_stage27_01001, ap_predicate_op248_write_state45, p_Result_13_fu_549_p1, ap_block_pp0_stage43_01001, ap_predicate_op251_write_state46, p_Result_8_fu_554_p1, ap_block_pp0_stage44_01001, ap_predicate_op303_write_state62, p_Result_9_fu_585_p1, ap_block_pp0_stage60_01001, ap_predicate_op330_write_state78, p_Result_10_fu_603_p1, ap_block_pp0_stage76_01001, ap_block_pp0_stage9_01001)
    begin
        if (((ap_enable_reg_pp0_iter1 = ap_const_logic_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage9) and (ap_const_boolean_0 = ap_block_pp0_stage9_01001))) then 
            gmem_WDATA <= ap_phi_reg_pp0_iter1_storemerge_reg_250;
        elsif (((ap_const_logic_1 = ap_CS_fsm_pp0_stage76) and (ap_const_boolean_0 = ap_block_pp0_stage76_01001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op330_write_state78 = ap_const_boolean_1))) then 
            gmem_WDATA <= p_Result_10_fu_603_p1;
        elsif (((ap_const_logic_1 = ap_CS_fsm_pp0_stage60) and (ap_const_boolean_0 = ap_block_pp0_stage60_01001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op303_write_state62 = ap_const_boolean_1))) then 
            gmem_WDATA <= p_Result_9_fu_585_p1;
        elsif (((ap_const_logic_1 = ap_CS_fsm_pp0_stage44) and (ap_const_boolean_0 = ap_block_pp0_stage44_01001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op251_write_state46 = ap_const_boolean_1))) then 
            gmem_WDATA <= p_Result_8_fu_554_p1;
        elsif (((ap_const_logic_1 = ap_CS_fsm_pp0_stage43) and (ap_const_boolean_0 = ap_block_pp0_stage43_01001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op248_write_state45 = ap_const_boolean_1))) then 
            gmem_WDATA <= p_Result_13_fu_549_p1;
        elsif (((ap_const_logic_1 = ap_CS_fsm_pp0_stage27) and (ap_const_boolean_0 = ap_block_pp0_stage27_01001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op221_write_state29 = ap_const_boolean_1))) then 
            gmem_WDATA <= p_Result_12_fu_531_p1;
        elsif (((ap_const_logic_1 = ap_CS_fsm_pp0_stage11) and (ap_const_boolean_0 = ap_block_pp0_stage11_01001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op194_write_state13 = ap_const_boolean_1))) then 
            gmem_WDATA <= p_Result_11_fu_515_p1;
        else 
            gmem_WDATA <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
        end if; 
    end process;


    gmem_WSTRB_assign_proc : process(ap_enable_reg_pp0_iter0, ap_enable_reg_pp0_iter1, ap_CS_fsm_pp0_stage9, ap_CS_fsm_pp0_stage44, ap_CS_fsm_pp0_stage60, ap_CS_fsm_pp0_stage76, ap_CS_fsm_pp0_stage11, ap_CS_fsm_pp0_stage27, ap_CS_fsm_pp0_stage43, ap_predicate_op194_write_state13, ap_block_pp0_stage11_01001, ap_predicate_op221_write_state29, ap_block_pp0_stage27_01001, ap_predicate_op248_write_state45, ap_block_pp0_stage43_01001, ap_predicate_op251_write_state46, ap_block_pp0_stage44_01001, ap_predicate_op303_write_state62, ap_block_pp0_stage60_01001, ap_predicate_op330_write_state78, ap_block_pp0_stage76_01001, ap_block_pp0_stage9_01001)
    begin
        if ((((ap_const_logic_1 = ap_CS_fsm_pp0_stage43) and (ap_const_boolean_0 = ap_block_pp0_stage43_01001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op248_write_state45 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage27) and (ap_const_boolean_0 = ap_block_pp0_stage27_01001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op221_write_state29 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage76) and (ap_const_boolean_0 = ap_block_pp0_stage76_01001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op330_write_state78 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage60) and (ap_const_boolean_0 = ap_block_pp0_stage60_01001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op303_write_state62 = ap_const_boolean_1)) or ((ap_enable_reg_pp0_iter1 = ap_const_logic_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage9) and (ap_const_boolean_0 = ap_block_pp0_stage9_01001)))) then 
            gmem_WSTRB <= ap_const_lv16_FFFF;
        elsif ((((ap_const_logic_1 = ap_CS_fsm_pp0_stage11) and (ap_const_boolean_0 = ap_block_pp0_stage11_01001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op194_write_state13 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage44) and (ap_const_boolean_0 = ap_block_pp0_stage44_01001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op251_write_state46 = ap_const_boolean_1)))) then 
            gmem_WSTRB <= ap_const_lv16_F;
        else 
            gmem_WSTRB <= "XXXXXXXXXXXXXXXX";
        end if; 
    end process;


    gmem_WVALID_assign_proc : process(ap_enable_reg_pp0_iter0, ap_enable_reg_pp0_iter1, ap_CS_fsm_pp0_stage9, ap_CS_fsm_pp0_stage44, ap_CS_fsm_pp0_stage60, ap_CS_fsm_pp0_stage76, ap_CS_fsm_pp0_stage11, ap_CS_fsm_pp0_stage27, ap_CS_fsm_pp0_stage43, ap_block_pp0_stage9_11001, ap_predicate_op194_write_state13, ap_block_pp0_stage11_11001, ap_predicate_op221_write_state29, ap_block_pp0_stage27_11001, ap_predicate_op248_write_state45, ap_block_pp0_stage43_11001, ap_predicate_op251_write_state46, ap_block_pp0_stage44_11001, ap_predicate_op303_write_state62, ap_block_pp0_stage60_11001, ap_predicate_op330_write_state78, ap_block_pp0_stage76_11001)
    begin
        if ((((ap_const_logic_1 = ap_CS_fsm_pp0_stage43) and (ap_const_boolean_0 = ap_block_pp0_stage43_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op248_write_state45 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage27) and (ap_const_boolean_0 = ap_block_pp0_stage27_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op221_write_state29 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage11) and (ap_const_boolean_0 = ap_block_pp0_stage11_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op194_write_state13 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage76) and (ap_const_boolean_0 = ap_block_pp0_stage76_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op330_write_state78 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage60) and (ap_const_boolean_0 = ap_block_pp0_stage60_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op303_write_state62 = ap_const_boolean_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage44) and (ap_const_boolean_0 = ap_block_pp0_stage44_11001) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1) and (ap_predicate_op251_write_state46 = ap_const_boolean_1)) or ((ap_enable_reg_pp0_iter1 = ap_const_logic_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage9) and (ap_const_boolean_0 = ap_block_pp0_stage9_11001)))) then 
            gmem_WVALID <= ap_const_logic_1;
        else 
            gmem_WVALID <= ap_const_logic_0;
        end if; 
    end process;


    gmem_blk_n_AR_assign_proc : process(m_axi_gmem_ARREADY, ap_CS_fsm_pp0_stage1, ap_enable_reg_pp0_iter0, ap_block_pp0_stage1, icmp_ln1073_reg_676, ap_CS_fsm_pp0_stage50, ap_block_pp0_stage50, op_read_reg_640, ap_CS_fsm_pp0_stage66, ap_block_pp0_stage66, ap_CS_fsm_pp0_stage82, ap_block_pp0_stage82, ap_enable_reg_pp0_iter1, ap_CS_fsm_pp0_stage17, ap_block_pp0_stage17, ap_CS_fsm_pp0_stage33, ap_block_pp0_stage33, ap_CS_fsm_pp0_stage49, ap_block_pp0_stage49, ap_CS_fsm_pp0_stage2, ap_block_pp0_stage2, ap_CS_fsm_pp0_stage51, ap_block_pp0_stage51, ap_CS_fsm_pp0_stage67, ap_block_pp0_stage67, ap_CS_fsm_pp0_stage0, ap_block_pp0_stage0, ap_CS_fsm_pp0_stage18, ap_block_pp0_stage18, ap_CS_fsm_pp0_stage34, ap_block_pp0_stage34)
    begin
        if ((((ap_const_logic_1 = ap_CS_fsm_pp0_stage2) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage2) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage34) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage34) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage18) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage18) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage49) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage49) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage33) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage33) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage17) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage17) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage50) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage50) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((ap_enable_reg_pp0_iter1 = ap_const_logic_1) and (op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage0) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage0)) or ((op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage67) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage67) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage51) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage51) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage82) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage82) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage66) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage66) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage50) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage50) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage1) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage1) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)))) then 
            gmem_blk_n_AR <= m_axi_gmem_ARREADY;
        else 
            gmem_blk_n_AR <= ap_const_logic_1;
        end if; 
    end process;


    gmem_blk_n_AW_assign_proc : process(m_axi_gmem_AWREADY, ap_CS_fsm_pp0_stage1, ap_enable_reg_pp0_iter0, ap_block_pp0_stage1, icmp_ln1073_reg_676, op_read_reg_640, ap_CS_fsm_pp0_stage2, ap_block_pp0_stage2, ap_CS_fsm_pp0_stage3, ap_block_pp0_stage3, ap_CS_fsm_pp0_stage10, ap_block_pp0_stage10)
    begin
        if ((((ap_const_logic_1 = ap_CS_fsm_pp0_stage10) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage10) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage3) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage3) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage2) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage2) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage1) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage1) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage3) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage3) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage2) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage2) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage1) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage1) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)))) then 
            gmem_blk_n_AW <= m_axi_gmem_AWREADY;
        else 
            gmem_blk_n_AW <= ap_const_logic_1;
        end if; 
    end process;


    gmem_blk_n_B_assign_proc : process(m_axi_gmem_BVALID, ap_enable_reg_pp0_iter0, icmp_ln1073_reg_676, op_read_reg_640, ap_enable_reg_pp0_iter1, ap_CS_fsm_pp0_stage49, ap_block_pp0_stage49, ap_CS_fsm_pp0_stage65, ap_block_pp0_stage65, ap_CS_fsm_pp0_stage81, ap_block_pp0_stage81, ap_CS_fsm_pp0_stage16, ap_block_pp0_stage16, ap_CS_fsm_pp0_stage32, ap_block_pp0_stage32, ap_CS_fsm_pp0_stage48, ap_block_pp0_stage48, ap_CS_fsm_pp0_stage14, ap_block_pp0_stage14)
    begin
        if ((((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage48) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage48) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage32) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage32) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage16) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage16) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((ap_enable_reg_pp0_iter1 = ap_const_logic_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage14) and (ap_const_boolean_0 = ap_block_pp0_stage14)) or ((op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage81) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage81) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage65) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage65) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage49) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage49) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)))) then 
            gmem_blk_n_B <= m_axi_gmem_BVALID;
        else 
            gmem_blk_n_B <= ap_const_logic_1;
        end if; 
    end process;


    gmem_blk_n_R_assign_proc : process(m_axi_gmem_RVALID, ap_enable_reg_pp0_iter0, icmp_ln1073_reg_676, ap_CS_fsm_pp0_stage8, ap_block_pp0_stage8, op_read_reg_640, ap_CS_fsm_pp0_stage57, ap_block_pp0_stage57, ap_CS_fsm_pp0_stage73, ap_block_pp0_stage73, ap_CS_fsm_pp0_stage6, ap_enable_reg_pp0_iter1, ap_block_pp0_stage6, icmp_ln1073_reg_676_pp0_iter1_reg, ap_CS_fsm_pp0_stage24, ap_block_pp0_stage24, ap_CS_fsm_pp0_stage40, ap_block_pp0_stage40, ap_CS_fsm_pp0_stage56, ap_block_pp0_stage56, ap_CS_fsm_pp0_stage9, ap_block_pp0_stage9, ap_CS_fsm_pp0_stage58, ap_block_pp0_stage58, ap_CS_fsm_pp0_stage74, ap_block_pp0_stage74, ap_CS_fsm_pp0_stage7, ap_block_pp0_stage7, ap_CS_fsm_pp0_stage25, ap_block_pp0_stage25, ap_CS_fsm_pp0_stage41, ap_block_pp0_stage41)
    begin
        if ((((ap_const_logic_1 = ap_CS_fsm_pp0_stage9) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage9) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage41) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage41) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage25) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage25) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage56) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage56) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage40) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage40) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage24) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage24) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage57) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage57) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((icmp_ln1073_reg_676_pp0_iter1_reg = ap_const_lv1_1) and (ap_enable_reg_pp0_iter1 = ap_const_logic_1) and (op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage7) and (ap_const_boolean_0 = ap_block_pp0_stage7)) or ((icmp_ln1073_reg_676_pp0_iter1_reg = ap_const_lv1_1) and (ap_enable_reg_pp0_iter1 = ap_const_logic_1) and (op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage6) and (ap_const_boolean_0 = ap_block_pp0_stage6)) or ((op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage74) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage74) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage58) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage58) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage73) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage73) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage57) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage57) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((ap_const_logic_1 = ap_CS_fsm_pp0_stage8) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage8) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)))) then 
            gmem_blk_n_R <= m_axi_gmem_RVALID;
        else 
            gmem_blk_n_R <= ap_const_logic_1;
        end if; 
    end process;


    gmem_blk_n_W_assign_proc : process(m_axi_gmem_WREADY, ap_enable_reg_pp0_iter0, icmp_ln1073_reg_676, op_read_reg_640, ap_enable_reg_pp0_iter1, ap_CS_fsm_pp0_stage9, ap_block_pp0_stage9, ap_CS_fsm_pp0_stage44, ap_block_pp0_stage44, ap_CS_fsm_pp0_stage60, ap_block_pp0_stage60, ap_CS_fsm_pp0_stage76, ap_block_pp0_stage76, ap_CS_fsm_pp0_stage11, ap_block_pp0_stage11, ap_CS_fsm_pp0_stage27, ap_block_pp0_stage27, ap_CS_fsm_pp0_stage43, ap_block_pp0_stage43)
    begin
        if ((((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage43) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage43) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage27) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage27) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage11) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage11) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((ap_enable_reg_pp0_iter1 = ap_const_logic_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage9) and (ap_const_boolean_0 = ap_block_pp0_stage9)) or ((op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage76) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage76) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage60) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage60) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)) or ((op_read_reg_640 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_pp0_stage44) and (icmp_ln1073_reg_676 = ap_const_lv1_1) and (ap_const_boolean_0 = ap_block_pp0_stage44) and (ap_enable_reg_pp0_iter0 = ap_const_logic_1)))) then 
            gmem_blk_n_W <= m_axi_gmem_WREADY;
        else 
            gmem_blk_n_W <= ap_const_logic_1;
        end if; 
    end process;

    i_V_fu_608_p2 <= std_logic_vector(signed(i_V_2_reg_671) + signed(ap_const_lv32_10));
    icmp_ln1073_fu_364_p0 <= rhs_V_fu_122;
    icmp_ln1073_fu_364_p2 <= "1" when (unsigned(icmp_ln1073_fu_364_p0) < unsigned(size_read_reg_644)) else "0";
    lhs_5_fu_348_p1 <= std_logic_vector(IEEE.numeric_std.resize(unsigned(src_addr2),34));
    lhs_6_fu_352_p1 <= std_logic_vector(IEEE.numeric_std.resize(unsigned(dst_addr),34));
    lhs_fu_344_p1 <= std_logic_vector(IEEE.numeric_std.resize(unsigned(src_addr1),34));
    p_Result_10_fu_603_p1 <= std_logic_vector(IEEE.numeric_std.resize(unsigned(tmp_4_fu_596_p4),128));
    p_Result_11_fu_515_p1 <= std_logic_vector(IEEE.numeric_std.resize(unsigned(sub_ln414_reg_731),128));
    p_Result_12_fu_531_p1 <= std_logic_vector(IEEE.numeric_std.resize(unsigned(tmp_9_fu_525_p3),128));
    p_Result_13_fu_549_p1 <= std_logic_vector(IEEE.numeric_std.resize(unsigned(tmp_12_fu_542_p4),128));
    p_Result_4_fu_564_p5 <= (((sub_ln414_3_fu_558_p2 & sub_ln414_2_reg_754) & sub_ln414_1_reg_747) & sub_ln414_reg_731);
    p_Result_8_fu_554_p1 <= std_logic_vector(IEEE.numeric_std.resize(unsigned(add_ln414_1_reg_739),128));
    p_Result_9_fu_585_p1 <= std_logic_vector(IEEE.numeric_std.resize(unsigned(tmp_fu_579_p3),128));
    p_Result_s_fu_624_p5 <= (((add_ln414_4_fu_618_p2 & add_ln414_3_reg_772) & add_ln414_2_reg_765) & add_ln414_1_reg_739);
    ret_V_1_fu_378_p2 <= std_logic_vector(signed(sext_ln232_fu_369_p1) + signed(lhs_5_reg_661));
    ret_V_2_fu_417_p2 <= std_logic_vector(signed(sext_ln232_fu_369_p1) + signed(lhs_6_reg_666));
    ret_V_fu_373_p2 <= std_logic_vector(signed(sext_ln232_fu_369_p1) + signed(lhs_reg_656));
    sext_ln232_fu_369_p0 <= rhs_V_fu_122;
        sext_ln232_fu_369_p1 <= std_logic_vector(IEEE.numeric_std.resize(signed(sext_ln232_fu_369_p0),34));

        sext_ln357_1_fu_489_p1 <= std_logic_vector(IEEE.numeric_std.resize(signed(trunc_ln357_1_reg_685),64));

        sext_ln357_2_fu_391_p1 <= std_logic_vector(IEEE.numeric_std.resize(signed(shl_ln_fu_383_p3),64));

        sext_ln357_3_fu_408_p1 <= std_logic_vector(IEEE.numeric_std.resize(signed(shl_ln357_1_fu_400_p3),64));

        sext_ln357_fu_469_p1 <= std_logic_vector(IEEE.numeric_std.resize(signed(trunc_ln_reg_680),64));

        sext_ln414_1_fu_430_p1 <= std_logic_vector(IEEE.numeric_std.resize(signed(shl_ln1_fu_422_p3),64));

        sext_ln414_fu_479_p1 <= std_logic_vector(IEEE.numeric_std.resize(signed(trunc_ln1_reg_690),64));

    shl_ln1_fu_422_p3 <= (ret_V_2_fu_417_p2 & ap_const_lv4_0);
    shl_ln357_1_fu_400_p3 <= (ret_V_1_fu_378_p2 & ap_const_lv4_0);
    shl_ln_fu_383_p3 <= (ret_V_fu_373_p2 & ap_const_lv4_0);
    sub_ln414_1_fu_519_p2 <= std_logic_vector(unsigned(reg_320) - unsigned(reg_324));
    sub_ln414_2_fu_536_p2 <= std_logic_vector(unsigned(reg_328) - unsigned(reg_332));
    sub_ln414_3_fu_558_p2 <= std_logic_vector(unsigned(reg_336) - unsigned(reg_340));
    sub_ln414_fu_507_p2 <= std_logic_vector(unsigned(trunc_ln357_reg_719) - unsigned(trunc_ln357_2_reg_725));
    tmp_12_fu_542_p4 <= ((sub_ln414_2_reg_754 & sub_ln414_1_reg_747) & sub_ln414_reg_731);
    tmp_4_fu_596_p4 <= ((add_ln414_3_reg_772 & add_ln414_2_reg_765) & add_ln414_1_reg_739);
    tmp_9_fu_525_p3 <= (sub_ln414_1_reg_747 & sub_ln414_reg_731);
    tmp_fu_579_p3 <= (add_ln414_2_reg_765 & add_ln414_1_reg_739);
    trunc_ln357_2_fu_503_p1 <= gmem_RDATA(32 - 1 downto 0);
    trunc_ln357_fu_499_p1 <= gmem_RDATA(32 - 1 downto 0);
end behav;
