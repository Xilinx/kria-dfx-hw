-- Copyright (C) 2022, Advanced Micro Devices, Inc. All rights reserved.
-- SPDX-License-Identifier: MIT
-- ==============================================================
-- Version: 2022.1
-- 
-- ===========================================================

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity pp_pipeline_accel_Axi2AxiStream is
port (
    ap_clk : IN STD_LOGIC;
    ap_rst : IN STD_LOGIC;
    ap_start : IN STD_LOGIC;
    ap_done : OUT STD_LOGIC;
    ap_continue : IN STD_LOGIC;
    ap_idle : OUT STD_LOGIC;
    ap_ready : OUT STD_LOGIC;
    m_axi_gmem2_AWVALID : OUT STD_LOGIC;
    m_axi_gmem2_AWREADY : IN STD_LOGIC;
    m_axi_gmem2_AWADDR : OUT STD_LOGIC_VECTOR (63 downto 0);
    m_axi_gmem2_AWID : OUT STD_LOGIC_VECTOR (0 downto 0);
    m_axi_gmem2_AWLEN : OUT STD_LOGIC_VECTOR (31 downto 0);
    m_axi_gmem2_AWSIZE : OUT STD_LOGIC_VECTOR (2 downto 0);
    m_axi_gmem2_AWBURST : OUT STD_LOGIC_VECTOR (1 downto 0);
    m_axi_gmem2_AWLOCK : OUT STD_LOGIC_VECTOR (1 downto 0);
    m_axi_gmem2_AWCACHE : OUT STD_LOGIC_VECTOR (3 downto 0);
    m_axi_gmem2_AWPROT : OUT STD_LOGIC_VECTOR (2 downto 0);
    m_axi_gmem2_AWQOS : OUT STD_LOGIC_VECTOR (3 downto 0);
    m_axi_gmem2_AWREGION : OUT STD_LOGIC_VECTOR (3 downto 0);
    m_axi_gmem2_AWUSER : OUT STD_LOGIC_VECTOR (0 downto 0);
    m_axi_gmem2_WVALID : OUT STD_LOGIC;
    m_axi_gmem2_WREADY : IN STD_LOGIC;
    m_axi_gmem2_WDATA : OUT STD_LOGIC_VECTOR (63 downto 0);
    m_axi_gmem2_WSTRB : OUT STD_LOGIC_VECTOR (7 downto 0);
    m_axi_gmem2_WLAST : OUT STD_LOGIC;
    m_axi_gmem2_WID : OUT STD_LOGIC_VECTOR (0 downto 0);
    m_axi_gmem2_WUSER : OUT STD_LOGIC_VECTOR (0 downto 0);
    m_axi_gmem2_ARVALID : OUT STD_LOGIC;
    m_axi_gmem2_ARREADY : IN STD_LOGIC;
    m_axi_gmem2_ARADDR : OUT STD_LOGIC_VECTOR (63 downto 0);
    m_axi_gmem2_ARID : OUT STD_LOGIC_VECTOR (0 downto 0);
    m_axi_gmem2_ARLEN : OUT STD_LOGIC_VECTOR (31 downto 0);
    m_axi_gmem2_ARSIZE : OUT STD_LOGIC_VECTOR (2 downto 0);
    m_axi_gmem2_ARBURST : OUT STD_LOGIC_VECTOR (1 downto 0);
    m_axi_gmem2_ARLOCK : OUT STD_LOGIC_VECTOR (1 downto 0);
    m_axi_gmem2_ARCACHE : OUT STD_LOGIC_VECTOR (3 downto 0);
    m_axi_gmem2_ARPROT : OUT STD_LOGIC_VECTOR (2 downto 0);
    m_axi_gmem2_ARQOS : OUT STD_LOGIC_VECTOR (3 downto 0);
    m_axi_gmem2_ARREGION : OUT STD_LOGIC_VECTOR (3 downto 0);
    m_axi_gmem2_ARUSER : OUT STD_LOGIC_VECTOR (0 downto 0);
    m_axi_gmem2_RVALID : IN STD_LOGIC;
    m_axi_gmem2_RREADY : OUT STD_LOGIC;
    m_axi_gmem2_RDATA : IN STD_LOGIC_VECTOR (63 downto 0);
    m_axi_gmem2_RLAST : IN STD_LOGIC;
    m_axi_gmem2_RID : IN STD_LOGIC_VECTOR (0 downto 0);
    m_axi_gmem2_RFIFONUM : IN STD_LOGIC_VECTOR (8 downto 0);
    m_axi_gmem2_RUSER : IN STD_LOGIC_VECTOR (0 downto 0);
    m_axi_gmem2_RRESP : IN STD_LOGIC_VECTOR (1 downto 0);
    m_axi_gmem2_BVALID : IN STD_LOGIC;
    m_axi_gmem2_BREADY : OUT STD_LOGIC;
    m_axi_gmem2_BRESP : IN STD_LOGIC_VECTOR (1 downto 0);
    m_axi_gmem2_BID : IN STD_LOGIC_VECTOR (0 downto 0);
    m_axi_gmem2_BUSER : IN STD_LOGIC_VECTOR (0 downto 0);
    din : IN STD_LOGIC_VECTOR (63 downto 0);
    ldata_din : OUT STD_LOGIC_VECTOR (63 downto 0);
    ldata_num_data_valid : IN STD_LOGIC_VECTOR (1 downto 0);
    ldata_fifo_cap : IN STD_LOGIC_VECTOR (1 downto 0);
    ldata_full_n : IN STD_LOGIC;
    ldata_write : OUT STD_LOGIC;
    p_read : IN STD_LOGIC_VECTOR (10 downto 0);
    p_read1 : IN STD_LOGIC_VECTOR (10 downto 0);
    cols : IN STD_LOGIC_VECTOR (10 downto 0);
    stride : IN STD_LOGIC_VECTOR (31 downto 0);
    cols_c_din : OUT STD_LOGIC_VECTOR (10 downto 0);
    cols_c_num_data_valid : IN STD_LOGIC_VECTOR (1 downto 0);
    cols_c_fifo_cap : IN STD_LOGIC_VECTOR (1 downto 0);
    cols_c_full_n : IN STD_LOGIC;
    cols_c_write : OUT STD_LOGIC );
end;


architecture behav of pp_pipeline_accel_Axi2AxiStream is 
    constant ap_const_logic_1 : STD_LOGIC := '1';
    constant ap_const_logic_0 : STD_LOGIC := '0';
    constant ap_ST_fsm_state1 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000001";
    constant ap_ST_fsm_state2 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000010";
    constant ap_ST_fsm_state3 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000100";
    constant ap_ST_fsm_state4 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000001000";
    constant ap_ST_fsm_state5 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000010000";
    constant ap_ST_fsm_state6 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000100000";
    constant ap_ST_fsm_state7 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000001000000";
    constant ap_ST_fsm_state8 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000010000000";
    constant ap_ST_fsm_state9 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000100000000";
    constant ap_ST_fsm_state10 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000001000000000";
    constant ap_ST_fsm_state11 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000010000000000";
    constant ap_ST_fsm_state12 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000100000000000";
    constant ap_ST_fsm_state13 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000001000000000000";
    constant ap_ST_fsm_state14 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000010000000000000";
    constant ap_ST_fsm_state15 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000100000000000000";
    constant ap_ST_fsm_state16 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000000000000000001000000000000000";
    constant ap_ST_fsm_state17 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000000000000000010000000000000000";
    constant ap_ST_fsm_state18 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000000000000000100000000000000000";
    constant ap_ST_fsm_state19 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000000000000001000000000000000000";
    constant ap_ST_fsm_state20 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000000000000010000000000000000000";
    constant ap_ST_fsm_state21 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000000000000100000000000000000000";
    constant ap_ST_fsm_state22 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000000000001000000000000000000000";
    constant ap_ST_fsm_state23 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000000000010000000000000000000000";
    constant ap_ST_fsm_state24 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000000000100000000000000000000000";
    constant ap_ST_fsm_state25 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000000001000000000000000000000000";
    constant ap_ST_fsm_state26 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000000010000000000000000000000000";
    constant ap_ST_fsm_state27 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000000100000000000000000000000000";
    constant ap_ST_fsm_state28 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000001000000000000000000000000000";
    constant ap_ST_fsm_state29 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000010000000000000000000000000000";
    constant ap_ST_fsm_state30 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000100000000000000000000000000000";
    constant ap_ST_fsm_state31 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000001000000000000000000000000000000";
    constant ap_ST_fsm_state32 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000010000000000000000000000000000000";
    constant ap_ST_fsm_state33 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000100000000000000000000000000000000";
    constant ap_ST_fsm_state34 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000001000000000000000000000000000000000";
    constant ap_ST_fsm_state35 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000010000000000000000000000000000000000";
    constant ap_ST_fsm_state36 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000100000000000000000000000000000000000";
    constant ap_ST_fsm_state37 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000001000000000000000000000000000000000000";
    constant ap_ST_fsm_state38 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000010000000000000000000000000000000000000";
    constant ap_ST_fsm_state39 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000100000000000000000000000000000000000000";
    constant ap_ST_fsm_state40 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000001000000000000000000000000000000000000000";
    constant ap_ST_fsm_state41 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000010000000000000000000000000000000000000000";
    constant ap_ST_fsm_state42 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000100000000000000000000000000000000000000000";
    constant ap_ST_fsm_state43 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000001000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state44 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000010000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state45 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000100000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state46 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000001000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state47 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000010000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state48 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000100000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state49 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000001000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state50 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000010000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state51 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000100000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state52 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000001000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state53 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000010000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state54 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000100000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state55 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000001000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state56 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000010000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state57 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000100000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state58 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000001000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state59 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000010000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state60 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000100000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state61 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000001000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state62 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000010000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state63 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000100000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state64 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000001000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state65 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000010000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state66 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000100000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state67 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000001000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state68 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000010000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state69 : STD_LOGIC_VECTOR (80 downto 0) := "000000000000100000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state70 : STD_LOGIC_VECTOR (80 downto 0) := "000000000001000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state71 : STD_LOGIC_VECTOR (80 downto 0) := "000000000010000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state72 : STD_LOGIC_VECTOR (80 downto 0) := "000000000100000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state73 : STD_LOGIC_VECTOR (80 downto 0) := "000000001000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state74 : STD_LOGIC_VECTOR (80 downto 0) := "000000010000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state75 : STD_LOGIC_VECTOR (80 downto 0) := "000000100000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state76 : STD_LOGIC_VECTOR (80 downto 0) := "000001000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state77 : STD_LOGIC_VECTOR (80 downto 0) := "000010000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state78 : STD_LOGIC_VECTOR (80 downto 0) := "000100000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state79 : STD_LOGIC_VECTOR (80 downto 0) := "001000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state80 : STD_LOGIC_VECTOR (80 downto 0) := "010000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_ST_fsm_state81 : STD_LOGIC_VECTOR (80 downto 0) := "100000000000000000000000000000000000000000000000000000000000000000000000000000000";
    constant ap_const_lv32_0 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000000";
    constant ap_const_boolean_1 : BOOLEAN := true;
    constant ap_const_lv64_0 : STD_LOGIC_VECTOR (63 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000";
    constant ap_const_lv1_0 : STD_LOGIC_VECTOR (0 downto 0) := "0";
    constant ap_const_lv3_0 : STD_LOGIC_VECTOR (2 downto 0) := "000";
    constant ap_const_lv2_0 : STD_LOGIC_VECTOR (1 downto 0) := "00";
    constant ap_const_lv4_0 : STD_LOGIC_VECTOR (3 downto 0) := "0000";
    constant ap_const_lv8_0 : STD_LOGIC_VECTOR (7 downto 0) := "00000000";
    constant ap_const_lv32_9 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000001001";
    constant ap_const_lv32_1 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000001";
    constant ap_const_lv32_3 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000011";
    constant ap_const_lv32_4 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000100";
    constant ap_const_lv32_5 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000101";
    constant ap_const_lv32_8 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000001000";
    constant ap_const_lv32_4F : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000001001111";
    constant ap_const_lv32_50 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000001010000";
    constant ap_const_lv11_0 : STD_LOGIC_VECTOR (10 downto 0) := "00000000000";
    constant ap_const_boolean_0 : BOOLEAN := false;
    constant ap_const_lv32_FFFFFFFF : STD_LOGIC_VECTOR (31 downto 0) := "11111111111111111111111111111111";
    constant ap_const_lv26_3F : STD_LOGIC_VECTOR (25 downto 0) := "00000000000000000000111111";
    constant ap_const_lv32_6 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000000110";
    constant ap_const_lv32_19 : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000011001";
    constant ap_const_lv20_0 : STD_LOGIC_VECTOR (19 downto 0) := "00000000000000000000";
    constant ap_const_lv11_1 : STD_LOGIC_VECTOR (10 downto 0) := "00000000001";
    constant ap_const_lv32_3F : STD_LOGIC_VECTOR (31 downto 0) := "00000000000000000000000000111111";
    constant ap_const_lv1_1 : STD_LOGIC_VECTOR (0 downto 0) := "1";

attribute shreg_extract : string;
    signal ap_done_reg : STD_LOGIC := '0';
    signal ap_CS_fsm : STD_LOGIC_VECTOR (80 downto 0) := "000000000000000000000000000000000000000000000000000000000000000000000000000000001";
    attribute fsm_encoding : string;
    attribute fsm_encoding of ap_CS_fsm : signal is "none";
    signal ap_CS_fsm_state1 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_state1 : signal is "none";
    signal gmem2_blk_n_AR : STD_LOGIC;
    signal ap_CS_fsm_state10 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_state10 : signal is "none";
    signal cols_c_blk_n : STD_LOGIC;
    signal cols_int16_fu_174_p1 : STD_LOGIC_VECTOR (15 downto 0);
    signal cols_int16_reg_366 : STD_LOGIC_VECTOR (15 downto 0);
    signal icmp_ln1021_fu_178_p2 : STD_LOGIC_VECTOR (0 downto 0);
    signal icmp_ln1021_reg_371 : STD_LOGIC_VECTOR (0 downto 0);
    signal ap_CS_fsm_state2 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_state2 : signal is "none";
    signal grp_fu_329_p2 : STD_LOGIC_VECTOR (21 downto 0);
    signal ret_V_36_reg_396 : STD_LOGIC_VECTOR (21 downto 0);
    signal ap_CS_fsm_state4 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_state4 : signal is "none";
    signal trunc_ln1540_fu_201_p1 : STD_LOGIC_VECTOR (21 downto 0);
    signal trunc_ln1540_reg_401 : STD_LOGIC_VECTOR (21 downto 0);
    signal ap_CS_fsm_state5 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_state5 : signal is "none";
    signal cols_addrbound_fu_217_p4 : STD_LOGIC_VECTOR (19 downto 0);
    signal cols_addrbound_reg_416 : STD_LOGIC_VECTOR (19 downto 0);
    signal cmp_i82_i_fu_257_p2 : STD_LOGIC_VECTOR (0 downto 0);
    signal cmp_i82_i_reg_421 : STD_LOGIC_VECTOR (0 downto 0);
    signal zext_ln1028_fu_263_p1 : STD_LOGIC_VECTOR (30 downto 0);
    signal zext_ln1028_reg_425 : STD_LOGIC_VECTOR (30 downto 0);
    signal zext_ln1028_1_fu_267_p1 : STD_LOGIC_VECTOR (31 downto 0);
    signal zext_ln1028_1_reg_430 : STD_LOGIC_VECTOR (31 downto 0);
    signal r_4_fu_279_p2 : STD_LOGIC_VECTOR (10 downto 0);
    signal r_4_reg_438 : STD_LOGIC_VECTOR (10 downto 0);
    signal ap_CS_fsm_state6 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_state6 : signal is "none";
    signal icmp_ln1024_fu_274_p2 : STD_LOGIC_VECTOR (0 downto 0);
    signal trunc_ln_reg_448 : STD_LOGIC_VECTOR (60 downto 0);
    signal ap_CS_fsm_state9 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_state9 : signal is "none";
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_ap_start : STD_LOGIC;
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_ap_done : STD_LOGIC;
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_ap_idle : STD_LOGIC;
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_ap_ready : STD_LOGIC;
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_AWVALID : STD_LOGIC;
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_AWADDR : STD_LOGIC_VECTOR (63 downto 0);
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_AWID : STD_LOGIC_VECTOR (0 downto 0);
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_AWLEN : STD_LOGIC_VECTOR (31 downto 0);
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_AWSIZE : STD_LOGIC_VECTOR (2 downto 0);
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_AWBURST : STD_LOGIC_VECTOR (1 downto 0);
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_AWLOCK : STD_LOGIC_VECTOR (1 downto 0);
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_AWCACHE : STD_LOGIC_VECTOR (3 downto 0);
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_AWPROT : STD_LOGIC_VECTOR (2 downto 0);
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_AWQOS : STD_LOGIC_VECTOR (3 downto 0);
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_AWREGION : STD_LOGIC_VECTOR (3 downto 0);
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_AWUSER : STD_LOGIC_VECTOR (0 downto 0);
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_WVALID : STD_LOGIC;
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_WDATA : STD_LOGIC_VECTOR (63 downto 0);
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_WSTRB : STD_LOGIC_VECTOR (7 downto 0);
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_WLAST : STD_LOGIC;
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_WID : STD_LOGIC_VECTOR (0 downto 0);
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_WUSER : STD_LOGIC_VECTOR (0 downto 0);
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARVALID : STD_LOGIC;
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARADDR : STD_LOGIC_VECTOR (63 downto 0);
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARID : STD_LOGIC_VECTOR (0 downto 0);
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARLEN : STD_LOGIC_VECTOR (31 downto 0);
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARSIZE : STD_LOGIC_VECTOR (2 downto 0);
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARBURST : STD_LOGIC_VECTOR (1 downto 0);
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARLOCK : STD_LOGIC_VECTOR (1 downto 0);
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARCACHE : STD_LOGIC_VECTOR (3 downto 0);
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARPROT : STD_LOGIC_VECTOR (2 downto 0);
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARQOS : STD_LOGIC_VECTOR (3 downto 0);
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARREGION : STD_LOGIC_VECTOR (3 downto 0);
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARUSER : STD_LOGIC_VECTOR (0 downto 0);
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_RREADY : STD_LOGIC;
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_BREADY : STD_LOGIC;
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_ldata_din : STD_LOGIC_VECTOR (63 downto 0);
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_ldata_write : STD_LOGIC;
    signal grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_ap_start_reg : STD_LOGIC := '0';
    signal ap_CS_fsm_state80 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_state80 : signal is "none";
    signal ap_CS_fsm_state81 : STD_LOGIC;
    attribute fsm_encoding of ap_CS_fsm_state81 : signal is "none";
    signal sext_ln1028_fu_315_p1 : STD_LOGIC_VECTOR (63 downto 0);
    signal r_fu_116 : STD_LOGIC_VECTOR (10 downto 0);
    signal ap_block_state81_on_subcall_done : BOOLEAN;
    signal ap_block_state1 : BOOLEAN;
    signal trunc_ln1540_fu_201_p0 : STD_LOGIC_VECTOR (26 downto 0);
    signal grp_fu_335_p2 : STD_LOGIC_VECTOR (26 downto 0);
    signal ret_V_fu_204_p3 : STD_LOGIC_VECTOR (25 downto 0);
    signal add_ln587_fu_211_p2 : STD_LOGIC_VECTOR (25 downto 0);
    signal ret_V_7_fu_227_p3 : STD_LOGIC_VECTOR (25 downto 0);
    signal add_ln587_1_fu_234_p2 : STD_LOGIC_VECTOR (25 downto 0);
    signal stride_addrbound_fu_240_p4 : STD_LOGIC_VECTOR (19 downto 0);
    signal addrbound_V_fu_250_p3 : STD_LOGIC_VECTOR (19 downto 0);
    signal tmp_s_fu_289_p1 : STD_LOGIC_VECTOR (30 downto 0);
    signal grp_fu_342_p2 : STD_LOGIC_VECTOR (30 downto 0);
    signal tmp_s_fu_289_p3 : STD_LOGIC_VECTOR (33 downto 0);
    signal p_cast2_i_fu_296_p1 : STD_LOGIC_VECTOR (63 downto 0);
    signal empty_229_fu_300_p2 : STD_LOGIC_VECTOR (63 downto 0);
    signal grp_fu_329_p0 : STD_LOGIC_VECTOR (10 downto 0);
    signal grp_fu_329_p1 : STD_LOGIC_VECTOR (10 downto 0);
    signal grp_fu_335_p0 : STD_LOGIC_VECTOR (15 downto 0);
    signal grp_fu_335_p1 : STD_LOGIC_VECTOR (10 downto 0);
    signal grp_fu_342_p0 : STD_LOGIC_VECTOR (19 downto 0);
    signal grp_fu_342_p1 : STD_LOGIC_VECTOR (10 downto 0);
    signal ap_NS_fsm : STD_LOGIC_VECTOR (80 downto 0);
    signal ap_ST_fsm_state1_blk : STD_LOGIC;
    signal ap_ST_fsm_state2_blk : STD_LOGIC;
    signal ap_ST_fsm_state3_blk : STD_LOGIC;
    signal ap_ST_fsm_state4_blk : STD_LOGIC;
    signal ap_ST_fsm_state5_blk : STD_LOGIC;
    signal ap_ST_fsm_state6_blk : STD_LOGIC;
    signal ap_ST_fsm_state7_blk : STD_LOGIC;
    signal ap_ST_fsm_state8_blk : STD_LOGIC;
    signal ap_ST_fsm_state9_blk : STD_LOGIC;
    signal ap_ST_fsm_state10_blk : STD_LOGIC;
    signal ap_ST_fsm_state11_blk : STD_LOGIC;
    signal ap_ST_fsm_state12_blk : STD_LOGIC;
    signal ap_ST_fsm_state13_blk : STD_LOGIC;
    signal ap_ST_fsm_state14_blk : STD_LOGIC;
    signal ap_ST_fsm_state15_blk : STD_LOGIC;
    signal ap_ST_fsm_state16_blk : STD_LOGIC;
    signal ap_ST_fsm_state17_blk : STD_LOGIC;
    signal ap_ST_fsm_state18_blk : STD_LOGIC;
    signal ap_ST_fsm_state19_blk : STD_LOGIC;
    signal ap_ST_fsm_state20_blk : STD_LOGIC;
    signal ap_ST_fsm_state21_blk : STD_LOGIC;
    signal ap_ST_fsm_state22_blk : STD_LOGIC;
    signal ap_ST_fsm_state23_blk : STD_LOGIC;
    signal ap_ST_fsm_state24_blk : STD_LOGIC;
    signal ap_ST_fsm_state25_blk : STD_LOGIC;
    signal ap_ST_fsm_state26_blk : STD_LOGIC;
    signal ap_ST_fsm_state27_blk : STD_LOGIC;
    signal ap_ST_fsm_state28_blk : STD_LOGIC;
    signal ap_ST_fsm_state29_blk : STD_LOGIC;
    signal ap_ST_fsm_state30_blk : STD_LOGIC;
    signal ap_ST_fsm_state31_blk : STD_LOGIC;
    signal ap_ST_fsm_state32_blk : STD_LOGIC;
    signal ap_ST_fsm_state33_blk : STD_LOGIC;
    signal ap_ST_fsm_state34_blk : STD_LOGIC;
    signal ap_ST_fsm_state35_blk : STD_LOGIC;
    signal ap_ST_fsm_state36_blk : STD_LOGIC;
    signal ap_ST_fsm_state37_blk : STD_LOGIC;
    signal ap_ST_fsm_state38_blk : STD_LOGIC;
    signal ap_ST_fsm_state39_blk : STD_LOGIC;
    signal ap_ST_fsm_state40_blk : STD_LOGIC;
    signal ap_ST_fsm_state41_blk : STD_LOGIC;
    signal ap_ST_fsm_state42_blk : STD_LOGIC;
    signal ap_ST_fsm_state43_blk : STD_LOGIC;
    signal ap_ST_fsm_state44_blk : STD_LOGIC;
    signal ap_ST_fsm_state45_blk : STD_LOGIC;
    signal ap_ST_fsm_state46_blk : STD_LOGIC;
    signal ap_ST_fsm_state47_blk : STD_LOGIC;
    signal ap_ST_fsm_state48_blk : STD_LOGIC;
    signal ap_ST_fsm_state49_blk : STD_LOGIC;
    signal ap_ST_fsm_state50_blk : STD_LOGIC;
    signal ap_ST_fsm_state51_blk : STD_LOGIC;
    signal ap_ST_fsm_state52_blk : STD_LOGIC;
    signal ap_ST_fsm_state53_blk : STD_LOGIC;
    signal ap_ST_fsm_state54_blk : STD_LOGIC;
    signal ap_ST_fsm_state55_blk : STD_LOGIC;
    signal ap_ST_fsm_state56_blk : STD_LOGIC;
    signal ap_ST_fsm_state57_blk : STD_LOGIC;
    signal ap_ST_fsm_state58_blk : STD_LOGIC;
    signal ap_ST_fsm_state59_blk : STD_LOGIC;
    signal ap_ST_fsm_state60_blk : STD_LOGIC;
    signal ap_ST_fsm_state61_blk : STD_LOGIC;
    signal ap_ST_fsm_state62_blk : STD_LOGIC;
    signal ap_ST_fsm_state63_blk : STD_LOGIC;
    signal ap_ST_fsm_state64_blk : STD_LOGIC;
    signal ap_ST_fsm_state65_blk : STD_LOGIC;
    signal ap_ST_fsm_state66_blk : STD_LOGIC;
    signal ap_ST_fsm_state67_blk : STD_LOGIC;
    signal ap_ST_fsm_state68_blk : STD_LOGIC;
    signal ap_ST_fsm_state69_blk : STD_LOGIC;
    signal ap_ST_fsm_state70_blk : STD_LOGIC;
    signal ap_ST_fsm_state71_blk : STD_LOGIC;
    signal ap_ST_fsm_state72_blk : STD_LOGIC;
    signal ap_ST_fsm_state73_blk : STD_LOGIC;
    signal ap_ST_fsm_state74_blk : STD_LOGIC;
    signal ap_ST_fsm_state75_blk : STD_LOGIC;
    signal ap_ST_fsm_state76_blk : STD_LOGIC;
    signal ap_ST_fsm_state77_blk : STD_LOGIC;
    signal ap_ST_fsm_state78_blk : STD_LOGIC;
    signal ap_ST_fsm_state79_blk : STD_LOGIC;
    signal ap_ST_fsm_state80_blk : STD_LOGIC;
    signal ap_ST_fsm_state81_blk : STD_LOGIC;
    signal grp_fu_329_p00 : STD_LOGIC_VECTOR (21 downto 0);
    signal grp_fu_329_p10 : STD_LOGIC_VECTOR (21 downto 0);
    signal grp_fu_335_p00 : STD_LOGIC_VECTOR (26 downto 0);
    signal grp_fu_335_p10 : STD_LOGIC_VECTOR (26 downto 0);
    signal grp_fu_342_p10 : STD_LOGIC_VECTOR (30 downto 0);
    signal ap_ce_reg : STD_LOGIC;

    component pp_pipeline_accel_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1 IS
    port (
        ap_clk : IN STD_LOGIC;
        ap_rst : IN STD_LOGIC;
        ap_start : IN STD_LOGIC;
        ap_done : OUT STD_LOGIC;
        ap_idle : OUT STD_LOGIC;
        ap_ready : OUT STD_LOGIC;
        m_axi_gmem2_AWVALID : OUT STD_LOGIC;
        m_axi_gmem2_AWREADY : IN STD_LOGIC;
        m_axi_gmem2_AWADDR : OUT STD_LOGIC_VECTOR (63 downto 0);
        m_axi_gmem2_AWID : OUT STD_LOGIC_VECTOR (0 downto 0);
        m_axi_gmem2_AWLEN : OUT STD_LOGIC_VECTOR (31 downto 0);
        m_axi_gmem2_AWSIZE : OUT STD_LOGIC_VECTOR (2 downto 0);
        m_axi_gmem2_AWBURST : OUT STD_LOGIC_VECTOR (1 downto 0);
        m_axi_gmem2_AWLOCK : OUT STD_LOGIC_VECTOR (1 downto 0);
        m_axi_gmem2_AWCACHE : OUT STD_LOGIC_VECTOR (3 downto 0);
        m_axi_gmem2_AWPROT : OUT STD_LOGIC_VECTOR (2 downto 0);
        m_axi_gmem2_AWQOS : OUT STD_LOGIC_VECTOR (3 downto 0);
        m_axi_gmem2_AWREGION : OUT STD_LOGIC_VECTOR (3 downto 0);
        m_axi_gmem2_AWUSER : OUT STD_LOGIC_VECTOR (0 downto 0);
        m_axi_gmem2_WVALID : OUT STD_LOGIC;
        m_axi_gmem2_WREADY : IN STD_LOGIC;
        m_axi_gmem2_WDATA : OUT STD_LOGIC_VECTOR (63 downto 0);
        m_axi_gmem2_WSTRB : OUT STD_LOGIC_VECTOR (7 downto 0);
        m_axi_gmem2_WLAST : OUT STD_LOGIC;
        m_axi_gmem2_WID : OUT STD_LOGIC_VECTOR (0 downto 0);
        m_axi_gmem2_WUSER : OUT STD_LOGIC_VECTOR (0 downto 0);
        m_axi_gmem2_ARVALID : OUT STD_LOGIC;
        m_axi_gmem2_ARREADY : IN STD_LOGIC;
        m_axi_gmem2_ARADDR : OUT STD_LOGIC_VECTOR (63 downto 0);
        m_axi_gmem2_ARID : OUT STD_LOGIC_VECTOR (0 downto 0);
        m_axi_gmem2_ARLEN : OUT STD_LOGIC_VECTOR (31 downto 0);
        m_axi_gmem2_ARSIZE : OUT STD_LOGIC_VECTOR (2 downto 0);
        m_axi_gmem2_ARBURST : OUT STD_LOGIC_VECTOR (1 downto 0);
        m_axi_gmem2_ARLOCK : OUT STD_LOGIC_VECTOR (1 downto 0);
        m_axi_gmem2_ARCACHE : OUT STD_LOGIC_VECTOR (3 downto 0);
        m_axi_gmem2_ARPROT : OUT STD_LOGIC_VECTOR (2 downto 0);
        m_axi_gmem2_ARQOS : OUT STD_LOGIC_VECTOR (3 downto 0);
        m_axi_gmem2_ARREGION : OUT STD_LOGIC_VECTOR (3 downto 0);
        m_axi_gmem2_ARUSER : OUT STD_LOGIC_VECTOR (0 downto 0);
        m_axi_gmem2_RVALID : IN STD_LOGIC;
        m_axi_gmem2_RREADY : OUT STD_LOGIC;
        m_axi_gmem2_RDATA : IN STD_LOGIC_VECTOR (63 downto 0);
        m_axi_gmem2_RLAST : IN STD_LOGIC;
        m_axi_gmem2_RID : IN STD_LOGIC_VECTOR (0 downto 0);
        m_axi_gmem2_RFIFONUM : IN STD_LOGIC_VECTOR (8 downto 0);
        m_axi_gmem2_RUSER : IN STD_LOGIC_VECTOR (0 downto 0);
        m_axi_gmem2_RRESP : IN STD_LOGIC_VECTOR (1 downto 0);
        m_axi_gmem2_BVALID : IN STD_LOGIC;
        m_axi_gmem2_BREADY : OUT STD_LOGIC;
        m_axi_gmem2_BRESP : IN STD_LOGIC_VECTOR (1 downto 0);
        m_axi_gmem2_BID : IN STD_LOGIC_VECTOR (0 downto 0);
        m_axi_gmem2_BUSER : IN STD_LOGIC_VECTOR (0 downto 0);
        ldata_din : OUT STD_LOGIC_VECTOR (63 downto 0);
        ldata_num_data_valid : IN STD_LOGIC_VECTOR (1 downto 0);
        ldata_fifo_cap : IN STD_LOGIC_VECTOR (1 downto 0);
        ldata_full_n : IN STD_LOGIC;
        ldata_write : OUT STD_LOGIC;
        sext_ln1028 : IN STD_LOGIC_VECTOR (60 downto 0);
        cols_addrbound : IN STD_LOGIC_VECTOR (19 downto 0) );
    end component;


    component pp_pipeline_accel_mul_mul_11ns_11ns_22_3_1 IS
    generic (
        ID : INTEGER;
        NUM_STAGE : INTEGER;
        din0_WIDTH : INTEGER;
        din1_WIDTH : INTEGER;
        dout_WIDTH : INTEGER );
    port (
        clk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        din0 : IN STD_LOGIC_VECTOR (10 downto 0);
        din1 : IN STD_LOGIC_VECTOR (10 downto 0);
        ce : IN STD_LOGIC;
        dout : OUT STD_LOGIC_VECTOR (21 downto 0) );
    end component;


    component pp_pipeline_accel_mul_mul_16ns_11ns_27_3_1 IS
    generic (
        ID : INTEGER;
        NUM_STAGE : INTEGER;
        din0_WIDTH : INTEGER;
        din1_WIDTH : INTEGER;
        dout_WIDTH : INTEGER );
    port (
        clk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        din0 : IN STD_LOGIC_VECTOR (15 downto 0);
        din1 : IN STD_LOGIC_VECTOR (10 downto 0);
        ce : IN STD_LOGIC;
        dout : OUT STD_LOGIC_VECTOR (26 downto 0) );
    end component;


    component pp_pipeline_accel_mul_mul_20ns_11ns_31_4_1 IS
    generic (
        ID : INTEGER;
        NUM_STAGE : INTEGER;
        din0_WIDTH : INTEGER;
        din1_WIDTH : INTEGER;
        dout_WIDTH : INTEGER );
    port (
        clk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        din0 : IN STD_LOGIC_VECTOR (19 downto 0);
        din1 : IN STD_LOGIC_VECTOR (10 downto 0);
        ce : IN STD_LOGIC;
        dout : OUT STD_LOGIC_VECTOR (30 downto 0) );
    end component;



begin
    grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164 : component pp_pipeline_accel_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1
    port map (
        ap_clk => ap_clk,
        ap_rst => ap_rst,
        ap_start => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_ap_start,
        ap_done => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_ap_done,
        ap_idle => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_ap_idle,
        ap_ready => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_ap_ready,
        m_axi_gmem2_AWVALID => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_AWVALID,
        m_axi_gmem2_AWREADY => ap_const_logic_0,
        m_axi_gmem2_AWADDR => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_AWADDR,
        m_axi_gmem2_AWID => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_AWID,
        m_axi_gmem2_AWLEN => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_AWLEN,
        m_axi_gmem2_AWSIZE => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_AWSIZE,
        m_axi_gmem2_AWBURST => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_AWBURST,
        m_axi_gmem2_AWLOCK => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_AWLOCK,
        m_axi_gmem2_AWCACHE => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_AWCACHE,
        m_axi_gmem2_AWPROT => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_AWPROT,
        m_axi_gmem2_AWQOS => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_AWQOS,
        m_axi_gmem2_AWREGION => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_AWREGION,
        m_axi_gmem2_AWUSER => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_AWUSER,
        m_axi_gmem2_WVALID => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_WVALID,
        m_axi_gmem2_WREADY => ap_const_logic_0,
        m_axi_gmem2_WDATA => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_WDATA,
        m_axi_gmem2_WSTRB => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_WSTRB,
        m_axi_gmem2_WLAST => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_WLAST,
        m_axi_gmem2_WID => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_WID,
        m_axi_gmem2_WUSER => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_WUSER,
        m_axi_gmem2_ARVALID => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARVALID,
        m_axi_gmem2_ARREADY => m_axi_gmem2_ARREADY,
        m_axi_gmem2_ARADDR => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARADDR,
        m_axi_gmem2_ARID => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARID,
        m_axi_gmem2_ARLEN => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARLEN,
        m_axi_gmem2_ARSIZE => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARSIZE,
        m_axi_gmem2_ARBURST => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARBURST,
        m_axi_gmem2_ARLOCK => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARLOCK,
        m_axi_gmem2_ARCACHE => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARCACHE,
        m_axi_gmem2_ARPROT => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARPROT,
        m_axi_gmem2_ARQOS => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARQOS,
        m_axi_gmem2_ARREGION => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARREGION,
        m_axi_gmem2_ARUSER => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARUSER,
        m_axi_gmem2_RVALID => m_axi_gmem2_RVALID,
        m_axi_gmem2_RREADY => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_RREADY,
        m_axi_gmem2_RDATA => m_axi_gmem2_RDATA,
        m_axi_gmem2_RLAST => m_axi_gmem2_RLAST,
        m_axi_gmem2_RID => m_axi_gmem2_RID,
        m_axi_gmem2_RFIFONUM => m_axi_gmem2_RFIFONUM,
        m_axi_gmem2_RUSER => m_axi_gmem2_RUSER,
        m_axi_gmem2_RRESP => m_axi_gmem2_RRESP,
        m_axi_gmem2_BVALID => ap_const_logic_0,
        m_axi_gmem2_BREADY => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_BREADY,
        m_axi_gmem2_BRESP => ap_const_lv2_0,
        m_axi_gmem2_BID => ap_const_lv1_0,
        m_axi_gmem2_BUSER => ap_const_lv1_0,
        ldata_din => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_ldata_din,
        ldata_num_data_valid => ap_const_lv2_0,
        ldata_fifo_cap => ap_const_lv2_0,
        ldata_full_n => ldata_full_n,
        ldata_write => grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_ldata_write,
        sext_ln1028 => trunc_ln_reg_448,
        cols_addrbound => cols_addrbound_reg_416);

    mul_mul_11ns_11ns_22_3_1_U87 : component pp_pipeline_accel_mul_mul_11ns_11ns_22_3_1
    generic map (
        ID => 1,
        NUM_STAGE => 3,
        din0_WIDTH => 11,
        din1_WIDTH => 11,
        dout_WIDTH => 22)
    port map (
        clk => ap_clk,
        reset => ap_rst,
        din0 => grp_fu_329_p0,
        din1 => grp_fu_329_p1,
        ce => ap_const_logic_1,
        dout => grp_fu_329_p2);

    mul_mul_16ns_11ns_27_3_1_U88 : component pp_pipeline_accel_mul_mul_16ns_11ns_27_3_1
    generic map (
        ID => 1,
        NUM_STAGE => 3,
        din0_WIDTH => 16,
        din1_WIDTH => 11,
        dout_WIDTH => 27)
    port map (
        clk => ap_clk,
        reset => ap_rst,
        din0 => grp_fu_335_p0,
        din1 => grp_fu_335_p1,
        ce => ap_const_logic_1,
        dout => grp_fu_335_p2);

    mul_mul_20ns_11ns_31_4_1_U89 : component pp_pipeline_accel_mul_mul_20ns_11ns_31_4_1
    generic map (
        ID => 1,
        NUM_STAGE => 4,
        din0_WIDTH => 20,
        din1_WIDTH => 11,
        dout_WIDTH => 31)
    port map (
        clk => ap_clk,
        reset => ap_rst,
        din0 => grp_fu_342_p0,
        din1 => grp_fu_342_p1,
        ce => ap_const_logic_1,
        dout => grp_fu_342_p2);





    ap_CS_fsm_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_CS_fsm <= ap_ST_fsm_state1;
            else
                ap_CS_fsm <= ap_NS_fsm;
            end if;
        end if;
    end process;


    ap_done_reg_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                ap_done_reg <= ap_const_logic_0;
            else
                if ((ap_continue = ap_const_logic_1)) then 
                    ap_done_reg <= ap_const_logic_0;
                elsif (((icmp_ln1024_fu_274_p2 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_state6))) then 
                    ap_done_reg <= ap_const_logic_1;
                end if; 
            end if;
        end if;
    end process;


    grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_ap_start_reg_assign_proc : process(ap_clk)
    begin
        if (ap_clk'event and ap_clk =  '1') then
            if (ap_rst = '1') then
                grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_ap_start_reg <= ap_const_logic_0;
            else
                if ((ap_const_logic_1 = ap_CS_fsm_state80)) then 
                    grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_ap_start_reg <= ap_const_logic_1;
                elsif ((grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_ap_ready = ap_const_logic_1)) then 
                    grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_ap_start_reg <= ap_const_logic_0;
                end if; 
            end if;
        end if;
    end process;


    r_fu_116_assign_proc : process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if ((not(((ap_done_reg = ap_const_logic_1) or (ap_start = ap_const_logic_0) or (cols_c_full_n = ap_const_logic_0))) and (ap_const_logic_1 = ap_CS_fsm_state1))) then 
                r_fu_116 <= ap_const_lv11_0;
            elsif (((ap_const_boolean_0 = ap_block_state81_on_subcall_done) and (ap_const_logic_1 = ap_CS_fsm_state81))) then 
                r_fu_116 <= r_4_reg_438;
            end if; 
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if ((ap_const_logic_1 = ap_CS_fsm_state5)) then
                cmp_i82_i_reg_421 <= cmp_i82_i_fu_257_p2;
                cols_addrbound_reg_416 <= add_ln587_fu_211_p2(25 downto 6);
                    zext_ln1028_1_reg_430(19 downto 0) <= zext_ln1028_1_fu_267_p1(19 downto 0);
                    zext_ln1028_reg_425(19 downto 0) <= zext_ln1028_fu_263_p1(19 downto 0);
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if ((ap_const_logic_1 = ap_CS_fsm_state1)) then
                cols_int16_reg_366 <= cols_int16_fu_174_p1;
                icmp_ln1021_reg_371 <= icmp_ln1021_fu_178_p2;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if ((ap_const_logic_1 = ap_CS_fsm_state6)) then
                r_4_reg_438 <= r_4_fu_279_p2;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if ((ap_const_logic_1 = ap_CS_fsm_state4)) then
                ret_V_36_reg_396 <= grp_fu_329_p2;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((ap_const_logic_1 = ap_CS_fsm_state4) and (icmp_ln1021_reg_371 = ap_const_lv1_0))) then
                trunc_ln1540_reg_401 <= trunc_ln1540_fu_201_p1;
            end if;
        end if;
    end process;
    process (ap_clk)
    begin
        if (ap_clk'event and ap_clk = '1') then
            if (((cmp_i82_i_reg_421 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_state9))) then
                trunc_ln_reg_448 <= empty_229_fu_300_p2(63 downto 3);
            end if;
        end if;
    end process;
    zext_ln1028_reg_425(30 downto 20) <= "00000000000";
    zext_ln1028_1_reg_430(31 downto 20) <= "000000000000";

    ap_NS_fsm_assign_proc : process (ap_start, ap_done_reg, ap_CS_fsm, ap_CS_fsm_state1, m_axi_gmem2_ARREADY, cols_c_full_n, ap_CS_fsm_state10, cmp_i82_i_reg_421, ap_CS_fsm_state6, icmp_ln1024_fu_274_p2, ap_CS_fsm_state9, ap_CS_fsm_state81, ap_block_state81_on_subcall_done)
    begin
        case ap_CS_fsm is
            when ap_ST_fsm_state1 => 
                if ((not(((ap_done_reg = ap_const_logic_1) or (ap_start = ap_const_logic_0) or (cols_c_full_n = ap_const_logic_0))) and (ap_const_logic_1 = ap_CS_fsm_state1))) then
                    ap_NS_fsm <= ap_ST_fsm_state2;
                else
                    ap_NS_fsm <= ap_ST_fsm_state1;
                end if;
            when ap_ST_fsm_state2 => 
                ap_NS_fsm <= ap_ST_fsm_state3;
            when ap_ST_fsm_state3 => 
                ap_NS_fsm <= ap_ST_fsm_state4;
            when ap_ST_fsm_state4 => 
                ap_NS_fsm <= ap_ST_fsm_state5;
            when ap_ST_fsm_state5 => 
                ap_NS_fsm <= ap_ST_fsm_state6;
            when ap_ST_fsm_state6 => 
                if (((icmp_ln1024_fu_274_p2 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_state6))) then
                    ap_NS_fsm <= ap_ST_fsm_state1;
                else
                    ap_NS_fsm <= ap_ST_fsm_state7;
                end if;
            when ap_ST_fsm_state7 => 
                ap_NS_fsm <= ap_ST_fsm_state8;
            when ap_ST_fsm_state8 => 
                ap_NS_fsm <= ap_ST_fsm_state9;
            when ap_ST_fsm_state9 => 
                if (((cmp_i82_i_reg_421 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_state9))) then
                    ap_NS_fsm <= ap_ST_fsm_state81;
                else
                    ap_NS_fsm <= ap_ST_fsm_state10;
                end if;
            when ap_ST_fsm_state10 => 
                if (((ap_const_logic_1 = ap_CS_fsm_state10) and (m_axi_gmem2_ARREADY = ap_const_logic_1))) then
                    ap_NS_fsm <= ap_ST_fsm_state11;
                else
                    ap_NS_fsm <= ap_ST_fsm_state10;
                end if;
            when ap_ST_fsm_state11 => 
                ap_NS_fsm <= ap_ST_fsm_state12;
            when ap_ST_fsm_state12 => 
                ap_NS_fsm <= ap_ST_fsm_state13;
            when ap_ST_fsm_state13 => 
                ap_NS_fsm <= ap_ST_fsm_state14;
            when ap_ST_fsm_state14 => 
                ap_NS_fsm <= ap_ST_fsm_state15;
            when ap_ST_fsm_state15 => 
                ap_NS_fsm <= ap_ST_fsm_state16;
            when ap_ST_fsm_state16 => 
                ap_NS_fsm <= ap_ST_fsm_state17;
            when ap_ST_fsm_state17 => 
                ap_NS_fsm <= ap_ST_fsm_state18;
            when ap_ST_fsm_state18 => 
                ap_NS_fsm <= ap_ST_fsm_state19;
            when ap_ST_fsm_state19 => 
                ap_NS_fsm <= ap_ST_fsm_state20;
            when ap_ST_fsm_state20 => 
                ap_NS_fsm <= ap_ST_fsm_state21;
            when ap_ST_fsm_state21 => 
                ap_NS_fsm <= ap_ST_fsm_state22;
            when ap_ST_fsm_state22 => 
                ap_NS_fsm <= ap_ST_fsm_state23;
            when ap_ST_fsm_state23 => 
                ap_NS_fsm <= ap_ST_fsm_state24;
            when ap_ST_fsm_state24 => 
                ap_NS_fsm <= ap_ST_fsm_state25;
            when ap_ST_fsm_state25 => 
                ap_NS_fsm <= ap_ST_fsm_state26;
            when ap_ST_fsm_state26 => 
                ap_NS_fsm <= ap_ST_fsm_state27;
            when ap_ST_fsm_state27 => 
                ap_NS_fsm <= ap_ST_fsm_state28;
            when ap_ST_fsm_state28 => 
                ap_NS_fsm <= ap_ST_fsm_state29;
            when ap_ST_fsm_state29 => 
                ap_NS_fsm <= ap_ST_fsm_state30;
            when ap_ST_fsm_state30 => 
                ap_NS_fsm <= ap_ST_fsm_state31;
            when ap_ST_fsm_state31 => 
                ap_NS_fsm <= ap_ST_fsm_state32;
            when ap_ST_fsm_state32 => 
                ap_NS_fsm <= ap_ST_fsm_state33;
            when ap_ST_fsm_state33 => 
                ap_NS_fsm <= ap_ST_fsm_state34;
            when ap_ST_fsm_state34 => 
                ap_NS_fsm <= ap_ST_fsm_state35;
            when ap_ST_fsm_state35 => 
                ap_NS_fsm <= ap_ST_fsm_state36;
            when ap_ST_fsm_state36 => 
                ap_NS_fsm <= ap_ST_fsm_state37;
            when ap_ST_fsm_state37 => 
                ap_NS_fsm <= ap_ST_fsm_state38;
            when ap_ST_fsm_state38 => 
                ap_NS_fsm <= ap_ST_fsm_state39;
            when ap_ST_fsm_state39 => 
                ap_NS_fsm <= ap_ST_fsm_state40;
            when ap_ST_fsm_state40 => 
                ap_NS_fsm <= ap_ST_fsm_state41;
            when ap_ST_fsm_state41 => 
                ap_NS_fsm <= ap_ST_fsm_state42;
            when ap_ST_fsm_state42 => 
                ap_NS_fsm <= ap_ST_fsm_state43;
            when ap_ST_fsm_state43 => 
                ap_NS_fsm <= ap_ST_fsm_state44;
            when ap_ST_fsm_state44 => 
                ap_NS_fsm <= ap_ST_fsm_state45;
            when ap_ST_fsm_state45 => 
                ap_NS_fsm <= ap_ST_fsm_state46;
            when ap_ST_fsm_state46 => 
                ap_NS_fsm <= ap_ST_fsm_state47;
            when ap_ST_fsm_state47 => 
                ap_NS_fsm <= ap_ST_fsm_state48;
            when ap_ST_fsm_state48 => 
                ap_NS_fsm <= ap_ST_fsm_state49;
            when ap_ST_fsm_state49 => 
                ap_NS_fsm <= ap_ST_fsm_state50;
            when ap_ST_fsm_state50 => 
                ap_NS_fsm <= ap_ST_fsm_state51;
            when ap_ST_fsm_state51 => 
                ap_NS_fsm <= ap_ST_fsm_state52;
            when ap_ST_fsm_state52 => 
                ap_NS_fsm <= ap_ST_fsm_state53;
            when ap_ST_fsm_state53 => 
                ap_NS_fsm <= ap_ST_fsm_state54;
            when ap_ST_fsm_state54 => 
                ap_NS_fsm <= ap_ST_fsm_state55;
            when ap_ST_fsm_state55 => 
                ap_NS_fsm <= ap_ST_fsm_state56;
            when ap_ST_fsm_state56 => 
                ap_NS_fsm <= ap_ST_fsm_state57;
            when ap_ST_fsm_state57 => 
                ap_NS_fsm <= ap_ST_fsm_state58;
            when ap_ST_fsm_state58 => 
                ap_NS_fsm <= ap_ST_fsm_state59;
            when ap_ST_fsm_state59 => 
                ap_NS_fsm <= ap_ST_fsm_state60;
            when ap_ST_fsm_state60 => 
                ap_NS_fsm <= ap_ST_fsm_state61;
            when ap_ST_fsm_state61 => 
                ap_NS_fsm <= ap_ST_fsm_state62;
            when ap_ST_fsm_state62 => 
                ap_NS_fsm <= ap_ST_fsm_state63;
            when ap_ST_fsm_state63 => 
                ap_NS_fsm <= ap_ST_fsm_state64;
            when ap_ST_fsm_state64 => 
                ap_NS_fsm <= ap_ST_fsm_state65;
            when ap_ST_fsm_state65 => 
                ap_NS_fsm <= ap_ST_fsm_state66;
            when ap_ST_fsm_state66 => 
                ap_NS_fsm <= ap_ST_fsm_state67;
            when ap_ST_fsm_state67 => 
                ap_NS_fsm <= ap_ST_fsm_state68;
            when ap_ST_fsm_state68 => 
                ap_NS_fsm <= ap_ST_fsm_state69;
            when ap_ST_fsm_state69 => 
                ap_NS_fsm <= ap_ST_fsm_state70;
            when ap_ST_fsm_state70 => 
                ap_NS_fsm <= ap_ST_fsm_state71;
            when ap_ST_fsm_state71 => 
                ap_NS_fsm <= ap_ST_fsm_state72;
            when ap_ST_fsm_state72 => 
                ap_NS_fsm <= ap_ST_fsm_state73;
            when ap_ST_fsm_state73 => 
                ap_NS_fsm <= ap_ST_fsm_state74;
            when ap_ST_fsm_state74 => 
                ap_NS_fsm <= ap_ST_fsm_state75;
            when ap_ST_fsm_state75 => 
                ap_NS_fsm <= ap_ST_fsm_state76;
            when ap_ST_fsm_state76 => 
                ap_NS_fsm <= ap_ST_fsm_state77;
            when ap_ST_fsm_state77 => 
                ap_NS_fsm <= ap_ST_fsm_state78;
            when ap_ST_fsm_state78 => 
                ap_NS_fsm <= ap_ST_fsm_state79;
            when ap_ST_fsm_state79 => 
                ap_NS_fsm <= ap_ST_fsm_state80;
            when ap_ST_fsm_state80 => 
                ap_NS_fsm <= ap_ST_fsm_state81;
            when ap_ST_fsm_state81 => 
                if (((ap_const_boolean_0 = ap_block_state81_on_subcall_done) and (ap_const_logic_1 = ap_CS_fsm_state81))) then
                    ap_NS_fsm <= ap_ST_fsm_state6;
                else
                    ap_NS_fsm <= ap_ST_fsm_state81;
                end if;
            when others =>  
                ap_NS_fsm <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
        end case;
    end process;
    add_ln587_1_fu_234_p2 <= std_logic_vector(unsigned(ret_V_7_fu_227_p3) + unsigned(ap_const_lv26_3F));
    add_ln587_fu_211_p2 <= std_logic_vector(unsigned(ret_V_fu_204_p3) + unsigned(ap_const_lv26_3F));
    addrbound_V_fu_250_p3 <= 
        cols_addrbound_fu_217_p4 when (icmp_ln1021_reg_371(0) = '1') else 
        stride_addrbound_fu_240_p4;
    ap_CS_fsm_state1 <= ap_CS_fsm(0);
    ap_CS_fsm_state10 <= ap_CS_fsm(9);
    ap_CS_fsm_state2 <= ap_CS_fsm(1);
    ap_CS_fsm_state4 <= ap_CS_fsm(3);
    ap_CS_fsm_state5 <= ap_CS_fsm(4);
    ap_CS_fsm_state6 <= ap_CS_fsm(5);
    ap_CS_fsm_state80 <= ap_CS_fsm(79);
    ap_CS_fsm_state81 <= ap_CS_fsm(80);
    ap_CS_fsm_state9 <= ap_CS_fsm(8);

    ap_ST_fsm_state10_blk_assign_proc : process(m_axi_gmem2_ARREADY)
    begin
        if ((m_axi_gmem2_ARREADY = ap_const_logic_0)) then 
            ap_ST_fsm_state10_blk <= ap_const_logic_1;
        else 
            ap_ST_fsm_state10_blk <= ap_const_logic_0;
        end if; 
    end process;

    ap_ST_fsm_state11_blk <= ap_const_logic_0;
    ap_ST_fsm_state12_blk <= ap_const_logic_0;
    ap_ST_fsm_state13_blk <= ap_const_logic_0;
    ap_ST_fsm_state14_blk <= ap_const_logic_0;
    ap_ST_fsm_state15_blk <= ap_const_logic_0;
    ap_ST_fsm_state16_blk <= ap_const_logic_0;
    ap_ST_fsm_state17_blk <= ap_const_logic_0;
    ap_ST_fsm_state18_blk <= ap_const_logic_0;
    ap_ST_fsm_state19_blk <= ap_const_logic_0;

    ap_ST_fsm_state1_blk_assign_proc : process(ap_start, ap_done_reg, cols_c_full_n)
    begin
        if (((ap_done_reg = ap_const_logic_1) or (ap_start = ap_const_logic_0) or (cols_c_full_n = ap_const_logic_0))) then 
            ap_ST_fsm_state1_blk <= ap_const_logic_1;
        else 
            ap_ST_fsm_state1_blk <= ap_const_logic_0;
        end if; 
    end process;

    ap_ST_fsm_state20_blk <= ap_const_logic_0;
    ap_ST_fsm_state21_blk <= ap_const_logic_0;
    ap_ST_fsm_state22_blk <= ap_const_logic_0;
    ap_ST_fsm_state23_blk <= ap_const_logic_0;
    ap_ST_fsm_state24_blk <= ap_const_logic_0;
    ap_ST_fsm_state25_blk <= ap_const_logic_0;
    ap_ST_fsm_state26_blk <= ap_const_logic_0;
    ap_ST_fsm_state27_blk <= ap_const_logic_0;
    ap_ST_fsm_state28_blk <= ap_const_logic_0;
    ap_ST_fsm_state29_blk <= ap_const_logic_0;
    ap_ST_fsm_state2_blk <= ap_const_logic_0;
    ap_ST_fsm_state30_blk <= ap_const_logic_0;
    ap_ST_fsm_state31_blk <= ap_const_logic_0;
    ap_ST_fsm_state32_blk <= ap_const_logic_0;
    ap_ST_fsm_state33_blk <= ap_const_logic_0;
    ap_ST_fsm_state34_blk <= ap_const_logic_0;
    ap_ST_fsm_state35_blk <= ap_const_logic_0;
    ap_ST_fsm_state36_blk <= ap_const_logic_0;
    ap_ST_fsm_state37_blk <= ap_const_logic_0;
    ap_ST_fsm_state38_blk <= ap_const_logic_0;
    ap_ST_fsm_state39_blk <= ap_const_logic_0;
    ap_ST_fsm_state3_blk <= ap_const_logic_0;
    ap_ST_fsm_state40_blk <= ap_const_logic_0;
    ap_ST_fsm_state41_blk <= ap_const_logic_0;
    ap_ST_fsm_state42_blk <= ap_const_logic_0;
    ap_ST_fsm_state43_blk <= ap_const_logic_0;
    ap_ST_fsm_state44_blk <= ap_const_logic_0;
    ap_ST_fsm_state45_blk <= ap_const_logic_0;
    ap_ST_fsm_state46_blk <= ap_const_logic_0;
    ap_ST_fsm_state47_blk <= ap_const_logic_0;
    ap_ST_fsm_state48_blk <= ap_const_logic_0;
    ap_ST_fsm_state49_blk <= ap_const_logic_0;
    ap_ST_fsm_state4_blk <= ap_const_logic_0;
    ap_ST_fsm_state50_blk <= ap_const_logic_0;
    ap_ST_fsm_state51_blk <= ap_const_logic_0;
    ap_ST_fsm_state52_blk <= ap_const_logic_0;
    ap_ST_fsm_state53_blk <= ap_const_logic_0;
    ap_ST_fsm_state54_blk <= ap_const_logic_0;
    ap_ST_fsm_state55_blk <= ap_const_logic_0;
    ap_ST_fsm_state56_blk <= ap_const_logic_0;
    ap_ST_fsm_state57_blk <= ap_const_logic_0;
    ap_ST_fsm_state58_blk <= ap_const_logic_0;
    ap_ST_fsm_state59_blk <= ap_const_logic_0;
    ap_ST_fsm_state5_blk <= ap_const_logic_0;
    ap_ST_fsm_state60_blk <= ap_const_logic_0;
    ap_ST_fsm_state61_blk <= ap_const_logic_0;
    ap_ST_fsm_state62_blk <= ap_const_logic_0;
    ap_ST_fsm_state63_blk <= ap_const_logic_0;
    ap_ST_fsm_state64_blk <= ap_const_logic_0;
    ap_ST_fsm_state65_blk <= ap_const_logic_0;
    ap_ST_fsm_state66_blk <= ap_const_logic_0;
    ap_ST_fsm_state67_blk <= ap_const_logic_0;
    ap_ST_fsm_state68_blk <= ap_const_logic_0;
    ap_ST_fsm_state69_blk <= ap_const_logic_0;
    ap_ST_fsm_state6_blk <= ap_const_logic_0;
    ap_ST_fsm_state70_blk <= ap_const_logic_0;
    ap_ST_fsm_state71_blk <= ap_const_logic_0;
    ap_ST_fsm_state72_blk <= ap_const_logic_0;
    ap_ST_fsm_state73_blk <= ap_const_logic_0;
    ap_ST_fsm_state74_blk <= ap_const_logic_0;
    ap_ST_fsm_state75_blk <= ap_const_logic_0;
    ap_ST_fsm_state76_blk <= ap_const_logic_0;
    ap_ST_fsm_state77_blk <= ap_const_logic_0;
    ap_ST_fsm_state78_blk <= ap_const_logic_0;
    ap_ST_fsm_state79_blk <= ap_const_logic_0;
    ap_ST_fsm_state7_blk <= ap_const_logic_0;
    ap_ST_fsm_state80_blk <= ap_const_logic_0;

    ap_ST_fsm_state81_blk_assign_proc : process(ap_block_state81_on_subcall_done)
    begin
        if ((ap_const_boolean_1 = ap_block_state81_on_subcall_done)) then 
            ap_ST_fsm_state81_blk <= ap_const_logic_1;
        else 
            ap_ST_fsm_state81_blk <= ap_const_logic_0;
        end if; 
    end process;

    ap_ST_fsm_state8_blk <= ap_const_logic_0;
    ap_ST_fsm_state9_blk <= ap_const_logic_0;

    ap_block_state1_assign_proc : process(ap_start, ap_done_reg, cols_c_full_n)
    begin
                ap_block_state1 <= ((ap_done_reg = ap_const_logic_1) or (ap_start = ap_const_logic_0) or (cols_c_full_n = ap_const_logic_0));
    end process;


    ap_block_state81_on_subcall_done_assign_proc : process(cmp_i82_i_reg_421, grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_ap_done)
    begin
                ap_block_state81_on_subcall_done <= ((grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_ap_done = ap_const_logic_0) and (cmp_i82_i_reg_421 = ap_const_lv1_0));
    end process;


    ap_done_assign_proc : process(ap_done_reg, ap_CS_fsm_state6, icmp_ln1024_fu_274_p2)
    begin
        if (((icmp_ln1024_fu_274_p2 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_state6))) then 
            ap_done <= ap_const_logic_1;
        else 
            ap_done <= ap_done_reg;
        end if; 
    end process;


    ap_idle_assign_proc : process(ap_start, ap_CS_fsm_state1)
    begin
        if (((ap_start = ap_const_logic_0) and (ap_const_logic_1 = ap_CS_fsm_state1))) then 
            ap_idle <= ap_const_logic_1;
        else 
            ap_idle <= ap_const_logic_0;
        end if; 
    end process;


    ap_ready_assign_proc : process(ap_CS_fsm_state6, icmp_ln1024_fu_274_p2)
    begin
        if (((icmp_ln1024_fu_274_p2 = ap_const_lv1_1) and (ap_const_logic_1 = ap_CS_fsm_state6))) then 
            ap_ready <= ap_const_logic_1;
        else 
            ap_ready <= ap_const_logic_0;
        end if; 
    end process;

    cmp_i82_i_fu_257_p2 <= "1" when (cols_addrbound_fu_217_p4 = ap_const_lv20_0) else "0";
    cols_addrbound_fu_217_p4 <= add_ln587_fu_211_p2(25 downto 6);

    cols_c_blk_n_assign_proc : process(ap_start, ap_done_reg, ap_CS_fsm_state1, cols_c_full_n)
    begin
        if ((not(((ap_done_reg = ap_const_logic_1) or (ap_start = ap_const_logic_0))) and (ap_const_logic_1 = ap_CS_fsm_state1))) then 
            cols_c_blk_n <= cols_c_full_n;
        else 
            cols_c_blk_n <= ap_const_logic_1;
        end if; 
    end process;

    cols_c_din <= cols;

    cols_c_write_assign_proc : process(ap_start, ap_done_reg, ap_CS_fsm_state1, cols_c_full_n)
    begin
        if ((not(((ap_done_reg = ap_const_logic_1) or (ap_start = ap_const_logic_0) or (cols_c_full_n = ap_const_logic_0))) and (ap_const_logic_1 = ap_CS_fsm_state1))) then 
            cols_c_write <= ap_const_logic_1;
        else 
            cols_c_write <= ap_const_logic_0;
        end if; 
    end process;

    cols_int16_fu_174_p1 <= stride(16 - 1 downto 0);
    empty_229_fu_300_p2 <= std_logic_vector(unsigned(p_cast2_i_fu_296_p1) + unsigned(din));

    gmem2_blk_n_AR_assign_proc : process(m_axi_gmem2_ARREADY, ap_CS_fsm_state10)
    begin
        if ((ap_const_logic_1 = ap_CS_fsm_state10)) then 
            gmem2_blk_n_AR <= m_axi_gmem2_ARREADY;
        else 
            gmem2_blk_n_AR <= ap_const_logic_1;
        end if; 
    end process;

    grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_ap_start <= grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_ap_start_reg;
    grp_fu_329_p0 <= grp_fu_329_p00(11 - 1 downto 0);
    grp_fu_329_p00 <= std_logic_vector(IEEE.numeric_std.resize(unsigned(cols),22));
    grp_fu_329_p1 <= grp_fu_329_p10(11 - 1 downto 0);
    grp_fu_329_p10 <= std_logic_vector(IEEE.numeric_std.resize(unsigned(p_read),22));
    grp_fu_335_p0 <= grp_fu_335_p00(16 - 1 downto 0);
    grp_fu_335_p00 <= std_logic_vector(IEEE.numeric_std.resize(unsigned(cols_int16_reg_366),27));
    grp_fu_335_p1 <= grp_fu_335_p10(11 - 1 downto 0);
    grp_fu_335_p10 <= std_logic_vector(IEEE.numeric_std.resize(unsigned(p_read),27));
    grp_fu_342_p0 <= zext_ln1028_reg_425(20 - 1 downto 0);
    grp_fu_342_p1 <= grp_fu_342_p10(11 - 1 downto 0);
    grp_fu_342_p10 <= std_logic_vector(IEEE.numeric_std.resize(unsigned(r_fu_116),31));
    icmp_ln1021_fu_178_p2 <= "1" when (stride = ap_const_lv32_FFFFFFFF) else "0";
    icmp_ln1024_fu_274_p2 <= "1" when (r_fu_116 = p_read1) else "0";
    ldata_din <= grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_ldata_din;

    ldata_write_assign_proc : process(cmp_i82_i_reg_421, grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_ldata_write, ap_CS_fsm_state81)
    begin
        if (((cmp_i82_i_reg_421 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_state81))) then 
            ldata_write <= grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_ldata_write;
        else 
            ldata_write <= ap_const_logic_0;
        end if; 
    end process;


    m_axi_gmem2_ARADDR_assign_proc : process(m_axi_gmem2_ARREADY, ap_CS_fsm_state10, cmp_i82_i_reg_421, grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARADDR, ap_CS_fsm_state80, ap_CS_fsm_state81, sext_ln1028_fu_315_p1)
    begin
        if (((ap_const_logic_1 = ap_CS_fsm_state10) and (m_axi_gmem2_ARREADY = ap_const_logic_1))) then 
            m_axi_gmem2_ARADDR <= sext_ln1028_fu_315_p1;
        elsif (((ap_const_logic_1 = ap_CS_fsm_state80) or ((cmp_i82_i_reg_421 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_state81)))) then 
            m_axi_gmem2_ARADDR <= grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARADDR;
        else 
            m_axi_gmem2_ARADDR <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
        end if; 
    end process;


    m_axi_gmem2_ARBURST_assign_proc : process(cmp_i82_i_reg_421, grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARBURST, ap_CS_fsm_state80, ap_CS_fsm_state81)
    begin
        if (((ap_const_logic_1 = ap_CS_fsm_state80) or ((cmp_i82_i_reg_421 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_state81)))) then 
            m_axi_gmem2_ARBURST <= grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARBURST;
        else 
            m_axi_gmem2_ARBURST <= ap_const_lv2_0;
        end if; 
    end process;


    m_axi_gmem2_ARCACHE_assign_proc : process(cmp_i82_i_reg_421, grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARCACHE, ap_CS_fsm_state80, ap_CS_fsm_state81)
    begin
        if (((ap_const_logic_1 = ap_CS_fsm_state80) or ((cmp_i82_i_reg_421 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_state81)))) then 
            m_axi_gmem2_ARCACHE <= grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARCACHE;
        else 
            m_axi_gmem2_ARCACHE <= ap_const_lv4_0;
        end if; 
    end process;


    m_axi_gmem2_ARID_assign_proc : process(cmp_i82_i_reg_421, grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARID, ap_CS_fsm_state80, ap_CS_fsm_state81)
    begin
        if (((ap_const_logic_1 = ap_CS_fsm_state80) or ((cmp_i82_i_reg_421 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_state81)))) then 
            m_axi_gmem2_ARID <= grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARID;
        else 
            m_axi_gmem2_ARID <= ap_const_lv1_0;
        end if; 
    end process;


    m_axi_gmem2_ARLEN_assign_proc : process(m_axi_gmem2_ARREADY, ap_CS_fsm_state10, cmp_i82_i_reg_421, zext_ln1028_1_reg_430, grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARLEN, ap_CS_fsm_state80, ap_CS_fsm_state81)
    begin
        if (((ap_const_logic_1 = ap_CS_fsm_state10) and (m_axi_gmem2_ARREADY = ap_const_logic_1))) then 
            m_axi_gmem2_ARLEN <= zext_ln1028_1_reg_430;
        elsif (((ap_const_logic_1 = ap_CS_fsm_state80) or ((cmp_i82_i_reg_421 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_state81)))) then 
            m_axi_gmem2_ARLEN <= grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARLEN;
        else 
            m_axi_gmem2_ARLEN <= "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";
        end if; 
    end process;


    m_axi_gmem2_ARLOCK_assign_proc : process(cmp_i82_i_reg_421, grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARLOCK, ap_CS_fsm_state80, ap_CS_fsm_state81)
    begin
        if (((ap_const_logic_1 = ap_CS_fsm_state80) or ((cmp_i82_i_reg_421 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_state81)))) then 
            m_axi_gmem2_ARLOCK <= grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARLOCK;
        else 
            m_axi_gmem2_ARLOCK <= ap_const_lv2_0;
        end if; 
    end process;


    m_axi_gmem2_ARPROT_assign_proc : process(cmp_i82_i_reg_421, grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARPROT, ap_CS_fsm_state80, ap_CS_fsm_state81)
    begin
        if (((ap_const_logic_1 = ap_CS_fsm_state80) or ((cmp_i82_i_reg_421 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_state81)))) then 
            m_axi_gmem2_ARPROT <= grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARPROT;
        else 
            m_axi_gmem2_ARPROT <= ap_const_lv3_0;
        end if; 
    end process;


    m_axi_gmem2_ARQOS_assign_proc : process(cmp_i82_i_reg_421, grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARQOS, ap_CS_fsm_state80, ap_CS_fsm_state81)
    begin
        if (((ap_const_logic_1 = ap_CS_fsm_state80) or ((cmp_i82_i_reg_421 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_state81)))) then 
            m_axi_gmem2_ARQOS <= grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARQOS;
        else 
            m_axi_gmem2_ARQOS <= ap_const_lv4_0;
        end if; 
    end process;


    m_axi_gmem2_ARREGION_assign_proc : process(cmp_i82_i_reg_421, grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARREGION, ap_CS_fsm_state80, ap_CS_fsm_state81)
    begin
        if (((ap_const_logic_1 = ap_CS_fsm_state80) or ((cmp_i82_i_reg_421 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_state81)))) then 
            m_axi_gmem2_ARREGION <= grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARREGION;
        else 
            m_axi_gmem2_ARREGION <= ap_const_lv4_0;
        end if; 
    end process;


    m_axi_gmem2_ARSIZE_assign_proc : process(cmp_i82_i_reg_421, grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARSIZE, ap_CS_fsm_state80, ap_CS_fsm_state81)
    begin
        if (((ap_const_logic_1 = ap_CS_fsm_state80) or ((cmp_i82_i_reg_421 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_state81)))) then 
            m_axi_gmem2_ARSIZE <= grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARSIZE;
        else 
            m_axi_gmem2_ARSIZE <= ap_const_lv3_0;
        end if; 
    end process;


    m_axi_gmem2_ARUSER_assign_proc : process(cmp_i82_i_reg_421, grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARUSER, ap_CS_fsm_state80, ap_CS_fsm_state81)
    begin
        if (((ap_const_logic_1 = ap_CS_fsm_state80) or ((cmp_i82_i_reg_421 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_state81)))) then 
            m_axi_gmem2_ARUSER <= grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARUSER;
        else 
            m_axi_gmem2_ARUSER <= ap_const_lv1_0;
        end if; 
    end process;


    m_axi_gmem2_ARVALID_assign_proc : process(m_axi_gmem2_ARREADY, ap_CS_fsm_state10, cmp_i82_i_reg_421, grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARVALID, ap_CS_fsm_state80, ap_CS_fsm_state81)
    begin
        if (((ap_const_logic_1 = ap_CS_fsm_state10) and (m_axi_gmem2_ARREADY = ap_const_logic_1))) then 
            m_axi_gmem2_ARVALID <= ap_const_logic_1;
        elsif (((ap_const_logic_1 = ap_CS_fsm_state80) or ((cmp_i82_i_reg_421 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_state81)))) then 
            m_axi_gmem2_ARVALID <= grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_ARVALID;
        else 
            m_axi_gmem2_ARVALID <= ap_const_logic_0;
        end if; 
    end process;

    m_axi_gmem2_AWADDR <= ap_const_lv64_0;
    m_axi_gmem2_AWBURST <= ap_const_lv2_0;
    m_axi_gmem2_AWCACHE <= ap_const_lv4_0;
    m_axi_gmem2_AWID <= ap_const_lv1_0;
    m_axi_gmem2_AWLEN <= ap_const_lv32_0;
    m_axi_gmem2_AWLOCK <= ap_const_lv2_0;
    m_axi_gmem2_AWPROT <= ap_const_lv3_0;
    m_axi_gmem2_AWQOS <= ap_const_lv4_0;
    m_axi_gmem2_AWREGION <= ap_const_lv4_0;
    m_axi_gmem2_AWSIZE <= ap_const_lv3_0;
    m_axi_gmem2_AWUSER <= ap_const_lv1_0;
    m_axi_gmem2_AWVALID <= ap_const_logic_0;
    m_axi_gmem2_BREADY <= ap_const_logic_0;

    m_axi_gmem2_RREADY_assign_proc : process(cmp_i82_i_reg_421, grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_RREADY, ap_CS_fsm_state80, ap_CS_fsm_state81)
    begin
        if (((ap_const_logic_1 = ap_CS_fsm_state80) or ((cmp_i82_i_reg_421 = ap_const_lv1_0) and (ap_const_logic_1 = ap_CS_fsm_state81)))) then 
            m_axi_gmem2_RREADY <= grp_Axi2AxiStream_Pipeline_VITIS_LOOP_1028_1_fu_164_m_axi_gmem2_RREADY;
        else 
            m_axi_gmem2_RREADY <= ap_const_logic_0;
        end if; 
    end process;

    m_axi_gmem2_WDATA <= ap_const_lv64_0;
    m_axi_gmem2_WID <= ap_const_lv1_0;
    m_axi_gmem2_WLAST <= ap_const_logic_0;
    m_axi_gmem2_WSTRB <= ap_const_lv8_0;
    m_axi_gmem2_WUSER <= ap_const_lv1_0;
    m_axi_gmem2_WVALID <= ap_const_logic_0;
    p_cast2_i_fu_296_p1 <= std_logic_vector(IEEE.numeric_std.resize(unsigned(tmp_s_fu_289_p3),64));
    r_4_fu_279_p2 <= std_logic_vector(unsigned(r_fu_116) + unsigned(ap_const_lv11_1));
    ret_V_7_fu_227_p3 <= (trunc_ln1540_reg_401 & ap_const_lv4_0);
    ret_V_fu_204_p3 <= (ret_V_36_reg_396 & ap_const_lv4_0);
        sext_ln1028_fu_315_p1 <= std_logic_vector(IEEE.numeric_std.resize(signed(trunc_ln_reg_448),64));

    stride_addrbound_fu_240_p4 <= add_ln587_1_fu_234_p2(25 downto 6);
    tmp_s_fu_289_p1 <= grp_fu_342_p2;
    tmp_s_fu_289_p3 <= (tmp_s_fu_289_p1 & ap_const_lv3_0);
    trunc_ln1540_fu_201_p0 <= grp_fu_335_p2;
    trunc_ln1540_fu_201_p1 <= trunc_ln1540_fu_201_p0(22 - 1 downto 0);
    zext_ln1028_1_fu_267_p1 <= std_logic_vector(IEEE.numeric_std.resize(unsigned(cols_addrbound_fu_217_p4),32));
    zext_ln1028_fu_263_p1 <= std_logic_vector(IEEE.numeric_std.resize(unsigned(addrbound_V_fu_250_p3),31));
end behav;
