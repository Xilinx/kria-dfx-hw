// Copyright (C) 2022, Advanced Micro Devices, Inc. All rights reserved.
// SPDX-License-Identifier: MIT
// ==============================================================
// Version: 2022.1.0
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module testEnc_process_r (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        p_read,
        p_read1,
        p_read2,
        p_read3,
        p_read4,
        p_read5,
        p_read6,
        p_read7,
        p_read8,
        p_read9,
        p_read10,
        plaintext,
        ap_return
);

parameter    ap_ST_fsm_pp0_stage0 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [127:0] p_read;
input  [127:0] p_read1;
input  [127:0] p_read2;
input  [127:0] p_read3;
input  [127:0] p_read4;
input  [127:0] p_read5;
input  [127:0] p_read6;
input  [127:0] p_read7;
input  [127:0] p_read8;
input  [127:0] p_read9;
input  [127:0] p_read10;
input  [127:0] plaintext;
output  [127:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;

(* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg    ap_enable_reg_pp0_iter5;
reg    ap_enable_reg_pp0_iter6;
reg    ap_enable_reg_pp0_iter7;
reg    ap_enable_reg_pp0_iter8;
reg    ap_enable_reg_pp0_iter9;
reg    ap_enable_reg_pp0_iter10;
reg    ap_enable_reg_pp0_iter11;
reg    ap_enable_reg_pp0_iter12;
reg    ap_enable_reg_pp0_iter13;
reg    ap_enable_reg_pp0_iter14;
reg    ap_enable_reg_pp0_iter15;
reg    ap_enable_reg_pp0_iter16;
reg    ap_enable_reg_pp0_iter17;
reg    ap_enable_reg_pp0_iter18;
reg    ap_enable_reg_pp0_iter19;
reg    ap_idle_pp0;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_state4_pp0_stage0_iter3;
wire    ap_block_state5_pp0_stage0_iter4;
wire    ap_block_state6_pp0_stage0_iter5;
wire    ap_block_state7_pp0_stage0_iter6;
wire    ap_block_state8_pp0_stage0_iter7;
wire    ap_block_state9_pp0_stage0_iter8;
wire    ap_block_state10_pp0_stage0_iter9;
wire    ap_block_state11_pp0_stage0_iter10;
wire    ap_block_state12_pp0_stage0_iter11;
wire    ap_block_state13_pp0_stage0_iter12;
wire    ap_block_state14_pp0_stage0_iter13;
wire    ap_block_state15_pp0_stage0_iter14;
wire    ap_block_state16_pp0_stage0_iter15;
wire    ap_block_state17_pp0_stage0_iter16;
wire    ap_block_state18_pp0_stage0_iter17;
wire    ap_block_state19_pp0_stage0_iter18;
wire    ap_block_state20_pp0_stage0_iter19;
wire    ap_block_pp0_stage0_subdone;
wire   [7:0] cipher_0_ssbox_address0;
reg    cipher_0_ssbox_ce0;
wire   [7:0] cipher_0_ssbox_q0;
wire   [7:0] cipher_0_ssbox_address1;
reg    cipher_0_ssbox_ce1;
wire   [7:0] cipher_0_ssbox_q1;
wire   [7:0] cipher_0_ssbox_address2;
reg    cipher_0_ssbox_ce2;
wire   [7:0] cipher_0_ssbox_q2;
wire   [7:0] cipher_0_ssbox_address3;
reg    cipher_0_ssbox_ce3;
wire   [7:0] cipher_0_ssbox_q3;
wire   [7:0] cipher_0_ssbox_address4;
reg    cipher_0_ssbox_ce4;
wire   [7:0] cipher_0_ssbox_q4;
wire   [7:0] cipher_0_ssbox_address5;
reg    cipher_0_ssbox_ce5;
wire   [7:0] cipher_0_ssbox_q5;
wire   [7:0] cipher_0_ssbox_address6;
reg    cipher_0_ssbox_ce6;
wire   [7:0] cipher_0_ssbox_q6;
wire   [7:0] cipher_0_ssbox_address7;
reg    cipher_0_ssbox_ce7;
wire   [7:0] cipher_0_ssbox_q7;
wire   [7:0] cipher_0_ssbox_address8;
reg    cipher_0_ssbox_ce8;
wire   [7:0] cipher_0_ssbox_q8;
wire   [7:0] cipher_0_ssbox_address9;
reg    cipher_0_ssbox_ce9;
wire   [7:0] cipher_0_ssbox_q9;
wire   [7:0] cipher_0_ssbox_address10;
reg    cipher_0_ssbox_ce10;
wire   [7:0] cipher_0_ssbox_q10;
wire   [7:0] cipher_0_ssbox_address11;
reg    cipher_0_ssbox_ce11;
wire   [7:0] cipher_0_ssbox_q11;
wire   [7:0] cipher_0_ssbox_address12;
reg    cipher_0_ssbox_ce12;
wire   [7:0] cipher_0_ssbox_q12;
wire   [7:0] cipher_0_ssbox_address13;
reg    cipher_0_ssbox_ce13;
wire   [7:0] cipher_0_ssbox_q13;
wire   [7:0] cipher_0_ssbox_address14;
reg    cipher_0_ssbox_ce14;
wire   [7:0] cipher_0_ssbox_q14;
wire   [7:0] cipher_0_ssbox_address15;
reg    cipher_0_ssbox_ce15;
wire   [7:0] cipher_0_ssbox_q15;
wire   [7:0] cipher_0_ssbox_address16;
reg    cipher_0_ssbox_ce16;
wire   [7:0] cipher_0_ssbox_q16;
wire   [7:0] cipher_0_ssbox_address17;
reg    cipher_0_ssbox_ce17;
wire   [7:0] cipher_0_ssbox_q17;
wire   [7:0] cipher_0_ssbox_address18;
reg    cipher_0_ssbox_ce18;
wire   [7:0] cipher_0_ssbox_q18;
wire   [7:0] cipher_0_ssbox_address19;
reg    cipher_0_ssbox_ce19;
wire   [7:0] cipher_0_ssbox_q19;
wire   [7:0] cipher_0_ssbox_address20;
reg    cipher_0_ssbox_ce20;
wire   [7:0] cipher_0_ssbox_q20;
wire   [7:0] cipher_0_ssbox_address21;
reg    cipher_0_ssbox_ce21;
wire   [7:0] cipher_0_ssbox_q21;
wire   [7:0] cipher_0_ssbox_address22;
reg    cipher_0_ssbox_ce22;
wire   [7:0] cipher_0_ssbox_q22;
wire   [7:0] cipher_0_ssbox_address23;
reg    cipher_0_ssbox_ce23;
wire   [7:0] cipher_0_ssbox_q23;
wire   [7:0] cipher_0_ssbox_address24;
reg    cipher_0_ssbox_ce24;
wire   [7:0] cipher_0_ssbox_q24;
wire   [7:0] cipher_0_ssbox_address25;
reg    cipher_0_ssbox_ce25;
wire   [7:0] cipher_0_ssbox_q25;
wire   [7:0] cipher_0_ssbox_address26;
reg    cipher_0_ssbox_ce26;
wire   [7:0] cipher_0_ssbox_q26;
wire   [7:0] cipher_0_ssbox_address27;
reg    cipher_0_ssbox_ce27;
wire   [7:0] cipher_0_ssbox_q27;
wire   [7:0] cipher_0_ssbox_address28;
reg    cipher_0_ssbox_ce28;
wire   [7:0] cipher_0_ssbox_q28;
wire   [7:0] cipher_0_ssbox_address29;
reg    cipher_0_ssbox_ce29;
wire   [7:0] cipher_0_ssbox_q29;
wire   [7:0] cipher_0_ssbox_address30;
reg    cipher_0_ssbox_ce30;
wire   [7:0] cipher_0_ssbox_q30;
wire   [7:0] cipher_0_ssbox_address31;
reg    cipher_0_ssbox_ce31;
wire   [7:0] cipher_0_ssbox_q31;
wire   [7:0] cipher_0_ssbox_address32;
reg    cipher_0_ssbox_ce32;
wire   [7:0] cipher_0_ssbox_q32;
wire   [7:0] cipher_0_ssbox_address33;
reg    cipher_0_ssbox_ce33;
wire   [7:0] cipher_0_ssbox_q33;
wire   [7:0] cipher_0_ssbox_address34;
reg    cipher_0_ssbox_ce34;
wire   [7:0] cipher_0_ssbox_q34;
wire   [7:0] cipher_0_ssbox_address35;
reg    cipher_0_ssbox_ce35;
wire   [7:0] cipher_0_ssbox_q35;
wire   [7:0] cipher_0_ssbox_address36;
reg    cipher_0_ssbox_ce36;
wire   [7:0] cipher_0_ssbox_q36;
wire   [7:0] cipher_0_ssbox_address37;
reg    cipher_0_ssbox_ce37;
wire   [7:0] cipher_0_ssbox_q37;
wire   [7:0] cipher_0_ssbox_address38;
reg    cipher_0_ssbox_ce38;
wire   [7:0] cipher_0_ssbox_q38;
wire   [7:0] cipher_0_ssbox_address39;
reg    cipher_0_ssbox_ce39;
wire   [7:0] cipher_0_ssbox_q39;
wire   [7:0] cipher_0_ssbox_address40;
reg    cipher_0_ssbox_ce40;
wire   [7:0] cipher_0_ssbox_q40;
wire   [7:0] cipher_0_ssbox_address41;
reg    cipher_0_ssbox_ce41;
wire   [7:0] cipher_0_ssbox_q41;
wire   [7:0] cipher_0_ssbox_address42;
reg    cipher_0_ssbox_ce42;
wire   [7:0] cipher_0_ssbox_q42;
wire   [7:0] cipher_0_ssbox_address43;
reg    cipher_0_ssbox_ce43;
wire   [7:0] cipher_0_ssbox_q43;
wire   [7:0] cipher_0_ssbox_address44;
reg    cipher_0_ssbox_ce44;
wire   [7:0] cipher_0_ssbox_q44;
wire   [7:0] cipher_0_ssbox_address45;
reg    cipher_0_ssbox_ce45;
wire   [7:0] cipher_0_ssbox_q45;
wire   [7:0] cipher_0_ssbox_address46;
reg    cipher_0_ssbox_ce46;
wire   [7:0] cipher_0_ssbox_q46;
wire   [7:0] cipher_0_ssbox_address47;
reg    cipher_0_ssbox_ce47;
wire   [7:0] cipher_0_ssbox_q47;
wire   [7:0] cipher_0_ssbox_address48;
reg    cipher_0_ssbox_ce48;
wire   [7:0] cipher_0_ssbox_q48;
wire   [7:0] cipher_0_ssbox_address49;
reg    cipher_0_ssbox_ce49;
wire   [7:0] cipher_0_ssbox_q49;
wire   [7:0] cipher_0_ssbox_address50;
reg    cipher_0_ssbox_ce50;
wire   [7:0] cipher_0_ssbox_q50;
wire   [7:0] cipher_0_ssbox_address51;
reg    cipher_0_ssbox_ce51;
wire   [7:0] cipher_0_ssbox_q51;
wire   [7:0] cipher_0_ssbox_address52;
reg    cipher_0_ssbox_ce52;
wire   [7:0] cipher_0_ssbox_q52;
wire   [7:0] cipher_0_ssbox_address53;
reg    cipher_0_ssbox_ce53;
wire   [7:0] cipher_0_ssbox_q53;
wire   [7:0] cipher_0_ssbox_address54;
reg    cipher_0_ssbox_ce54;
wire   [7:0] cipher_0_ssbox_q54;
wire   [7:0] cipher_0_ssbox_address55;
reg    cipher_0_ssbox_ce55;
wire   [7:0] cipher_0_ssbox_q55;
wire   [7:0] cipher_0_ssbox_address56;
reg    cipher_0_ssbox_ce56;
wire   [7:0] cipher_0_ssbox_q56;
wire   [7:0] cipher_0_ssbox_address57;
reg    cipher_0_ssbox_ce57;
wire   [7:0] cipher_0_ssbox_q57;
wire   [7:0] cipher_0_ssbox_address58;
reg    cipher_0_ssbox_ce58;
wire   [7:0] cipher_0_ssbox_q58;
wire   [7:0] cipher_0_ssbox_address59;
reg    cipher_0_ssbox_ce59;
wire   [7:0] cipher_0_ssbox_q59;
wire   [7:0] cipher_0_ssbox_address60;
reg    cipher_0_ssbox_ce60;
wire   [7:0] cipher_0_ssbox_q60;
wire   [7:0] cipher_0_ssbox_address61;
reg    cipher_0_ssbox_ce61;
wire   [7:0] cipher_0_ssbox_q61;
wire   [7:0] cipher_0_ssbox_address62;
reg    cipher_0_ssbox_ce62;
wire   [7:0] cipher_0_ssbox_q62;
wire   [7:0] cipher_0_ssbox_address63;
reg    cipher_0_ssbox_ce63;
wire   [7:0] cipher_0_ssbox_q63;
wire   [7:0] cipher_0_ssbox_address64;
reg    cipher_0_ssbox_ce64;
wire   [7:0] cipher_0_ssbox_q64;
wire   [7:0] cipher_0_ssbox_address65;
reg    cipher_0_ssbox_ce65;
wire   [7:0] cipher_0_ssbox_q65;
wire   [7:0] cipher_0_ssbox_address66;
reg    cipher_0_ssbox_ce66;
wire   [7:0] cipher_0_ssbox_q66;
wire   [7:0] cipher_0_ssbox_address67;
reg    cipher_0_ssbox_ce67;
wire   [7:0] cipher_0_ssbox_q67;
wire   [7:0] cipher_0_ssbox_address68;
reg    cipher_0_ssbox_ce68;
wire   [7:0] cipher_0_ssbox_q68;
wire   [7:0] cipher_0_ssbox_address69;
reg    cipher_0_ssbox_ce69;
wire   [7:0] cipher_0_ssbox_q69;
wire   [7:0] cipher_0_ssbox_address70;
reg    cipher_0_ssbox_ce70;
wire   [7:0] cipher_0_ssbox_q70;
wire   [7:0] cipher_0_ssbox_address71;
reg    cipher_0_ssbox_ce71;
wire   [7:0] cipher_0_ssbox_q71;
wire   [7:0] cipher_0_ssbox_address72;
reg    cipher_0_ssbox_ce72;
wire   [7:0] cipher_0_ssbox_q72;
wire   [7:0] cipher_0_ssbox_address73;
reg    cipher_0_ssbox_ce73;
wire   [7:0] cipher_0_ssbox_q73;
wire   [7:0] cipher_0_ssbox_address74;
reg    cipher_0_ssbox_ce74;
wire   [7:0] cipher_0_ssbox_q74;
wire   [7:0] cipher_0_ssbox_address75;
reg    cipher_0_ssbox_ce75;
wire   [7:0] cipher_0_ssbox_q75;
wire   [7:0] cipher_0_ssbox_address76;
reg    cipher_0_ssbox_ce76;
wire   [7:0] cipher_0_ssbox_q76;
wire   [7:0] cipher_0_ssbox_address77;
reg    cipher_0_ssbox_ce77;
wire   [7:0] cipher_0_ssbox_q77;
wire   [7:0] cipher_0_ssbox_address78;
reg    cipher_0_ssbox_ce78;
wire   [7:0] cipher_0_ssbox_q78;
wire   [7:0] cipher_0_ssbox_address79;
reg    cipher_0_ssbox_ce79;
wire   [7:0] cipher_0_ssbox_q79;
wire   [7:0] cipher_0_ssbox_address80;
reg    cipher_0_ssbox_ce80;
wire   [7:0] cipher_0_ssbox_q80;
wire   [7:0] cipher_0_ssbox_address81;
reg    cipher_0_ssbox_ce81;
wire   [7:0] cipher_0_ssbox_q81;
wire   [7:0] cipher_0_ssbox_address82;
reg    cipher_0_ssbox_ce82;
wire   [7:0] cipher_0_ssbox_q82;
wire   [7:0] cipher_0_ssbox_address83;
reg    cipher_0_ssbox_ce83;
wire   [7:0] cipher_0_ssbox_q83;
wire   [7:0] cipher_0_ssbox_address84;
reg    cipher_0_ssbox_ce84;
wire   [7:0] cipher_0_ssbox_q84;
wire   [7:0] cipher_0_ssbox_address85;
reg    cipher_0_ssbox_ce85;
wire   [7:0] cipher_0_ssbox_q85;
wire   [7:0] cipher_0_ssbox_address86;
reg    cipher_0_ssbox_ce86;
wire   [7:0] cipher_0_ssbox_q86;
wire   [7:0] cipher_0_ssbox_address87;
reg    cipher_0_ssbox_ce87;
wire   [7:0] cipher_0_ssbox_q87;
wire   [7:0] cipher_0_ssbox_address88;
reg    cipher_0_ssbox_ce88;
wire   [7:0] cipher_0_ssbox_q88;
wire   [7:0] cipher_0_ssbox_address89;
reg    cipher_0_ssbox_ce89;
wire   [7:0] cipher_0_ssbox_q89;
wire   [7:0] cipher_0_ssbox_address90;
reg    cipher_0_ssbox_ce90;
wire   [7:0] cipher_0_ssbox_q90;
wire   [7:0] cipher_0_ssbox_address91;
reg    cipher_0_ssbox_ce91;
wire   [7:0] cipher_0_ssbox_q91;
wire   [7:0] cipher_0_ssbox_address92;
reg    cipher_0_ssbox_ce92;
wire   [7:0] cipher_0_ssbox_q92;
wire   [7:0] cipher_0_ssbox_address93;
reg    cipher_0_ssbox_ce93;
wire   [7:0] cipher_0_ssbox_q93;
wire   [7:0] cipher_0_ssbox_address94;
reg    cipher_0_ssbox_ce94;
wire   [7:0] cipher_0_ssbox_q94;
wire   [7:0] cipher_0_ssbox_address95;
reg    cipher_0_ssbox_ce95;
wire   [7:0] cipher_0_ssbox_q95;
wire   [7:0] cipher_0_ssbox_address96;
reg    cipher_0_ssbox_ce96;
wire   [7:0] cipher_0_ssbox_q96;
wire   [7:0] cipher_0_ssbox_address97;
reg    cipher_0_ssbox_ce97;
wire   [7:0] cipher_0_ssbox_q97;
wire   [7:0] cipher_0_ssbox_address98;
reg    cipher_0_ssbox_ce98;
wire   [7:0] cipher_0_ssbox_q98;
wire   [7:0] cipher_0_ssbox_address99;
reg    cipher_0_ssbox_ce99;
wire   [7:0] cipher_0_ssbox_q99;
wire   [7:0] cipher_0_ssbox_address100;
reg    cipher_0_ssbox_ce100;
wire   [7:0] cipher_0_ssbox_q100;
wire   [7:0] cipher_0_ssbox_address101;
reg    cipher_0_ssbox_ce101;
wire   [7:0] cipher_0_ssbox_q101;
wire   [7:0] cipher_0_ssbox_address102;
reg    cipher_0_ssbox_ce102;
wire   [7:0] cipher_0_ssbox_q102;
wire   [7:0] cipher_0_ssbox_address103;
reg    cipher_0_ssbox_ce103;
wire   [7:0] cipher_0_ssbox_q103;
wire   [7:0] cipher_0_ssbox_address104;
reg    cipher_0_ssbox_ce104;
wire   [7:0] cipher_0_ssbox_q104;
wire   [7:0] cipher_0_ssbox_address105;
reg    cipher_0_ssbox_ce105;
wire   [7:0] cipher_0_ssbox_q105;
wire   [7:0] cipher_0_ssbox_address106;
reg    cipher_0_ssbox_ce106;
wire   [7:0] cipher_0_ssbox_q106;
wire   [7:0] cipher_0_ssbox_address107;
reg    cipher_0_ssbox_ce107;
wire   [7:0] cipher_0_ssbox_q107;
wire   [7:0] cipher_0_ssbox_address108;
reg    cipher_0_ssbox_ce108;
wire   [7:0] cipher_0_ssbox_q108;
wire   [7:0] cipher_0_ssbox_address109;
reg    cipher_0_ssbox_ce109;
wire   [7:0] cipher_0_ssbox_q109;
wire   [7:0] cipher_0_ssbox_address110;
reg    cipher_0_ssbox_ce110;
wire   [7:0] cipher_0_ssbox_q110;
wire   [7:0] cipher_0_ssbox_address111;
reg    cipher_0_ssbox_ce111;
wire   [7:0] cipher_0_ssbox_q111;
wire   [7:0] cipher_0_ssbox_address112;
reg    cipher_0_ssbox_ce112;
wire   [7:0] cipher_0_ssbox_q112;
wire   [7:0] cipher_0_ssbox_address113;
reg    cipher_0_ssbox_ce113;
wire   [7:0] cipher_0_ssbox_q113;
wire   [7:0] cipher_0_ssbox_address114;
reg    cipher_0_ssbox_ce114;
wire   [7:0] cipher_0_ssbox_q114;
wire   [7:0] cipher_0_ssbox_address115;
reg    cipher_0_ssbox_ce115;
wire   [7:0] cipher_0_ssbox_q115;
wire   [7:0] cipher_0_ssbox_address116;
reg    cipher_0_ssbox_ce116;
wire   [7:0] cipher_0_ssbox_q116;
wire   [7:0] cipher_0_ssbox_address117;
reg    cipher_0_ssbox_ce117;
wire   [7:0] cipher_0_ssbox_q117;
wire   [7:0] cipher_0_ssbox_address118;
reg    cipher_0_ssbox_ce118;
wire   [7:0] cipher_0_ssbox_q118;
wire   [7:0] cipher_0_ssbox_address119;
reg    cipher_0_ssbox_ce119;
wire   [7:0] cipher_0_ssbox_q119;
wire   [7:0] cipher_0_ssbox_address120;
reg    cipher_0_ssbox_ce120;
wire   [7:0] cipher_0_ssbox_q120;
wire   [7:0] cipher_0_ssbox_address121;
reg    cipher_0_ssbox_ce121;
wire   [7:0] cipher_0_ssbox_q121;
wire   [7:0] cipher_0_ssbox_address122;
reg    cipher_0_ssbox_ce122;
wire   [7:0] cipher_0_ssbox_q122;
wire   [7:0] cipher_0_ssbox_address123;
reg    cipher_0_ssbox_ce123;
wire   [7:0] cipher_0_ssbox_q123;
wire   [7:0] cipher_0_ssbox_address124;
reg    cipher_0_ssbox_ce124;
wire   [7:0] cipher_0_ssbox_q124;
wire   [7:0] cipher_0_ssbox_address125;
reg    cipher_0_ssbox_ce125;
wire   [7:0] cipher_0_ssbox_q125;
wire   [7:0] cipher_0_ssbox_address126;
reg    cipher_0_ssbox_ce126;
wire   [7:0] cipher_0_ssbox_q126;
wire   [7:0] cipher_0_ssbox_address127;
reg    cipher_0_ssbox_ce127;
wire   [7:0] cipher_0_ssbox_q127;
wire   [7:0] cipher_0_ssbox_address128;
reg    cipher_0_ssbox_ce128;
wire   [7:0] cipher_0_ssbox_q128;
wire   [7:0] cipher_0_ssbox_address129;
reg    cipher_0_ssbox_ce129;
wire   [7:0] cipher_0_ssbox_q129;
wire   [7:0] cipher_0_ssbox_address130;
reg    cipher_0_ssbox_ce130;
wire   [7:0] cipher_0_ssbox_q130;
wire   [7:0] cipher_0_ssbox_address131;
reg    cipher_0_ssbox_ce131;
wire   [7:0] cipher_0_ssbox_q131;
wire   [7:0] cipher_0_ssbox_address132;
reg    cipher_0_ssbox_ce132;
wire   [7:0] cipher_0_ssbox_q132;
wire   [7:0] cipher_0_ssbox_address133;
reg    cipher_0_ssbox_ce133;
wire   [7:0] cipher_0_ssbox_q133;
wire   [7:0] cipher_0_ssbox_address134;
reg    cipher_0_ssbox_ce134;
wire   [7:0] cipher_0_ssbox_q134;
wire   [7:0] cipher_0_ssbox_address135;
reg    cipher_0_ssbox_ce135;
wire   [7:0] cipher_0_ssbox_q135;
wire   [7:0] cipher_0_ssbox_address136;
reg    cipher_0_ssbox_ce136;
wire   [7:0] cipher_0_ssbox_q136;
wire   [7:0] cipher_0_ssbox_address137;
reg    cipher_0_ssbox_ce137;
wire   [7:0] cipher_0_ssbox_q137;
wire   [7:0] cipher_0_ssbox_address138;
reg    cipher_0_ssbox_ce138;
wire   [7:0] cipher_0_ssbox_q138;
wire   [7:0] cipher_0_ssbox_address139;
reg    cipher_0_ssbox_ce139;
wire   [7:0] cipher_0_ssbox_q139;
wire   [7:0] cipher_0_ssbox_address140;
reg    cipher_0_ssbox_ce140;
wire   [7:0] cipher_0_ssbox_q140;
wire   [7:0] cipher_0_ssbox_address141;
reg    cipher_0_ssbox_ce141;
wire   [7:0] cipher_0_ssbox_q141;
wire   [7:0] cipher_0_ssbox_address142;
reg    cipher_0_ssbox_ce142;
wire   [7:0] cipher_0_ssbox_q142;
wire   [7:0] cipher_0_ssbox_address143;
reg    cipher_0_ssbox_ce143;
wire   [7:0] cipher_0_ssbox_q143;
wire   [7:0] cipher_0_ssbox_address144;
reg    cipher_0_ssbox_ce144;
wire   [7:0] cipher_0_ssbox_q144;
wire   [7:0] cipher_0_ssbox_address145;
reg    cipher_0_ssbox_ce145;
wire   [7:0] cipher_0_ssbox_q145;
wire   [7:0] cipher_0_ssbox_address146;
reg    cipher_0_ssbox_ce146;
wire   [7:0] cipher_0_ssbox_q146;
wire   [7:0] cipher_0_ssbox_address147;
reg    cipher_0_ssbox_ce147;
wire   [7:0] cipher_0_ssbox_q147;
wire   [7:0] cipher_0_ssbox_address148;
reg    cipher_0_ssbox_ce148;
wire   [7:0] cipher_0_ssbox_q148;
wire   [7:0] cipher_0_ssbox_address149;
reg    cipher_0_ssbox_ce149;
wire   [7:0] cipher_0_ssbox_q149;
wire   [7:0] cipher_0_ssbox_address150;
reg    cipher_0_ssbox_ce150;
wire   [7:0] cipher_0_ssbox_q150;
wire   [7:0] cipher_0_ssbox_address151;
reg    cipher_0_ssbox_ce151;
wire   [7:0] cipher_0_ssbox_q151;
wire   [7:0] cipher_0_ssbox_address152;
reg    cipher_0_ssbox_ce152;
wire   [7:0] cipher_0_ssbox_q152;
wire   [7:0] cipher_0_ssbox_address153;
reg    cipher_0_ssbox_ce153;
wire   [7:0] cipher_0_ssbox_q153;
wire   [7:0] cipher_0_ssbox_address154;
reg    cipher_0_ssbox_ce154;
wire   [7:0] cipher_0_ssbox_q154;
wire   [7:0] cipher_0_ssbox_address155;
reg    cipher_0_ssbox_ce155;
wire   [7:0] cipher_0_ssbox_q155;
wire   [7:0] cipher_0_ssbox_address156;
reg    cipher_0_ssbox_ce156;
wire   [7:0] cipher_0_ssbox_q156;
wire   [7:0] cipher_0_ssbox_address157;
reg    cipher_0_ssbox_ce157;
wire   [7:0] cipher_0_ssbox_q157;
wire   [7:0] cipher_0_ssbox_address158;
reg    cipher_0_ssbox_ce158;
wire   [7:0] cipher_0_ssbox_q158;
wire   [7:0] cipher_0_ssbox_address159;
reg    cipher_0_ssbox_ce159;
wire   [7:0] cipher_0_ssbox_q159;
wire   [7:0] cipher_0_p16box_address0;
reg    cipher_0_p16box_ce0;
wire   [15:0] cipher_0_p16box_q0;
wire   [7:0] cipher_0_p16box_address1;
reg    cipher_0_p16box_ce1;
wire   [15:0] cipher_0_p16box_q1;
wire   [7:0] cipher_0_p16box_address2;
reg    cipher_0_p16box_ce2;
wire   [15:0] cipher_0_p16box_q2;
wire   [7:0] cipher_0_p16box_address3;
reg    cipher_0_p16box_ce3;
wire   [15:0] cipher_0_p16box_q3;
wire   [7:0] cipher_0_p16box_address4;
reg    cipher_0_p16box_ce4;
wire   [15:0] cipher_0_p16box_q4;
wire   [7:0] cipher_0_p16box_address5;
reg    cipher_0_p16box_ce5;
wire   [15:0] cipher_0_p16box_q5;
wire   [7:0] cipher_0_p16box_address6;
reg    cipher_0_p16box_ce6;
wire   [15:0] cipher_0_p16box_q6;
wire   [7:0] cipher_0_p16box_address7;
reg    cipher_0_p16box_ce7;
wire   [15:0] cipher_0_p16box_q7;
wire   [7:0] cipher_0_p16box_address8;
reg    cipher_0_p16box_ce8;
wire   [15:0] cipher_0_p16box_q8;
wire   [7:0] cipher_0_p16box_address9;
reg    cipher_0_p16box_ce9;
wire   [15:0] cipher_0_p16box_q9;
wire   [7:0] cipher_0_p16box_address10;
reg    cipher_0_p16box_ce10;
wire   [15:0] cipher_0_p16box_q10;
wire   [7:0] cipher_0_p16box_address11;
reg    cipher_0_p16box_ce11;
wire   [15:0] cipher_0_p16box_q11;
wire   [7:0] cipher_0_p16box_address12;
reg    cipher_0_p16box_ce12;
wire   [15:0] cipher_0_p16box_q12;
wire   [7:0] cipher_0_p16box_address13;
reg    cipher_0_p16box_ce13;
wire   [15:0] cipher_0_p16box_q13;
wire   [7:0] cipher_0_p16box_address14;
reg    cipher_0_p16box_ce14;
wire   [15:0] cipher_0_p16box_q14;
wire   [7:0] cipher_0_p16box_address15;
reg    cipher_0_p16box_ce15;
wire   [15:0] cipher_0_p16box_q15;
wire   [7:0] cipher_0_p16box_address16;
reg    cipher_0_p16box_ce16;
wire   [15:0] cipher_0_p16box_q16;
wire   [7:0] cipher_0_p16box_address17;
reg    cipher_0_p16box_ce17;
wire   [15:0] cipher_0_p16box_q17;
wire   [7:0] cipher_0_p16box_address18;
reg    cipher_0_p16box_ce18;
wire   [15:0] cipher_0_p16box_q18;
wire   [7:0] cipher_0_p16box_address19;
reg    cipher_0_p16box_ce19;
wire   [15:0] cipher_0_p16box_q19;
wire   [7:0] cipher_0_p16box_address20;
reg    cipher_0_p16box_ce20;
wire   [15:0] cipher_0_p16box_q20;
wire   [7:0] cipher_0_p16box_address21;
reg    cipher_0_p16box_ce21;
wire   [15:0] cipher_0_p16box_q21;
wire   [7:0] cipher_0_p16box_address22;
reg    cipher_0_p16box_ce22;
wire   [15:0] cipher_0_p16box_q22;
wire   [7:0] cipher_0_p16box_address23;
reg    cipher_0_p16box_ce23;
wire   [15:0] cipher_0_p16box_q23;
wire   [7:0] cipher_0_p16box_address24;
reg    cipher_0_p16box_ce24;
wire   [15:0] cipher_0_p16box_q24;
wire   [7:0] cipher_0_p16box_address25;
reg    cipher_0_p16box_ce25;
wire   [15:0] cipher_0_p16box_q25;
wire   [7:0] cipher_0_p16box_address26;
reg    cipher_0_p16box_ce26;
wire   [15:0] cipher_0_p16box_q26;
wire   [7:0] cipher_0_p16box_address27;
reg    cipher_0_p16box_ce27;
wire   [15:0] cipher_0_p16box_q27;
wire   [7:0] cipher_0_p16box_address28;
reg    cipher_0_p16box_ce28;
wire   [15:0] cipher_0_p16box_q28;
wire   [7:0] cipher_0_p16box_address29;
reg    cipher_0_p16box_ce29;
wire   [15:0] cipher_0_p16box_q29;
wire   [7:0] cipher_0_p16box_address30;
reg    cipher_0_p16box_ce30;
wire   [15:0] cipher_0_p16box_q30;
wire   [7:0] cipher_0_p16box_address31;
reg    cipher_0_p16box_ce31;
wire   [15:0] cipher_0_p16box_q31;
wire   [7:0] cipher_0_p16box_address32;
reg    cipher_0_p16box_ce32;
wire   [15:0] cipher_0_p16box_q32;
wire   [7:0] cipher_0_p16box_address33;
reg    cipher_0_p16box_ce33;
wire   [15:0] cipher_0_p16box_q33;
wire   [7:0] cipher_0_p16box_address34;
reg    cipher_0_p16box_ce34;
wire   [15:0] cipher_0_p16box_q34;
wire   [7:0] cipher_0_p16box_address35;
reg    cipher_0_p16box_ce35;
wire   [15:0] cipher_0_p16box_q35;
wire   [7:0] cipher_0_p16box_address36;
reg    cipher_0_p16box_ce36;
wire   [15:0] cipher_0_p16box_q36;
wire   [7:0] cipher_0_p16box_address37;
reg    cipher_0_p16box_ce37;
wire   [15:0] cipher_0_p16box_q37;
wire   [7:0] cipher_0_p16box_address38;
reg    cipher_0_p16box_ce38;
wire   [15:0] cipher_0_p16box_q38;
wire   [7:0] cipher_0_p16box_address39;
reg    cipher_0_p16box_ce39;
wire   [15:0] cipher_0_p16box_q39;
wire   [7:0] cipher_0_p16box_address40;
reg    cipher_0_p16box_ce40;
wire   [15:0] cipher_0_p16box_q40;
wire   [7:0] cipher_0_p16box_address41;
reg    cipher_0_p16box_ce41;
wire   [15:0] cipher_0_p16box_q41;
wire   [7:0] cipher_0_p16box_address42;
reg    cipher_0_p16box_ce42;
wire   [15:0] cipher_0_p16box_q42;
wire   [7:0] cipher_0_p16box_address43;
reg    cipher_0_p16box_ce43;
wire   [15:0] cipher_0_p16box_q43;
wire   [7:0] cipher_0_p16box_address44;
reg    cipher_0_p16box_ce44;
wire   [15:0] cipher_0_p16box_q44;
wire   [7:0] cipher_0_p16box_address45;
reg    cipher_0_p16box_ce45;
wire   [15:0] cipher_0_p16box_q45;
wire   [7:0] cipher_0_p16box_address46;
reg    cipher_0_p16box_ce46;
wire   [15:0] cipher_0_p16box_q46;
wire   [7:0] cipher_0_p16box_address47;
reg    cipher_0_p16box_ce47;
wire   [15:0] cipher_0_p16box_q47;
wire   [7:0] cipher_0_p16box_address48;
reg    cipher_0_p16box_ce48;
wire   [15:0] cipher_0_p16box_q48;
wire   [7:0] cipher_0_p16box_address49;
reg    cipher_0_p16box_ce49;
wire   [15:0] cipher_0_p16box_q49;
wire   [7:0] cipher_0_p16box_address50;
reg    cipher_0_p16box_ce50;
wire   [15:0] cipher_0_p16box_q50;
wire   [7:0] cipher_0_p16box_address51;
reg    cipher_0_p16box_ce51;
wire   [15:0] cipher_0_p16box_q51;
wire   [7:0] cipher_0_p16box_address52;
reg    cipher_0_p16box_ce52;
wire   [15:0] cipher_0_p16box_q52;
wire   [7:0] cipher_0_p16box_address53;
reg    cipher_0_p16box_ce53;
wire   [15:0] cipher_0_p16box_q53;
wire   [7:0] cipher_0_p16box_address54;
reg    cipher_0_p16box_ce54;
wire   [15:0] cipher_0_p16box_q54;
wire   [7:0] cipher_0_p16box_address55;
reg    cipher_0_p16box_ce55;
wire   [15:0] cipher_0_p16box_q55;
wire   [7:0] cipher_0_p16box_address56;
reg    cipher_0_p16box_ce56;
wire   [15:0] cipher_0_p16box_q56;
wire   [7:0] cipher_0_p16box_address57;
reg    cipher_0_p16box_ce57;
wire   [15:0] cipher_0_p16box_q57;
wire   [7:0] cipher_0_p16box_address58;
reg    cipher_0_p16box_ce58;
wire   [15:0] cipher_0_p16box_q58;
wire   [7:0] cipher_0_p16box_address59;
reg    cipher_0_p16box_ce59;
wire   [15:0] cipher_0_p16box_q59;
wire   [7:0] cipher_0_p16box_address60;
reg    cipher_0_p16box_ce60;
wire   [15:0] cipher_0_p16box_q60;
wire   [7:0] cipher_0_p16box_address61;
reg    cipher_0_p16box_ce61;
wire   [15:0] cipher_0_p16box_q61;
wire   [7:0] cipher_0_p16box_address62;
reg    cipher_0_p16box_ce62;
wire   [15:0] cipher_0_p16box_q62;
wire   [7:0] cipher_0_p16box_address63;
reg    cipher_0_p16box_ce63;
wire   [15:0] cipher_0_p16box_q63;
wire   [7:0] cipher_0_p16box_address64;
reg    cipher_0_p16box_ce64;
wire   [15:0] cipher_0_p16box_q64;
wire   [7:0] cipher_0_p16box_address65;
reg    cipher_0_p16box_ce65;
wire   [15:0] cipher_0_p16box_q65;
wire   [7:0] cipher_0_p16box_address66;
reg    cipher_0_p16box_ce66;
wire   [15:0] cipher_0_p16box_q66;
wire   [7:0] cipher_0_p16box_address67;
reg    cipher_0_p16box_ce67;
wire   [15:0] cipher_0_p16box_q67;
wire   [7:0] cipher_0_p16box_address68;
reg    cipher_0_p16box_ce68;
wire   [15:0] cipher_0_p16box_q68;
wire   [7:0] cipher_0_p16box_address69;
reg    cipher_0_p16box_ce69;
wire   [15:0] cipher_0_p16box_q69;
wire   [7:0] cipher_0_p16box_address70;
reg    cipher_0_p16box_ce70;
wire   [15:0] cipher_0_p16box_q70;
wire   [7:0] cipher_0_p16box_address71;
reg    cipher_0_p16box_ce71;
wire   [15:0] cipher_0_p16box_q71;
wire   [7:0] cipher_0_p16box_address72;
reg    cipher_0_p16box_ce72;
wire   [15:0] cipher_0_p16box_q72;
wire   [7:0] cipher_0_p16box_address73;
reg    cipher_0_p16box_ce73;
wire   [15:0] cipher_0_p16box_q73;
wire   [7:0] cipher_0_p16box_address74;
reg    cipher_0_p16box_ce74;
wire   [15:0] cipher_0_p16box_q74;
wire   [7:0] cipher_0_p16box_address75;
reg    cipher_0_p16box_ce75;
wire   [15:0] cipher_0_p16box_q75;
wire   [7:0] cipher_0_p16box_address76;
reg    cipher_0_p16box_ce76;
wire   [15:0] cipher_0_p16box_q76;
wire   [7:0] cipher_0_p16box_address77;
reg    cipher_0_p16box_ce77;
wire   [15:0] cipher_0_p16box_q77;
wire   [7:0] cipher_0_p16box_address78;
reg    cipher_0_p16box_ce78;
wire   [15:0] cipher_0_p16box_q78;
wire   [7:0] cipher_0_p16box_address79;
reg    cipher_0_p16box_ce79;
wire   [15:0] cipher_0_p16box_q79;
wire   [7:0] cipher_0_p16box_address80;
reg    cipher_0_p16box_ce80;
wire   [15:0] cipher_0_p16box_q80;
wire   [7:0] cipher_0_p16box_address81;
reg    cipher_0_p16box_ce81;
wire   [15:0] cipher_0_p16box_q81;
wire   [7:0] cipher_0_p16box_address82;
reg    cipher_0_p16box_ce82;
wire   [15:0] cipher_0_p16box_q82;
wire   [7:0] cipher_0_p16box_address83;
reg    cipher_0_p16box_ce83;
wire   [15:0] cipher_0_p16box_q83;
wire   [7:0] cipher_0_p16box_address84;
reg    cipher_0_p16box_ce84;
wire   [15:0] cipher_0_p16box_q84;
wire   [7:0] cipher_0_p16box_address85;
reg    cipher_0_p16box_ce85;
wire   [15:0] cipher_0_p16box_q85;
wire   [7:0] cipher_0_p16box_address86;
reg    cipher_0_p16box_ce86;
wire   [15:0] cipher_0_p16box_q86;
wire   [7:0] cipher_0_p16box_address87;
reg    cipher_0_p16box_ce87;
wire   [15:0] cipher_0_p16box_q87;
wire   [7:0] cipher_0_p16box_address88;
reg    cipher_0_p16box_ce88;
wire   [15:0] cipher_0_p16box_q88;
wire   [7:0] cipher_0_p16box_address89;
reg    cipher_0_p16box_ce89;
wire   [15:0] cipher_0_p16box_q89;
wire   [7:0] cipher_0_p16box_address90;
reg    cipher_0_p16box_ce90;
wire   [15:0] cipher_0_p16box_q90;
wire   [7:0] cipher_0_p16box_address91;
reg    cipher_0_p16box_ce91;
wire   [15:0] cipher_0_p16box_q91;
wire   [7:0] cipher_0_p16box_address92;
reg    cipher_0_p16box_ce92;
wire   [15:0] cipher_0_p16box_q92;
wire   [7:0] cipher_0_p16box_address93;
reg    cipher_0_p16box_ce93;
wire   [15:0] cipher_0_p16box_q93;
wire   [7:0] cipher_0_p16box_address94;
reg    cipher_0_p16box_ce94;
wire   [15:0] cipher_0_p16box_q94;
wire   [7:0] cipher_0_p16box_address95;
reg    cipher_0_p16box_ce95;
wire   [15:0] cipher_0_p16box_q95;
wire   [7:0] cipher_0_p16box_address96;
reg    cipher_0_p16box_ce96;
wire   [15:0] cipher_0_p16box_q96;
wire   [7:0] cipher_0_p16box_address97;
reg    cipher_0_p16box_ce97;
wire   [15:0] cipher_0_p16box_q97;
wire   [7:0] cipher_0_p16box_address98;
reg    cipher_0_p16box_ce98;
wire   [15:0] cipher_0_p16box_q98;
wire   [7:0] cipher_0_p16box_address99;
reg    cipher_0_p16box_ce99;
wire   [15:0] cipher_0_p16box_q99;
wire   [7:0] cipher_0_p16box_address100;
reg    cipher_0_p16box_ce100;
wire   [15:0] cipher_0_p16box_q100;
wire   [7:0] cipher_0_p16box_address101;
reg    cipher_0_p16box_ce101;
wire   [15:0] cipher_0_p16box_q101;
wire   [7:0] cipher_0_p16box_address102;
reg    cipher_0_p16box_ce102;
wire   [15:0] cipher_0_p16box_q102;
wire   [7:0] cipher_0_p16box_address103;
reg    cipher_0_p16box_ce103;
wire   [15:0] cipher_0_p16box_q103;
wire   [7:0] cipher_0_p16box_address104;
reg    cipher_0_p16box_ce104;
wire   [15:0] cipher_0_p16box_q104;
wire   [7:0] cipher_0_p16box_address105;
reg    cipher_0_p16box_ce105;
wire   [15:0] cipher_0_p16box_q105;
wire   [7:0] cipher_0_p16box_address106;
reg    cipher_0_p16box_ce106;
wire   [15:0] cipher_0_p16box_q106;
wire   [7:0] cipher_0_p16box_address107;
reg    cipher_0_p16box_ce107;
wire   [15:0] cipher_0_p16box_q107;
wire   [7:0] cipher_0_p16box_address108;
reg    cipher_0_p16box_ce108;
wire   [15:0] cipher_0_p16box_q108;
wire   [7:0] cipher_0_p16box_address109;
reg    cipher_0_p16box_ce109;
wire   [15:0] cipher_0_p16box_q109;
wire   [7:0] cipher_0_p16box_address110;
reg    cipher_0_p16box_ce110;
wire   [15:0] cipher_0_p16box_q110;
wire   [7:0] cipher_0_p16box_address111;
reg    cipher_0_p16box_ce111;
wire   [15:0] cipher_0_p16box_q111;
wire   [7:0] cipher_0_p16box_address112;
reg    cipher_0_p16box_ce112;
wire   [15:0] cipher_0_p16box_q112;
wire   [7:0] cipher_0_p16box_address113;
reg    cipher_0_p16box_ce113;
wire   [15:0] cipher_0_p16box_q113;
wire   [7:0] cipher_0_p16box_address114;
reg    cipher_0_p16box_ce114;
wire   [15:0] cipher_0_p16box_q114;
wire   [7:0] cipher_0_p16box_address115;
reg    cipher_0_p16box_ce115;
wire   [15:0] cipher_0_p16box_q115;
wire   [7:0] cipher_0_p16box_address116;
reg    cipher_0_p16box_ce116;
wire   [15:0] cipher_0_p16box_q116;
wire   [7:0] cipher_0_p16box_address117;
reg    cipher_0_p16box_ce117;
wire   [15:0] cipher_0_p16box_q117;
wire   [7:0] cipher_0_p16box_address118;
reg    cipher_0_p16box_ce118;
wire   [15:0] cipher_0_p16box_q118;
wire   [7:0] cipher_0_p16box_address119;
reg    cipher_0_p16box_ce119;
wire   [15:0] cipher_0_p16box_q119;
wire   [7:0] cipher_0_p16box_address120;
reg    cipher_0_p16box_ce120;
wire   [15:0] cipher_0_p16box_q120;
wire   [7:0] cipher_0_p16box_address121;
reg    cipher_0_p16box_ce121;
wire   [15:0] cipher_0_p16box_q121;
wire   [7:0] cipher_0_p16box_address122;
reg    cipher_0_p16box_ce122;
wire   [15:0] cipher_0_p16box_q122;
wire   [7:0] cipher_0_p16box_address123;
reg    cipher_0_p16box_ce123;
wire   [15:0] cipher_0_p16box_q123;
wire   [7:0] cipher_0_p16box_address124;
reg    cipher_0_p16box_ce124;
wire   [15:0] cipher_0_p16box_q124;
wire   [7:0] cipher_0_p16box_address125;
reg    cipher_0_p16box_ce125;
wire   [15:0] cipher_0_p16box_q125;
wire   [7:0] cipher_0_p16box_address126;
reg    cipher_0_p16box_ce126;
wire   [15:0] cipher_0_p16box_q126;
wire   [7:0] cipher_0_p16box_address127;
reg    cipher_0_p16box_ce127;
wire   [15:0] cipher_0_p16box_q127;
wire   [7:0] cipher_0_p16box_address128;
reg    cipher_0_p16box_ce128;
wire   [15:0] cipher_0_p16box_q128;
wire   [7:0] cipher_0_p16box_address129;
reg    cipher_0_p16box_ce129;
wire   [15:0] cipher_0_p16box_q129;
wire   [7:0] cipher_0_p16box_address130;
reg    cipher_0_p16box_ce130;
wire   [15:0] cipher_0_p16box_q130;
wire   [7:0] cipher_0_p16box_address131;
reg    cipher_0_p16box_ce131;
wire   [15:0] cipher_0_p16box_q131;
wire   [7:0] cipher_0_p16box_address132;
reg    cipher_0_p16box_ce132;
wire   [15:0] cipher_0_p16box_q132;
wire   [7:0] cipher_0_p16box_address133;
reg    cipher_0_p16box_ce133;
wire   [15:0] cipher_0_p16box_q133;
wire   [7:0] cipher_0_p16box_address134;
reg    cipher_0_p16box_ce134;
wire   [15:0] cipher_0_p16box_q134;
wire   [7:0] cipher_0_p16box_address135;
reg    cipher_0_p16box_ce135;
wire   [15:0] cipher_0_p16box_q135;
wire   [7:0] cipher_0_p16box_address136;
reg    cipher_0_p16box_ce136;
wire   [15:0] cipher_0_p16box_q136;
wire   [7:0] cipher_0_p16box_address137;
reg    cipher_0_p16box_ce137;
wire   [15:0] cipher_0_p16box_q137;
wire   [7:0] cipher_0_p16box_address138;
reg    cipher_0_p16box_ce138;
wire   [15:0] cipher_0_p16box_q138;
wire   [7:0] cipher_0_p16box_address139;
reg    cipher_0_p16box_ce139;
wire   [15:0] cipher_0_p16box_q139;
wire   [7:0] cipher_0_p16box_address140;
reg    cipher_0_p16box_ce140;
wire   [15:0] cipher_0_p16box_q140;
wire   [7:0] cipher_0_p16box_address141;
reg    cipher_0_p16box_ce141;
wire   [15:0] cipher_0_p16box_q141;
wire   [7:0] cipher_0_p16box_address142;
reg    cipher_0_p16box_ce142;
wire   [15:0] cipher_0_p16box_q142;
wire   [7:0] cipher_0_p16box_address143;
reg    cipher_0_p16box_ce143;
wire   [15:0] cipher_0_p16box_q143;
reg   [127:0] p_read_1_reg_11624;
wire    ap_block_pp0_stage0_11001;
reg   [127:0] p_read_1_reg_11624_pp0_iter1_reg;
reg   [127:0] p_read_1_reg_11624_pp0_iter2_reg;
reg   [127:0] p_read_1_reg_11624_pp0_iter3_reg;
reg   [127:0] p_read_1_reg_11624_pp0_iter4_reg;
reg   [127:0] p_read_1_reg_11624_pp0_iter5_reg;
reg   [127:0] p_read_1_reg_11624_pp0_iter6_reg;
reg   [127:0] p_read_1_reg_11624_pp0_iter7_reg;
reg   [127:0] p_read_1_reg_11624_pp0_iter8_reg;
reg   [127:0] p_read_1_reg_11624_pp0_iter9_reg;
reg   [127:0] p_read_1_reg_11624_pp0_iter10_reg;
reg   [127:0] p_read_1_reg_11624_pp0_iter11_reg;
reg   [127:0] p_read_1_reg_11624_pp0_iter12_reg;
reg   [127:0] p_read_1_reg_11624_pp0_iter13_reg;
reg   [127:0] p_read_1_reg_11624_pp0_iter14_reg;
reg   [127:0] p_read_1_reg_11624_pp0_iter15_reg;
reg   [127:0] p_read_1_reg_11624_pp0_iter16_reg;
reg   [127:0] p_read_1_reg_11624_pp0_iter17_reg;
reg   [127:0] p_read_1_reg_11624_pp0_iter18_reg;
reg   [127:0] p_read_2_reg_11629;
reg   [127:0] p_read_2_reg_11629_pp0_iter1_reg;
reg   [127:0] p_read_2_reg_11629_pp0_iter2_reg;
reg   [127:0] p_read_2_reg_11629_pp0_iter3_reg;
reg   [127:0] p_read_2_reg_11629_pp0_iter4_reg;
reg   [127:0] p_read_2_reg_11629_pp0_iter5_reg;
reg   [127:0] p_read_2_reg_11629_pp0_iter6_reg;
reg   [127:0] p_read_2_reg_11629_pp0_iter7_reg;
reg   [127:0] p_read_2_reg_11629_pp0_iter8_reg;
reg   [127:0] p_read_2_reg_11629_pp0_iter9_reg;
reg   [127:0] p_read_2_reg_11629_pp0_iter10_reg;
reg   [127:0] p_read_2_reg_11629_pp0_iter11_reg;
reg   [127:0] p_read_2_reg_11629_pp0_iter12_reg;
reg   [127:0] p_read_2_reg_11629_pp0_iter13_reg;
reg   [127:0] p_read_2_reg_11629_pp0_iter14_reg;
reg   [127:0] p_read_2_reg_11629_pp0_iter15_reg;
reg   [127:0] p_read_2_reg_11629_pp0_iter16_reg;
reg   [127:0] p_read_2_reg_11629_pp0_iter17_reg;
reg   [127:0] p_read_3_reg_11634;
reg   [127:0] p_read_3_reg_11634_pp0_iter1_reg;
reg   [127:0] p_read_3_reg_11634_pp0_iter2_reg;
reg   [127:0] p_read_3_reg_11634_pp0_iter3_reg;
reg   [127:0] p_read_3_reg_11634_pp0_iter4_reg;
reg   [127:0] p_read_3_reg_11634_pp0_iter5_reg;
reg   [127:0] p_read_3_reg_11634_pp0_iter6_reg;
reg   [127:0] p_read_3_reg_11634_pp0_iter7_reg;
reg   [127:0] p_read_3_reg_11634_pp0_iter8_reg;
reg   [127:0] p_read_3_reg_11634_pp0_iter9_reg;
reg   [127:0] p_read_3_reg_11634_pp0_iter10_reg;
reg   [127:0] p_read_3_reg_11634_pp0_iter11_reg;
reg   [127:0] p_read_3_reg_11634_pp0_iter12_reg;
reg   [127:0] p_read_3_reg_11634_pp0_iter13_reg;
reg   [127:0] p_read_3_reg_11634_pp0_iter14_reg;
reg   [127:0] p_read_3_reg_11634_pp0_iter15_reg;
reg   [127:0] p_read_4_reg_11639;
reg   [127:0] p_read_4_reg_11639_pp0_iter1_reg;
reg   [127:0] p_read_4_reg_11639_pp0_iter2_reg;
reg   [127:0] p_read_4_reg_11639_pp0_iter3_reg;
reg   [127:0] p_read_4_reg_11639_pp0_iter4_reg;
reg   [127:0] p_read_4_reg_11639_pp0_iter5_reg;
reg   [127:0] p_read_4_reg_11639_pp0_iter6_reg;
reg   [127:0] p_read_4_reg_11639_pp0_iter7_reg;
reg   [127:0] p_read_4_reg_11639_pp0_iter8_reg;
reg   [127:0] p_read_4_reg_11639_pp0_iter9_reg;
reg   [127:0] p_read_4_reg_11639_pp0_iter10_reg;
reg   [127:0] p_read_4_reg_11639_pp0_iter11_reg;
reg   [127:0] p_read_4_reg_11639_pp0_iter12_reg;
reg   [127:0] p_read_4_reg_11639_pp0_iter13_reg;
reg   [127:0] p_read_5_reg_11644;
reg   [127:0] p_read_5_reg_11644_pp0_iter1_reg;
reg   [127:0] p_read_5_reg_11644_pp0_iter2_reg;
reg   [127:0] p_read_5_reg_11644_pp0_iter3_reg;
reg   [127:0] p_read_5_reg_11644_pp0_iter4_reg;
reg   [127:0] p_read_5_reg_11644_pp0_iter5_reg;
reg   [127:0] p_read_5_reg_11644_pp0_iter6_reg;
reg   [127:0] p_read_5_reg_11644_pp0_iter7_reg;
reg   [127:0] p_read_5_reg_11644_pp0_iter8_reg;
reg   [127:0] p_read_5_reg_11644_pp0_iter9_reg;
reg   [127:0] p_read_5_reg_11644_pp0_iter10_reg;
reg   [127:0] p_read_5_reg_11644_pp0_iter11_reg;
reg   [127:0] p_read_6_reg_11649;
reg   [127:0] p_read_6_reg_11649_pp0_iter1_reg;
reg   [127:0] p_read_6_reg_11649_pp0_iter2_reg;
reg   [127:0] p_read_6_reg_11649_pp0_iter3_reg;
reg   [127:0] p_read_6_reg_11649_pp0_iter4_reg;
reg   [127:0] p_read_6_reg_11649_pp0_iter5_reg;
reg   [127:0] p_read_6_reg_11649_pp0_iter6_reg;
reg   [127:0] p_read_6_reg_11649_pp0_iter7_reg;
reg   [127:0] p_read_6_reg_11649_pp0_iter8_reg;
reg   [127:0] p_read_6_reg_11649_pp0_iter9_reg;
reg   [127:0] p_read_7_reg_11654;
reg   [127:0] p_read_7_reg_11654_pp0_iter1_reg;
reg   [127:0] p_read_7_reg_11654_pp0_iter2_reg;
reg   [127:0] p_read_7_reg_11654_pp0_iter3_reg;
reg   [127:0] p_read_7_reg_11654_pp0_iter4_reg;
reg   [127:0] p_read_7_reg_11654_pp0_iter5_reg;
reg   [127:0] p_read_7_reg_11654_pp0_iter6_reg;
reg   [127:0] p_read_7_reg_11654_pp0_iter7_reg;
reg   [127:0] p_read_8_reg_11659;
reg   [127:0] p_read_8_reg_11659_pp0_iter1_reg;
reg   [127:0] p_read_8_reg_11659_pp0_iter2_reg;
reg   [127:0] p_read_8_reg_11659_pp0_iter3_reg;
reg   [127:0] p_read_8_reg_11659_pp0_iter4_reg;
reg   [127:0] p_read_8_reg_11659_pp0_iter5_reg;
reg   [127:0] p_read_9_reg_11664;
reg   [127:0] p_read_9_reg_11664_pp0_iter1_reg;
reg   [127:0] p_read_9_reg_11664_pp0_iter2_reg;
reg   [127:0] p_read_9_reg_11664_pp0_iter3_reg;
reg   [127:0] p_read_10_reg_11669;
reg   [127:0] p_read_10_reg_11669_pp0_iter1_reg;
reg   [7:0] tmp_V_reg_11754;
reg   [7:0] tmp_1_V_10_reg_11760;
reg   [7:0] tmp_2_1_V_10_reg_11766;
reg   [7:0] tmp_V_7_reg_11772;
reg   [7:0] tmp_V_4_reg_11778;
reg   [7:0] tmp_V_1_reg_11784;
reg   [7:0] tmp_2_2_V_10_reg_11790;
reg   [7:0] tmp_V_11_reg_11796;
reg   [7:0] tmp_V_8_reg_11802;
reg   [7:0] tmp_V_5_reg_11808;
reg   [7:0] tmp_V_2_reg_11814;
reg   [7:0] tmp_V_15_reg_11820;
reg   [7:0] tmp_V_12_reg_11826;
reg   [7:0] tmp_V_9_reg_11832;
reg   [7:0] tmp_V_6_reg_11838;
reg   [7:0] tmp_3_V_10_reg_11844;
reg   [7:0] tmp_V_16_reg_12010;
reg   [7:0] tmp_1_V_11_reg_12016;
reg   [7:0] tmp_2_1_V_11_reg_12022;
reg   [7:0] tmp_V_23_reg_12028;
reg   [7:0] tmp_V_20_reg_12034;
reg   [7:0] tmp_V_17_reg_12040;
reg   [7:0] tmp_2_2_V_11_reg_12046;
reg   [7:0] tmp_V_27_reg_12052;
reg   [7:0] tmp_V_24_reg_12058;
reg   [7:0] tmp_V_21_reg_12064;
reg   [7:0] tmp_V_18_reg_12070;
reg   [7:0] tmp_V_31_reg_12076;
reg   [7:0] tmp_V_28_reg_12082;
reg   [7:0] tmp_V_25_reg_12088;
reg   [7:0] tmp_V_22_reg_12094;
reg   [7:0] tmp_3_V_11_reg_12100;
reg   [7:0] tmp_V_32_reg_12266;
reg   [7:0] tmp_1_V_12_reg_12272;
reg   [7:0] tmp_2_1_V_12_reg_12278;
reg   [7:0] tmp_V_39_reg_12284;
reg   [7:0] tmp_V_36_reg_12290;
reg   [7:0] tmp_V_33_reg_12296;
reg   [7:0] tmp_2_2_V_12_reg_12302;
reg   [7:0] tmp_V_43_reg_12308;
reg   [7:0] tmp_V_40_reg_12314;
reg   [7:0] tmp_V_37_reg_12320;
reg   [7:0] tmp_V_34_reg_12326;
reg   [7:0] tmp_V_47_reg_12332;
reg   [7:0] tmp_V_44_reg_12338;
reg   [7:0] tmp_V_41_reg_12344;
reg   [7:0] tmp_V_38_reg_12350;
reg   [7:0] tmp_3_V_12_reg_12356;
reg   [7:0] tmp_V_48_reg_12522;
reg   [7:0] tmp_1_V_13_reg_12528;
reg   [7:0] tmp_2_1_V_13_reg_12534;
reg   [7:0] tmp_V_55_reg_12540;
reg   [7:0] tmp_V_52_reg_12546;
reg   [7:0] tmp_V_49_reg_12552;
reg   [7:0] tmp_2_2_V_13_reg_12558;
reg   [7:0] tmp_V_59_reg_12564;
reg   [7:0] tmp_V_56_reg_12570;
reg   [7:0] tmp_V_53_reg_12576;
reg   [7:0] tmp_V_50_reg_12582;
reg   [7:0] tmp_V_63_reg_12588;
reg   [7:0] tmp_V_60_reg_12594;
reg   [7:0] tmp_V_57_reg_12600;
reg   [7:0] tmp_V_54_reg_12606;
reg   [7:0] tmp_3_V_13_reg_12612;
reg   [7:0] tmp_V_64_reg_12778;
reg   [7:0] tmp_1_V_14_reg_12784;
reg   [7:0] tmp_2_1_V_14_reg_12790;
reg   [7:0] tmp_V_71_reg_12796;
reg   [7:0] tmp_V_68_reg_12802;
reg   [7:0] tmp_V_65_reg_12808;
reg   [7:0] tmp_2_2_V_14_reg_12814;
reg   [7:0] tmp_V_75_reg_12820;
reg   [7:0] tmp_V_72_reg_12826;
reg   [7:0] tmp_V_69_reg_12832;
reg   [7:0] tmp_V_66_reg_12838;
reg   [7:0] tmp_V_79_reg_12844;
reg   [7:0] tmp_V_76_reg_12850;
reg   [7:0] tmp_V_73_reg_12856;
reg   [7:0] tmp_V_70_reg_12862;
reg   [7:0] tmp_3_V_14_reg_12868;
reg   [7:0] tmp_V_80_reg_13034;
reg   [7:0] tmp_1_V_15_reg_13040;
reg   [7:0] tmp_2_1_V_15_reg_13046;
reg   [7:0] tmp_V_87_reg_13052;
reg   [7:0] tmp_V_84_reg_13058;
reg   [7:0] tmp_V_81_reg_13064;
reg   [7:0] tmp_2_2_V_15_reg_13070;
reg   [7:0] tmp_V_91_reg_13076;
reg   [7:0] tmp_V_88_reg_13082;
reg   [7:0] tmp_V_85_reg_13088;
reg   [7:0] tmp_V_82_reg_13094;
reg   [7:0] tmp_V_95_reg_13100;
reg   [7:0] tmp_V_92_reg_13106;
reg   [7:0] tmp_V_89_reg_13112;
reg   [7:0] tmp_V_86_reg_13118;
reg   [7:0] tmp_3_V_15_reg_13124;
reg   [7:0] tmp_V_96_reg_13290;
reg   [7:0] tmp_1_V_16_reg_13296;
reg   [7:0] tmp_2_1_V_16_reg_13302;
reg   [7:0] tmp_V_103_reg_13308;
reg   [7:0] tmp_V_100_reg_13314;
reg   [7:0] tmp_V_97_reg_13320;
reg   [7:0] tmp_2_2_V_16_reg_13326;
reg   [7:0] tmp_V_107_reg_13332;
reg   [7:0] tmp_V_104_reg_13338;
reg   [7:0] tmp_V_101_reg_13344;
reg   [7:0] tmp_V_98_reg_13350;
reg   [7:0] tmp_V_111_reg_13356;
reg   [7:0] tmp_V_108_reg_13362;
reg   [7:0] tmp_V_105_reg_13368;
reg   [7:0] tmp_V_102_reg_13374;
reg   [7:0] tmp_3_V_16_reg_13380;
reg   [7:0] tmp_V_112_reg_13546;
reg   [7:0] tmp_1_V_17_reg_13552;
reg   [7:0] tmp_2_1_V_17_reg_13558;
reg   [7:0] tmp_V_119_reg_13564;
reg   [7:0] tmp_V_116_reg_13570;
reg   [7:0] tmp_V_113_reg_13576;
reg   [7:0] tmp_2_2_V_17_reg_13582;
reg   [7:0] tmp_V_123_reg_13588;
reg   [7:0] tmp_V_120_reg_13594;
reg   [7:0] tmp_V_117_reg_13600;
reg   [7:0] tmp_V_114_reg_13606;
reg   [7:0] tmp_V_127_reg_13612;
reg   [7:0] tmp_V_124_reg_13618;
reg   [7:0] tmp_V_121_reg_13624;
reg   [7:0] tmp_V_118_reg_13630;
reg   [7:0] tmp_3_V_17_reg_13636;
reg   [7:0] tmp_V_128_reg_13802;
reg   [7:0] tmp_1_V_18_reg_13808;
reg   [7:0] tmp_2_1_V_18_reg_13814;
reg   [7:0] tmp_V_135_reg_13820;
reg   [7:0] tmp_V_132_reg_13826;
reg   [7:0] tmp_V_129_reg_13832;
reg   [7:0] tmp_2_2_V_18_reg_13838;
reg   [7:0] tmp_V_139_reg_13844;
reg   [7:0] tmp_V_136_reg_13850;
reg   [7:0] tmp_V_133_reg_13856;
reg   [7:0] tmp_V_130_reg_13862;
reg   [7:0] tmp_V_143_reg_13868;
reg   [7:0] tmp_V_140_reg_13874;
reg   [7:0] tmp_V_137_reg_13880;
reg   [7:0] tmp_V_134_reg_13886;
reg   [7:0] tmp_3_V_18_reg_13892;
wire   [63:0] zext_ln708_fu_3838_p1;
wire    ap_block_pp0_stage0;
wire   [63:0] zext_ln708_4_fu_3853_p1;
wire   [63:0] zext_ln708_5_fu_3868_p1;
wire   [63:0] zext_ln708_6_fu_3883_p1;
wire   [63:0] zext_ln708_7_fu_3898_p1;
wire   [63:0] zext_ln708_8_fu_3913_p1;
wire   [63:0] zext_ln708_9_fu_3928_p1;
wire   [63:0] zext_ln708_10_fu_3943_p1;
wire   [63:0] zext_ln708_11_fu_3958_p1;
wire   [63:0] zext_ln708_12_fu_3973_p1;
wire   [63:0] zext_ln708_13_fu_3988_p1;
wire   [63:0] zext_ln708_14_fu_4003_p1;
wire   [63:0] zext_ln708_15_fu_4018_p1;
wire   [63:0] zext_ln708_16_fu_4033_p1;
wire   [63:0] zext_ln708_17_fu_4048_p1;
wire   [63:0] zext_ln708_18_fu_4063_p1;
wire   [63:0] zext_ln587_fu_4068_p1;
wire   [63:0] zext_ln587_1_fu_4073_p1;
wire   [63:0] zext_ln587_2_fu_4078_p1;
wire   [63:0] zext_ln587_3_fu_4083_p1;
wire   [63:0] zext_ln587_4_fu_4088_p1;
wire   [63:0] zext_ln587_5_fu_4093_p1;
wire   [63:0] zext_ln587_6_fu_4098_p1;
wire   [63:0] zext_ln587_7_fu_4103_p1;
wire   [63:0] zext_ln587_8_fu_4108_p1;
wire   [63:0] zext_ln587_9_fu_4113_p1;
wire   [63:0] zext_ln587_10_fu_4118_p1;
wire   [63:0] zext_ln587_11_fu_4123_p1;
wire   [63:0] zext_ln587_12_fu_4128_p1;
wire   [63:0] zext_ln587_13_fu_4133_p1;
wire   [63:0] zext_ln587_14_fu_4138_p1;
wire   [63:0] zext_ln587_15_fu_4143_p1;
wire   [63:0] zext_ln708_19_fu_4673_p1;
wire   [63:0] zext_ln708_20_fu_4688_p1;
wire   [63:0] zext_ln708_21_fu_4703_p1;
wire   [63:0] zext_ln708_22_fu_4718_p1;
wire   [63:0] zext_ln708_23_fu_4733_p1;
wire   [63:0] zext_ln708_24_fu_4748_p1;
wire   [63:0] zext_ln708_25_fu_4763_p1;
wire   [63:0] zext_ln708_26_fu_4778_p1;
wire   [63:0] zext_ln708_27_fu_4793_p1;
wire   [63:0] zext_ln708_28_fu_4808_p1;
wire   [63:0] zext_ln708_29_fu_4823_p1;
wire   [63:0] zext_ln708_30_fu_4838_p1;
wire   [63:0] zext_ln708_31_fu_4853_p1;
wire   [63:0] zext_ln708_32_fu_4868_p1;
wire   [63:0] zext_ln708_33_fu_4883_p1;
wire   [63:0] zext_ln708_34_fu_4898_p1;
wire   [63:0] zext_ln587_16_fu_4903_p1;
wire   [63:0] zext_ln587_17_fu_4908_p1;
wire   [63:0] zext_ln587_18_fu_4913_p1;
wire   [63:0] zext_ln587_19_fu_4918_p1;
wire   [63:0] zext_ln587_20_fu_4923_p1;
wire   [63:0] zext_ln587_21_fu_4928_p1;
wire   [63:0] zext_ln587_22_fu_4933_p1;
wire   [63:0] zext_ln587_23_fu_4938_p1;
wire   [63:0] zext_ln587_24_fu_4943_p1;
wire   [63:0] zext_ln587_25_fu_4948_p1;
wire   [63:0] zext_ln587_26_fu_4953_p1;
wire   [63:0] zext_ln587_27_fu_4958_p1;
wire   [63:0] zext_ln587_28_fu_4963_p1;
wire   [63:0] zext_ln587_29_fu_4968_p1;
wire   [63:0] zext_ln587_30_fu_4973_p1;
wire   [63:0] zext_ln587_31_fu_4978_p1;
wire   [63:0] zext_ln708_35_fu_5508_p1;
wire   [63:0] zext_ln708_36_fu_5523_p1;
wire   [63:0] zext_ln708_37_fu_5538_p1;
wire   [63:0] zext_ln708_38_fu_5553_p1;
wire   [63:0] zext_ln708_39_fu_5568_p1;
wire   [63:0] zext_ln708_40_fu_5583_p1;
wire   [63:0] zext_ln708_41_fu_5598_p1;
wire   [63:0] zext_ln708_42_fu_5613_p1;
wire   [63:0] zext_ln708_43_fu_5628_p1;
wire   [63:0] zext_ln708_44_fu_5643_p1;
wire   [63:0] zext_ln708_45_fu_5658_p1;
wire   [63:0] zext_ln708_46_fu_5673_p1;
wire   [63:0] zext_ln708_47_fu_5688_p1;
wire   [63:0] zext_ln708_48_fu_5703_p1;
wire   [63:0] zext_ln708_49_fu_5718_p1;
wire   [63:0] zext_ln708_50_fu_5733_p1;
wire   [63:0] zext_ln587_32_fu_5738_p1;
wire   [63:0] zext_ln587_33_fu_5743_p1;
wire   [63:0] zext_ln587_34_fu_5748_p1;
wire   [63:0] zext_ln587_35_fu_5753_p1;
wire   [63:0] zext_ln587_36_fu_5758_p1;
wire   [63:0] zext_ln587_37_fu_5763_p1;
wire   [63:0] zext_ln587_38_fu_5768_p1;
wire   [63:0] zext_ln587_39_fu_5773_p1;
wire   [63:0] zext_ln587_40_fu_5778_p1;
wire   [63:0] zext_ln587_41_fu_5783_p1;
wire   [63:0] zext_ln587_42_fu_5788_p1;
wire   [63:0] zext_ln587_43_fu_5793_p1;
wire   [63:0] zext_ln587_44_fu_5798_p1;
wire   [63:0] zext_ln587_45_fu_5803_p1;
wire   [63:0] zext_ln587_46_fu_5808_p1;
wire   [63:0] zext_ln587_47_fu_5813_p1;
wire   [63:0] zext_ln708_51_fu_6343_p1;
wire   [63:0] zext_ln708_52_fu_6358_p1;
wire   [63:0] zext_ln708_53_fu_6373_p1;
wire   [63:0] zext_ln708_54_fu_6388_p1;
wire   [63:0] zext_ln708_55_fu_6403_p1;
wire   [63:0] zext_ln708_56_fu_6418_p1;
wire   [63:0] zext_ln708_57_fu_6433_p1;
wire   [63:0] zext_ln708_58_fu_6448_p1;
wire   [63:0] zext_ln708_59_fu_6463_p1;
wire   [63:0] zext_ln708_60_fu_6478_p1;
wire   [63:0] zext_ln708_61_fu_6493_p1;
wire   [63:0] zext_ln708_62_fu_6508_p1;
wire   [63:0] zext_ln708_63_fu_6523_p1;
wire   [63:0] zext_ln708_64_fu_6538_p1;
wire   [63:0] zext_ln708_65_fu_6553_p1;
wire   [63:0] zext_ln708_66_fu_6568_p1;
wire   [63:0] zext_ln587_48_fu_6573_p1;
wire   [63:0] zext_ln587_49_fu_6578_p1;
wire   [63:0] zext_ln587_50_fu_6583_p1;
wire   [63:0] zext_ln587_51_fu_6588_p1;
wire   [63:0] zext_ln587_52_fu_6593_p1;
wire   [63:0] zext_ln587_53_fu_6598_p1;
wire   [63:0] zext_ln587_54_fu_6603_p1;
wire   [63:0] zext_ln587_55_fu_6608_p1;
wire   [63:0] zext_ln587_56_fu_6613_p1;
wire   [63:0] zext_ln587_57_fu_6618_p1;
wire   [63:0] zext_ln587_58_fu_6623_p1;
wire   [63:0] zext_ln587_59_fu_6628_p1;
wire   [63:0] zext_ln587_60_fu_6633_p1;
wire   [63:0] zext_ln587_61_fu_6638_p1;
wire   [63:0] zext_ln587_62_fu_6643_p1;
wire   [63:0] zext_ln587_63_fu_6648_p1;
wire   [63:0] zext_ln708_67_fu_7178_p1;
wire   [63:0] zext_ln708_68_fu_7193_p1;
wire   [63:0] zext_ln708_69_fu_7208_p1;
wire   [63:0] zext_ln708_70_fu_7223_p1;
wire   [63:0] zext_ln708_71_fu_7238_p1;
wire   [63:0] zext_ln708_72_fu_7253_p1;
wire   [63:0] zext_ln708_73_fu_7268_p1;
wire   [63:0] zext_ln708_74_fu_7283_p1;
wire   [63:0] zext_ln708_75_fu_7298_p1;
wire   [63:0] zext_ln708_76_fu_7313_p1;
wire   [63:0] zext_ln708_77_fu_7328_p1;
wire   [63:0] zext_ln708_78_fu_7343_p1;
wire   [63:0] zext_ln708_79_fu_7358_p1;
wire   [63:0] zext_ln708_80_fu_7373_p1;
wire   [63:0] zext_ln708_81_fu_7388_p1;
wire   [63:0] zext_ln708_82_fu_7403_p1;
wire   [63:0] zext_ln587_64_fu_7408_p1;
wire   [63:0] zext_ln587_65_fu_7413_p1;
wire   [63:0] zext_ln587_66_fu_7418_p1;
wire   [63:0] zext_ln587_67_fu_7423_p1;
wire   [63:0] zext_ln587_68_fu_7428_p1;
wire   [63:0] zext_ln587_69_fu_7433_p1;
wire   [63:0] zext_ln587_70_fu_7438_p1;
wire   [63:0] zext_ln587_71_fu_7443_p1;
wire   [63:0] zext_ln587_72_fu_7448_p1;
wire   [63:0] zext_ln587_73_fu_7453_p1;
wire   [63:0] zext_ln587_74_fu_7458_p1;
wire   [63:0] zext_ln587_75_fu_7463_p1;
wire   [63:0] zext_ln587_76_fu_7468_p1;
wire   [63:0] zext_ln587_77_fu_7473_p1;
wire   [63:0] zext_ln587_78_fu_7478_p1;
wire   [63:0] zext_ln587_79_fu_7483_p1;
wire   [63:0] zext_ln708_83_fu_8013_p1;
wire   [63:0] zext_ln708_84_fu_8028_p1;
wire   [63:0] zext_ln708_85_fu_8043_p1;
wire   [63:0] zext_ln708_86_fu_8058_p1;
wire   [63:0] zext_ln708_87_fu_8073_p1;
wire   [63:0] zext_ln708_88_fu_8088_p1;
wire   [63:0] zext_ln708_89_fu_8103_p1;
wire   [63:0] zext_ln708_90_fu_8118_p1;
wire   [63:0] zext_ln708_91_fu_8133_p1;
wire   [63:0] zext_ln708_92_fu_8148_p1;
wire   [63:0] zext_ln708_93_fu_8163_p1;
wire   [63:0] zext_ln708_94_fu_8178_p1;
wire   [63:0] zext_ln708_95_fu_8193_p1;
wire   [63:0] zext_ln708_96_fu_8208_p1;
wire   [63:0] zext_ln708_97_fu_8223_p1;
wire   [63:0] zext_ln708_98_fu_8238_p1;
wire   [63:0] zext_ln587_80_fu_8243_p1;
wire   [63:0] zext_ln587_81_fu_8248_p1;
wire   [63:0] zext_ln587_82_fu_8253_p1;
wire   [63:0] zext_ln587_83_fu_8258_p1;
wire   [63:0] zext_ln587_84_fu_8263_p1;
wire   [63:0] zext_ln587_85_fu_8268_p1;
wire   [63:0] zext_ln587_86_fu_8273_p1;
wire   [63:0] zext_ln587_87_fu_8278_p1;
wire   [63:0] zext_ln587_88_fu_8283_p1;
wire   [63:0] zext_ln587_89_fu_8288_p1;
wire   [63:0] zext_ln587_90_fu_8293_p1;
wire   [63:0] zext_ln587_91_fu_8298_p1;
wire   [63:0] zext_ln587_92_fu_8303_p1;
wire   [63:0] zext_ln587_93_fu_8308_p1;
wire   [63:0] zext_ln587_94_fu_8313_p1;
wire   [63:0] zext_ln587_95_fu_8318_p1;
wire   [63:0] zext_ln708_99_fu_8848_p1;
wire   [63:0] zext_ln708_100_fu_8863_p1;
wire   [63:0] zext_ln708_101_fu_8878_p1;
wire   [63:0] zext_ln708_102_fu_8893_p1;
wire   [63:0] zext_ln708_103_fu_8908_p1;
wire   [63:0] zext_ln708_104_fu_8923_p1;
wire   [63:0] zext_ln708_105_fu_8938_p1;
wire   [63:0] zext_ln708_106_fu_8953_p1;
wire   [63:0] zext_ln708_107_fu_8968_p1;
wire   [63:0] zext_ln708_108_fu_8983_p1;
wire   [63:0] zext_ln708_109_fu_8998_p1;
wire   [63:0] zext_ln708_110_fu_9013_p1;
wire   [63:0] zext_ln708_111_fu_9028_p1;
wire   [63:0] zext_ln708_112_fu_9043_p1;
wire   [63:0] zext_ln708_113_fu_9058_p1;
wire   [63:0] zext_ln708_114_fu_9073_p1;
wire   [63:0] zext_ln587_96_fu_9078_p1;
wire   [63:0] zext_ln587_97_fu_9083_p1;
wire   [63:0] zext_ln587_98_fu_9088_p1;
wire   [63:0] zext_ln587_99_fu_9093_p1;
wire   [63:0] zext_ln587_100_fu_9098_p1;
wire   [63:0] zext_ln587_101_fu_9103_p1;
wire   [63:0] zext_ln587_102_fu_9108_p1;
wire   [63:0] zext_ln587_103_fu_9113_p1;
wire   [63:0] zext_ln587_104_fu_9118_p1;
wire   [63:0] zext_ln587_105_fu_9123_p1;
wire   [63:0] zext_ln587_106_fu_9128_p1;
wire   [63:0] zext_ln587_107_fu_9133_p1;
wire   [63:0] zext_ln587_108_fu_9138_p1;
wire   [63:0] zext_ln587_109_fu_9143_p1;
wire   [63:0] zext_ln587_110_fu_9148_p1;
wire   [63:0] zext_ln587_111_fu_9153_p1;
wire   [63:0] zext_ln708_115_fu_9683_p1;
wire   [63:0] zext_ln708_116_fu_9698_p1;
wire   [63:0] zext_ln708_117_fu_9713_p1;
wire   [63:0] zext_ln708_118_fu_9728_p1;
wire   [63:0] zext_ln708_119_fu_9743_p1;
wire   [63:0] zext_ln708_120_fu_9758_p1;
wire   [63:0] zext_ln708_121_fu_9773_p1;
wire   [63:0] zext_ln708_122_fu_9788_p1;
wire   [63:0] zext_ln708_123_fu_9803_p1;
wire   [63:0] zext_ln708_124_fu_9818_p1;
wire   [63:0] zext_ln708_125_fu_9833_p1;
wire   [63:0] zext_ln708_126_fu_9848_p1;
wire   [63:0] zext_ln708_127_fu_9863_p1;
wire   [63:0] zext_ln708_128_fu_9878_p1;
wire   [63:0] zext_ln708_129_fu_9893_p1;
wire   [63:0] zext_ln708_130_fu_9908_p1;
wire   [63:0] zext_ln587_112_fu_9913_p1;
wire   [63:0] zext_ln587_113_fu_9918_p1;
wire   [63:0] zext_ln587_114_fu_9923_p1;
wire   [63:0] zext_ln587_115_fu_9928_p1;
wire   [63:0] zext_ln587_116_fu_9933_p1;
wire   [63:0] zext_ln587_117_fu_9938_p1;
wire   [63:0] zext_ln587_118_fu_9943_p1;
wire   [63:0] zext_ln587_119_fu_9948_p1;
wire   [63:0] zext_ln587_120_fu_9953_p1;
wire   [63:0] zext_ln587_121_fu_9958_p1;
wire   [63:0] zext_ln587_122_fu_9963_p1;
wire   [63:0] zext_ln587_123_fu_9968_p1;
wire   [63:0] zext_ln587_124_fu_9973_p1;
wire   [63:0] zext_ln587_125_fu_9978_p1;
wire   [63:0] zext_ln587_126_fu_9983_p1;
wire   [63:0] zext_ln587_127_fu_9988_p1;
wire   [63:0] zext_ln708_131_fu_10518_p1;
wire   [63:0] zext_ln708_132_fu_10533_p1;
wire   [63:0] zext_ln708_133_fu_10548_p1;
wire   [63:0] zext_ln708_134_fu_10563_p1;
wire   [63:0] zext_ln708_135_fu_10578_p1;
wire   [63:0] zext_ln708_136_fu_10593_p1;
wire   [63:0] zext_ln708_137_fu_10608_p1;
wire   [63:0] zext_ln708_138_fu_10623_p1;
wire   [63:0] zext_ln708_139_fu_10638_p1;
wire   [63:0] zext_ln708_140_fu_10653_p1;
wire   [63:0] zext_ln708_141_fu_10668_p1;
wire   [63:0] zext_ln708_142_fu_10683_p1;
wire   [63:0] zext_ln708_143_fu_10698_p1;
wire   [63:0] zext_ln708_144_fu_10713_p1;
wire   [63:0] zext_ln708_145_fu_10728_p1;
wire   [63:0] zext_ln708_146_fu_10743_p1;
wire   [63:0] zext_ln587_128_fu_10748_p1;
wire   [63:0] zext_ln587_129_fu_10753_p1;
wire   [63:0] zext_ln587_130_fu_10758_p1;
wire   [63:0] zext_ln587_131_fu_10763_p1;
wire   [63:0] zext_ln587_132_fu_10768_p1;
wire   [63:0] zext_ln587_133_fu_10773_p1;
wire   [63:0] zext_ln587_134_fu_10778_p1;
wire   [63:0] zext_ln587_135_fu_10783_p1;
wire   [63:0] zext_ln587_136_fu_10788_p1;
wire   [63:0] zext_ln587_137_fu_10793_p1;
wire   [63:0] zext_ln587_138_fu_10798_p1;
wire   [63:0] zext_ln587_139_fu_10803_p1;
wire   [63:0] zext_ln587_140_fu_10808_p1;
wire   [63:0] zext_ln587_141_fu_10813_p1;
wire   [63:0] zext_ln587_142_fu_10818_p1;
wire   [63:0] zext_ln587_143_fu_10823_p1;
wire   [63:0] zext_ln708_147_fu_11353_p1;
wire   [63:0] zext_ln708_148_fu_11368_p1;
wire   [63:0] zext_ln708_149_fu_11383_p1;
wire   [63:0] zext_ln708_150_fu_11398_p1;
wire   [63:0] zext_ln708_151_fu_11413_p1;
wire   [63:0] zext_ln708_152_fu_11428_p1;
wire   [63:0] zext_ln708_153_fu_11443_p1;
wire   [63:0] zext_ln708_154_fu_11458_p1;
wire   [63:0] zext_ln708_155_fu_11473_p1;
wire   [63:0] zext_ln708_156_fu_11488_p1;
wire   [63:0] zext_ln708_157_fu_11503_p1;
wire   [63:0] zext_ln708_158_fu_11518_p1;
wire   [63:0] zext_ln708_159_fu_11533_p1;
wire   [63:0] zext_ln708_160_fu_11548_p1;
wire   [63:0] zext_ln708_161_fu_11563_p1;
wire   [63:0] zext_ln708_162_fu_11578_p1;
wire   [127:0] ret_V_fu_3828_p2;
wire   [7:0] trunc_ln708_fu_3834_p1;
wire   [7:0] tmp_s_fu_3843_p4;
wire   [7:0] tmp_4_fu_3858_p4;
wire   [7:0] tmp_5_fu_3873_p4;
wire   [7:0] tmp_6_fu_3888_p4;
wire   [7:0] tmp_7_fu_3903_p4;
wire   [7:0] tmp_8_fu_3918_p4;
wire   [7:0] tmp_9_fu_3933_p4;
wire   [7:0] tmp_10_fu_3948_p4;
wire   [7:0] tmp_11_fu_3963_p4;
wire   [7:0] tmp_12_fu_3978_p4;
wire   [7:0] tmp_13_fu_3993_p4;
wire   [7:0] tmp_14_fu_4008_p4;
wire   [7:0] tmp_15_fu_4023_p4;
wire   [7:0] tmp_16_fu_4038_p4;
wire   [7:0] tmp_17_fu_4053_p4;
wire   [7:0] tmp_19_fu_4166_p4;
wire   [7:0] trunc_ln674_fu_4148_p1;
wire   [7:0] xor_ln1545_6_fu_4376_p2;
wire   [7:0] xor_ln1545_fu_4372_p2;
wire   [7:0] trunc_ln674_1_fu_4162_p1;
wire   [7:0] tmp_20_fu_4180_p4;
wire   [7:0] xor_ln1545_9_fu_4392_p2;
wire   [7:0] xor_ln1545_7_fu_4388_p2;
wire   [7:0] trunc_ln674_2_fu_4176_p1;
wire   [7:0] tmp_21_fu_4194_p4;
wire   [7:0] xor_ln1545_12_fu_4408_p2;
wire   [7:0] xor_ln1545_10_fu_4404_p2;
wire   [7:0] tmp_18_fu_4152_p4;
wire   [7:0] trunc_ln674_3_fu_4190_p1;
wire   [7:0] xor_ln1545_15_fu_4424_p2;
wire   [7:0] xor_ln1545_13_fu_4420_p2;
wire   [7:0] tmp_23_fu_4222_p4;
wire   [7:0] trunc_ln674_4_fu_4204_p1;
wire   [7:0] xor_ln1545_18_fu_4440_p2;
wire   [7:0] xor_ln1545_16_fu_4436_p2;
wire   [7:0] trunc_ln674_5_fu_4218_p1;
wire   [7:0] tmp_24_fu_4236_p4;
wire   [7:0] xor_ln1545_21_fu_4456_p2;
wire   [7:0] xor_ln1545_19_fu_4452_p2;
wire   [7:0] trunc_ln674_6_fu_4232_p1;
wire   [7:0] tmp_25_fu_4250_p4;
wire   [7:0] xor_ln1545_24_fu_4472_p2;
wire   [7:0] xor_ln1545_22_fu_4468_p2;
wire   [7:0] tmp_22_fu_4208_p4;
wire   [7:0] trunc_ln674_7_fu_4246_p1;
wire   [7:0] xor_ln1545_27_fu_4488_p2;
wire   [7:0] xor_ln1545_25_fu_4484_p2;
wire   [7:0] tmp_27_fu_4278_p4;
wire   [7:0] trunc_ln674_8_fu_4260_p1;
wire   [7:0] xor_ln1545_30_fu_4504_p2;
wire   [7:0] xor_ln1545_28_fu_4500_p2;
wire   [7:0] trunc_ln674_9_fu_4274_p1;
wire   [7:0] tmp_28_fu_4292_p4;
wire   [7:0] xor_ln1545_33_fu_4520_p2;
wire   [7:0] xor_ln1545_31_fu_4516_p2;
wire   [7:0] trunc_ln674_10_fu_4288_p1;
wire   [7:0] tmp_29_fu_4306_p4;
wire   [7:0] xor_ln1545_36_fu_4536_p2;
wire   [7:0] xor_ln1545_34_fu_4532_p2;
wire   [7:0] tmp_26_fu_4264_p4;
wire   [7:0] trunc_ln674_11_fu_4302_p1;
wire   [7:0] xor_ln1545_39_fu_4552_p2;
wire   [7:0] xor_ln1545_37_fu_4548_p2;
wire   [7:0] tmp_31_fu_4334_p4;
wire   [7:0] trunc_ln674_12_fu_4316_p1;
wire   [7:0] xor_ln1545_42_fu_4568_p2;
wire   [7:0] xor_ln1545_40_fu_4564_p2;
wire   [7:0] trunc_ln674_13_fu_4330_p1;
wire   [7:0] tmp_32_fu_4348_p4;
wire   [7:0] xor_ln1545_45_fu_4584_p2;
wire   [7:0] xor_ln1545_43_fu_4580_p2;
wire   [7:0] trunc_ln674_14_fu_4344_p1;
wire   [7:0] tmp_33_fu_4362_p4;
wire   [7:0] xor_ln1545_48_fu_4600_p2;
wire   [7:0] xor_ln1545_46_fu_4596_p2;
wire   [7:0] tmp_30_fu_4320_p4;
wire   [7:0] trunc_ln674_15_fu_4358_p1;
wire   [7:0] xor_ln1545_51_fu_4616_p2;
wire   [7:0] xor_ln1545_49_fu_4612_p2;
wire   [7:0] xor_ln1545_50_fu_4622_p2;
wire   [7:0] xor_ln1545_47_fu_4606_p2;
wire   [7:0] xor_ln1545_44_fu_4590_p2;
wire   [7:0] xor_ln1545_41_fu_4574_p2;
wire   [7:0] xor_ln1545_38_fu_4558_p2;
wire   [7:0] xor_ln1545_35_fu_4542_p2;
wire   [7:0] xor_ln1545_32_fu_4526_p2;
wire   [7:0] xor_ln1545_29_fu_4510_p2;
wire   [7:0] xor_ln1545_26_fu_4494_p2;
wire   [7:0] xor_ln1545_23_fu_4478_p2;
wire   [7:0] xor_ln1545_20_fu_4462_p2;
wire   [7:0] xor_ln1545_17_fu_4446_p2;
wire   [7:0] xor_ln1545_14_fu_4430_p2;
wire   [7:0] xor_ln1545_11_fu_4414_p2;
wire   [7:0] xor_ln1545_8_fu_4398_p2;
wire   [7:0] xor_ln1545_5_fu_4382_p2;
wire   [127:0] p_Result_s_fu_4628_p17;
wire   [127:0] state_V_20_fu_4664_p2;
wire   [7:0] trunc_ln708_1_fu_4669_p1;
wire   [7:0] tmp_34_fu_4678_p4;
wire   [7:0] tmp_35_fu_4693_p4;
wire   [7:0] tmp_36_fu_4708_p4;
wire   [7:0] tmp_37_fu_4723_p4;
wire   [7:0] tmp_38_fu_4738_p4;
wire   [7:0] tmp_39_fu_4753_p4;
wire   [7:0] tmp_40_fu_4768_p4;
wire   [7:0] tmp_41_fu_4783_p4;
wire   [7:0] tmp_42_fu_4798_p4;
wire   [7:0] tmp_43_fu_4813_p4;
wire   [7:0] tmp_44_fu_4828_p4;
wire   [7:0] tmp_45_fu_4843_p4;
wire   [7:0] tmp_46_fu_4858_p4;
wire   [7:0] tmp_47_fu_4873_p4;
wire   [7:0] tmp_48_fu_4888_p4;
wire   [7:0] tmp_50_fu_5001_p4;
wire   [7:0] trunc_ln674_16_fu_4983_p1;
wire   [7:0] xor_ln1545_54_fu_5211_p2;
wire   [7:0] xor_ln1545_52_fu_5207_p2;
wire   [7:0] trunc_ln674_17_fu_4997_p1;
wire   [7:0] tmp_51_fu_5015_p4;
wire   [7:0] xor_ln1545_57_fu_5227_p2;
wire   [7:0] xor_ln1545_55_fu_5223_p2;
wire   [7:0] trunc_ln674_18_fu_5011_p1;
wire   [7:0] tmp_52_fu_5029_p4;
wire   [7:0] xor_ln1545_60_fu_5243_p2;
wire   [7:0] xor_ln1545_58_fu_5239_p2;
wire   [7:0] tmp_49_fu_4987_p4;
wire   [7:0] trunc_ln674_19_fu_5025_p1;
wire   [7:0] xor_ln1545_63_fu_5259_p2;
wire   [7:0] xor_ln1545_61_fu_5255_p2;
wire   [7:0] tmp_54_fu_5057_p4;
wire   [7:0] trunc_ln674_20_fu_5039_p1;
wire   [7:0] xor_ln1545_66_fu_5275_p2;
wire   [7:0] xor_ln1545_64_fu_5271_p2;
wire   [7:0] trunc_ln674_21_fu_5053_p1;
wire   [7:0] tmp_55_fu_5071_p4;
wire   [7:0] xor_ln1545_69_fu_5291_p2;
wire   [7:0] xor_ln1545_67_fu_5287_p2;
wire   [7:0] trunc_ln674_22_fu_5067_p1;
wire   [7:0] tmp_56_fu_5085_p4;
wire   [7:0] xor_ln1545_72_fu_5307_p2;
wire   [7:0] xor_ln1545_70_fu_5303_p2;
wire   [7:0] tmp_53_fu_5043_p4;
wire   [7:0] trunc_ln674_23_fu_5081_p1;
wire   [7:0] xor_ln1545_75_fu_5323_p2;
wire   [7:0] xor_ln1545_73_fu_5319_p2;
wire   [7:0] tmp_58_fu_5113_p4;
wire   [7:0] trunc_ln674_24_fu_5095_p1;
wire   [7:0] xor_ln1545_78_fu_5339_p2;
wire   [7:0] xor_ln1545_76_fu_5335_p2;
wire   [7:0] trunc_ln674_25_fu_5109_p1;
wire   [7:0] tmp_59_fu_5127_p4;
wire   [7:0] xor_ln1545_81_fu_5355_p2;
wire   [7:0] xor_ln1545_79_fu_5351_p2;
wire   [7:0] trunc_ln674_26_fu_5123_p1;
wire   [7:0] tmp_60_fu_5141_p4;
wire   [7:0] xor_ln1545_84_fu_5371_p2;
wire   [7:0] xor_ln1545_82_fu_5367_p2;
wire   [7:0] tmp_57_fu_5099_p4;
wire   [7:0] trunc_ln674_27_fu_5137_p1;
wire   [7:0] xor_ln1545_87_fu_5387_p2;
wire   [7:0] xor_ln1545_85_fu_5383_p2;
wire   [7:0] tmp_62_fu_5169_p4;
wire   [7:0] trunc_ln674_28_fu_5151_p1;
wire   [7:0] xor_ln1545_90_fu_5403_p2;
wire   [7:0] xor_ln1545_88_fu_5399_p2;
wire   [7:0] trunc_ln674_29_fu_5165_p1;
wire   [7:0] tmp_63_fu_5183_p4;
wire   [7:0] xor_ln1545_93_fu_5419_p2;
wire   [7:0] xor_ln1545_91_fu_5415_p2;
wire   [7:0] trunc_ln674_30_fu_5179_p1;
wire   [7:0] tmp_64_fu_5197_p4;
wire   [7:0] xor_ln1545_96_fu_5435_p2;
wire   [7:0] xor_ln1545_94_fu_5431_p2;
wire   [7:0] tmp_61_fu_5155_p4;
wire   [7:0] trunc_ln674_31_fu_5193_p1;
wire   [7:0] xor_ln1545_99_fu_5451_p2;
wire   [7:0] xor_ln1545_97_fu_5447_p2;
wire   [7:0] xor_ln1545_98_fu_5457_p2;
wire   [7:0] xor_ln1545_95_fu_5441_p2;
wire   [7:0] xor_ln1545_92_fu_5425_p2;
wire   [7:0] xor_ln1545_89_fu_5409_p2;
wire   [7:0] xor_ln1545_86_fu_5393_p2;
wire   [7:0] xor_ln1545_83_fu_5377_p2;
wire   [7:0] xor_ln1545_80_fu_5361_p2;
wire   [7:0] xor_ln1545_77_fu_5345_p2;
wire   [7:0] xor_ln1545_74_fu_5329_p2;
wire   [7:0] xor_ln1545_71_fu_5313_p2;
wire   [7:0] xor_ln1545_68_fu_5297_p2;
wire   [7:0] xor_ln1545_65_fu_5281_p2;
wire   [7:0] xor_ln1545_62_fu_5265_p2;
wire   [7:0] xor_ln1545_59_fu_5249_p2;
wire   [7:0] xor_ln1545_56_fu_5233_p2;
wire   [7:0] xor_ln1545_53_fu_5217_p2;
wire   [127:0] p_Result_2_fu_5463_p17;
wire   [127:0] state_V_21_fu_5499_p2;
wire   [7:0] trunc_ln708_2_fu_5504_p1;
wire   [7:0] tmp_65_fu_5513_p4;
wire   [7:0] tmp_66_fu_5528_p4;
wire   [7:0] tmp_67_fu_5543_p4;
wire   [7:0] tmp_68_fu_5558_p4;
wire   [7:0] tmp_69_fu_5573_p4;
wire   [7:0] tmp_70_fu_5588_p4;
wire   [7:0] tmp_71_fu_5603_p4;
wire   [7:0] tmp_72_fu_5618_p4;
wire   [7:0] tmp_73_fu_5633_p4;
wire   [7:0] tmp_74_fu_5648_p4;
wire   [7:0] tmp_75_fu_5663_p4;
wire   [7:0] tmp_76_fu_5678_p4;
wire   [7:0] tmp_77_fu_5693_p4;
wire   [7:0] tmp_78_fu_5708_p4;
wire   [7:0] tmp_79_fu_5723_p4;
wire   [7:0] tmp_81_fu_5836_p4;
wire   [7:0] trunc_ln674_32_fu_5818_p1;
wire   [7:0] xor_ln1545_102_fu_6046_p2;
wire   [7:0] xor_ln1545_100_fu_6042_p2;
wire   [7:0] trunc_ln674_33_fu_5832_p1;
wire   [7:0] tmp_82_fu_5850_p4;
wire   [7:0] xor_ln1545_105_fu_6062_p2;
wire   [7:0] xor_ln1545_103_fu_6058_p2;
wire   [7:0] trunc_ln674_34_fu_5846_p1;
wire   [7:0] tmp_83_fu_5864_p4;
wire   [7:0] xor_ln1545_108_fu_6078_p2;
wire   [7:0] xor_ln1545_106_fu_6074_p2;
wire   [7:0] tmp_80_fu_5822_p4;
wire   [7:0] trunc_ln674_35_fu_5860_p1;
wire   [7:0] xor_ln1545_111_fu_6094_p2;
wire   [7:0] xor_ln1545_109_fu_6090_p2;
wire   [7:0] tmp_85_fu_5892_p4;
wire   [7:0] trunc_ln674_36_fu_5874_p1;
wire   [7:0] xor_ln1545_114_fu_6110_p2;
wire   [7:0] xor_ln1545_112_fu_6106_p2;
wire   [7:0] trunc_ln674_37_fu_5888_p1;
wire   [7:0] tmp_86_fu_5906_p4;
wire   [7:0] xor_ln1545_117_fu_6126_p2;
wire   [7:0] xor_ln1545_115_fu_6122_p2;
wire   [7:0] trunc_ln674_38_fu_5902_p1;
wire   [7:0] tmp_87_fu_5920_p4;
wire   [7:0] xor_ln1545_120_fu_6142_p2;
wire   [7:0] xor_ln1545_118_fu_6138_p2;
wire   [7:0] tmp_84_fu_5878_p4;
wire   [7:0] trunc_ln674_39_fu_5916_p1;
wire   [7:0] xor_ln1545_123_fu_6158_p2;
wire   [7:0] xor_ln1545_121_fu_6154_p2;
wire   [7:0] tmp_89_fu_5948_p4;
wire   [7:0] trunc_ln674_40_fu_5930_p1;
wire   [7:0] xor_ln1545_126_fu_6174_p2;
wire   [7:0] xor_ln1545_124_fu_6170_p2;
wire   [7:0] trunc_ln674_41_fu_5944_p1;
wire   [7:0] tmp_90_fu_5962_p4;
wire   [7:0] xor_ln1545_129_fu_6190_p2;
wire   [7:0] xor_ln1545_127_fu_6186_p2;
wire   [7:0] trunc_ln674_42_fu_5958_p1;
wire   [7:0] tmp_91_fu_5976_p4;
wire   [7:0] xor_ln1545_132_fu_6206_p2;
wire   [7:0] xor_ln1545_130_fu_6202_p2;
wire   [7:0] tmp_88_fu_5934_p4;
wire   [7:0] trunc_ln674_43_fu_5972_p1;
wire   [7:0] xor_ln1545_135_fu_6222_p2;
wire   [7:0] xor_ln1545_133_fu_6218_p2;
wire   [7:0] tmp_93_fu_6004_p4;
wire   [7:0] trunc_ln674_44_fu_5986_p1;
wire   [7:0] xor_ln1545_138_fu_6238_p2;
wire   [7:0] xor_ln1545_136_fu_6234_p2;
wire   [7:0] trunc_ln674_45_fu_6000_p1;
wire   [7:0] tmp_94_fu_6018_p4;
wire   [7:0] xor_ln1545_141_fu_6254_p2;
wire   [7:0] xor_ln1545_139_fu_6250_p2;
wire   [7:0] trunc_ln674_46_fu_6014_p1;
wire   [7:0] tmp_95_fu_6032_p4;
wire   [7:0] xor_ln1545_144_fu_6270_p2;
wire   [7:0] xor_ln1545_142_fu_6266_p2;
wire   [7:0] tmp_92_fu_5990_p4;
wire   [7:0] trunc_ln674_47_fu_6028_p1;
wire   [7:0] xor_ln1545_147_fu_6286_p2;
wire   [7:0] xor_ln1545_145_fu_6282_p2;
wire   [7:0] xor_ln1545_146_fu_6292_p2;
wire   [7:0] xor_ln1545_143_fu_6276_p2;
wire   [7:0] xor_ln1545_140_fu_6260_p2;
wire   [7:0] xor_ln1545_137_fu_6244_p2;
wire   [7:0] xor_ln1545_134_fu_6228_p2;
wire   [7:0] xor_ln1545_131_fu_6212_p2;
wire   [7:0] xor_ln1545_128_fu_6196_p2;
wire   [7:0] xor_ln1545_125_fu_6180_p2;
wire   [7:0] xor_ln1545_122_fu_6164_p2;
wire   [7:0] xor_ln1545_119_fu_6148_p2;
wire   [7:0] xor_ln1545_116_fu_6132_p2;
wire   [7:0] xor_ln1545_113_fu_6116_p2;
wire   [7:0] xor_ln1545_110_fu_6100_p2;
wire   [7:0] xor_ln1545_107_fu_6084_p2;
wire   [7:0] xor_ln1545_104_fu_6068_p2;
wire   [7:0] xor_ln1545_101_fu_6052_p2;
wire   [127:0] p_Result_3_fu_6298_p17;
wire   [127:0] state_V_22_fu_6334_p2;
wire   [7:0] trunc_ln708_3_fu_6339_p1;
wire   [7:0] tmp_96_fu_6348_p4;
wire   [7:0] tmp_97_fu_6363_p4;
wire   [7:0] tmp_98_fu_6378_p4;
wire   [7:0] tmp_99_fu_6393_p4;
wire   [7:0] tmp_100_fu_6408_p4;
wire   [7:0] tmp_101_fu_6423_p4;
wire   [7:0] tmp_102_fu_6438_p4;
wire   [7:0] tmp_103_fu_6453_p4;
wire   [7:0] tmp_104_fu_6468_p4;
wire   [7:0] tmp_105_fu_6483_p4;
wire   [7:0] tmp_106_fu_6498_p4;
wire   [7:0] tmp_107_fu_6513_p4;
wire   [7:0] tmp_108_fu_6528_p4;
wire   [7:0] tmp_109_fu_6543_p4;
wire   [7:0] tmp_110_fu_6558_p4;
wire   [7:0] tmp_112_fu_6671_p4;
wire   [7:0] trunc_ln674_48_fu_6653_p1;
wire   [7:0] xor_ln1545_150_fu_6881_p2;
wire   [7:0] xor_ln1545_148_fu_6877_p2;
wire   [7:0] trunc_ln674_49_fu_6667_p1;
wire   [7:0] tmp_113_fu_6685_p4;
wire   [7:0] xor_ln1545_153_fu_6897_p2;
wire   [7:0] xor_ln1545_151_fu_6893_p2;
wire   [7:0] trunc_ln674_50_fu_6681_p1;
wire   [7:0] tmp_114_fu_6699_p4;
wire   [7:0] xor_ln1545_156_fu_6913_p2;
wire   [7:0] xor_ln1545_154_fu_6909_p2;
wire   [7:0] tmp_111_fu_6657_p4;
wire   [7:0] trunc_ln674_51_fu_6695_p1;
wire   [7:0] xor_ln1545_159_fu_6929_p2;
wire   [7:0] xor_ln1545_157_fu_6925_p2;
wire   [7:0] tmp_116_fu_6727_p4;
wire   [7:0] trunc_ln674_52_fu_6709_p1;
wire   [7:0] xor_ln1545_162_fu_6945_p2;
wire   [7:0] xor_ln1545_160_fu_6941_p2;
wire   [7:0] trunc_ln674_53_fu_6723_p1;
wire   [7:0] tmp_117_fu_6741_p4;
wire   [7:0] xor_ln1545_165_fu_6961_p2;
wire   [7:0] xor_ln1545_163_fu_6957_p2;
wire   [7:0] trunc_ln674_54_fu_6737_p1;
wire   [7:0] tmp_118_fu_6755_p4;
wire   [7:0] xor_ln1545_168_fu_6977_p2;
wire   [7:0] xor_ln1545_166_fu_6973_p2;
wire   [7:0] tmp_115_fu_6713_p4;
wire   [7:0] trunc_ln674_55_fu_6751_p1;
wire   [7:0] xor_ln1545_171_fu_6993_p2;
wire   [7:0] xor_ln1545_169_fu_6989_p2;
wire   [7:0] tmp_120_fu_6783_p4;
wire   [7:0] trunc_ln674_56_fu_6765_p1;
wire   [7:0] xor_ln1545_174_fu_7009_p2;
wire   [7:0] xor_ln1545_172_fu_7005_p2;
wire   [7:0] trunc_ln674_57_fu_6779_p1;
wire   [7:0] tmp_121_fu_6797_p4;
wire   [7:0] xor_ln1545_177_fu_7025_p2;
wire   [7:0] xor_ln1545_175_fu_7021_p2;
wire   [7:0] trunc_ln674_58_fu_6793_p1;
wire   [7:0] tmp_122_fu_6811_p4;
wire   [7:0] xor_ln1545_180_fu_7041_p2;
wire   [7:0] xor_ln1545_178_fu_7037_p2;
wire   [7:0] tmp_119_fu_6769_p4;
wire   [7:0] trunc_ln674_59_fu_6807_p1;
wire   [7:0] xor_ln1545_183_fu_7057_p2;
wire   [7:0] xor_ln1545_181_fu_7053_p2;
wire   [7:0] tmp_124_fu_6839_p4;
wire   [7:0] trunc_ln674_60_fu_6821_p1;
wire   [7:0] xor_ln1545_186_fu_7073_p2;
wire   [7:0] xor_ln1545_184_fu_7069_p2;
wire   [7:0] trunc_ln674_61_fu_6835_p1;
wire   [7:0] tmp_125_fu_6853_p4;
wire   [7:0] xor_ln1545_189_fu_7089_p2;
wire   [7:0] xor_ln1545_187_fu_7085_p2;
wire   [7:0] trunc_ln674_62_fu_6849_p1;
wire   [7:0] tmp_126_fu_6867_p4;
wire   [7:0] xor_ln1545_192_fu_7105_p2;
wire   [7:0] xor_ln1545_190_fu_7101_p2;
wire   [7:0] tmp_123_fu_6825_p4;
wire   [7:0] trunc_ln674_63_fu_6863_p1;
wire   [7:0] xor_ln1545_195_fu_7121_p2;
wire   [7:0] xor_ln1545_193_fu_7117_p2;
wire   [7:0] xor_ln1545_194_fu_7127_p2;
wire   [7:0] xor_ln1545_191_fu_7111_p2;
wire   [7:0] xor_ln1545_188_fu_7095_p2;
wire   [7:0] xor_ln1545_185_fu_7079_p2;
wire   [7:0] xor_ln1545_182_fu_7063_p2;
wire   [7:0] xor_ln1545_179_fu_7047_p2;
wire   [7:0] xor_ln1545_176_fu_7031_p2;
wire   [7:0] xor_ln1545_173_fu_7015_p2;
wire   [7:0] xor_ln1545_170_fu_6999_p2;
wire   [7:0] xor_ln1545_167_fu_6983_p2;
wire   [7:0] xor_ln1545_164_fu_6967_p2;
wire   [7:0] xor_ln1545_161_fu_6951_p2;
wire   [7:0] xor_ln1545_158_fu_6935_p2;
wire   [7:0] xor_ln1545_155_fu_6919_p2;
wire   [7:0] xor_ln1545_152_fu_6903_p2;
wire   [7:0] xor_ln1545_149_fu_6887_p2;
wire   [127:0] p_Result_4_fu_7133_p17;
wire   [127:0] state_V_23_fu_7169_p2;
wire   [7:0] trunc_ln708_4_fu_7174_p1;
wire   [7:0] tmp_127_fu_7183_p4;
wire   [7:0] tmp_128_fu_7198_p4;
wire   [7:0] tmp_129_fu_7213_p4;
wire   [7:0] tmp_130_fu_7228_p4;
wire   [7:0] tmp_131_fu_7243_p4;
wire   [7:0] tmp_132_fu_7258_p4;
wire   [7:0] tmp_133_fu_7273_p4;
wire   [7:0] tmp_134_fu_7288_p4;
wire   [7:0] tmp_135_fu_7303_p4;
wire   [7:0] tmp_136_fu_7318_p4;
wire   [7:0] tmp_137_fu_7333_p4;
wire   [7:0] tmp_138_fu_7348_p4;
wire   [7:0] tmp_139_fu_7363_p4;
wire   [7:0] tmp_140_fu_7378_p4;
wire   [7:0] tmp_141_fu_7393_p4;
wire   [7:0] tmp_143_fu_7506_p4;
wire   [7:0] trunc_ln674_64_fu_7488_p1;
wire   [7:0] xor_ln1545_198_fu_7716_p2;
wire   [7:0] xor_ln1545_196_fu_7712_p2;
wire   [7:0] trunc_ln674_65_fu_7502_p1;
wire   [7:0] tmp_144_fu_7520_p4;
wire   [7:0] xor_ln1545_201_fu_7732_p2;
wire   [7:0] xor_ln1545_199_fu_7728_p2;
wire   [7:0] trunc_ln674_66_fu_7516_p1;
wire   [7:0] tmp_145_fu_7534_p4;
wire   [7:0] xor_ln1545_204_fu_7748_p2;
wire   [7:0] xor_ln1545_202_fu_7744_p2;
wire   [7:0] tmp_142_fu_7492_p4;
wire   [7:0] trunc_ln674_67_fu_7530_p1;
wire   [7:0] xor_ln1545_207_fu_7764_p2;
wire   [7:0] xor_ln1545_205_fu_7760_p2;
wire   [7:0] tmp_147_fu_7562_p4;
wire   [7:0] trunc_ln674_68_fu_7544_p1;
wire   [7:0] xor_ln1545_210_fu_7780_p2;
wire   [7:0] xor_ln1545_208_fu_7776_p2;
wire   [7:0] trunc_ln674_69_fu_7558_p1;
wire   [7:0] tmp_148_fu_7576_p4;
wire   [7:0] xor_ln1545_213_fu_7796_p2;
wire   [7:0] xor_ln1545_211_fu_7792_p2;
wire   [7:0] trunc_ln674_70_fu_7572_p1;
wire   [7:0] tmp_149_fu_7590_p4;
wire   [7:0] xor_ln1545_216_fu_7812_p2;
wire   [7:0] xor_ln1545_214_fu_7808_p2;
wire   [7:0] tmp_146_fu_7548_p4;
wire   [7:0] trunc_ln674_71_fu_7586_p1;
wire   [7:0] xor_ln1545_219_fu_7828_p2;
wire   [7:0] xor_ln1545_217_fu_7824_p2;
wire   [7:0] tmp_151_fu_7618_p4;
wire   [7:0] trunc_ln674_72_fu_7600_p1;
wire   [7:0] xor_ln1545_222_fu_7844_p2;
wire   [7:0] xor_ln1545_220_fu_7840_p2;
wire   [7:0] trunc_ln674_73_fu_7614_p1;
wire   [7:0] tmp_152_fu_7632_p4;
wire   [7:0] xor_ln1545_225_fu_7860_p2;
wire   [7:0] xor_ln1545_223_fu_7856_p2;
wire   [7:0] trunc_ln674_74_fu_7628_p1;
wire   [7:0] tmp_153_fu_7646_p4;
wire   [7:0] xor_ln1545_228_fu_7876_p2;
wire   [7:0] xor_ln1545_226_fu_7872_p2;
wire   [7:0] tmp_150_fu_7604_p4;
wire   [7:0] trunc_ln674_75_fu_7642_p1;
wire   [7:0] xor_ln1545_231_fu_7892_p2;
wire   [7:0] xor_ln1545_229_fu_7888_p2;
wire   [7:0] tmp_155_fu_7674_p4;
wire   [7:0] trunc_ln674_76_fu_7656_p1;
wire   [7:0] xor_ln1545_234_fu_7908_p2;
wire   [7:0] xor_ln1545_232_fu_7904_p2;
wire   [7:0] trunc_ln674_77_fu_7670_p1;
wire   [7:0] tmp_156_fu_7688_p4;
wire   [7:0] xor_ln1545_237_fu_7924_p2;
wire   [7:0] xor_ln1545_235_fu_7920_p2;
wire   [7:0] trunc_ln674_78_fu_7684_p1;
wire   [7:0] tmp_157_fu_7702_p4;
wire   [7:0] xor_ln1545_240_fu_7940_p2;
wire   [7:0] xor_ln1545_238_fu_7936_p2;
wire   [7:0] tmp_154_fu_7660_p4;
wire   [7:0] trunc_ln674_79_fu_7698_p1;
wire   [7:0] xor_ln1545_243_fu_7956_p2;
wire   [7:0] xor_ln1545_241_fu_7952_p2;
wire   [7:0] xor_ln1545_242_fu_7962_p2;
wire   [7:0] xor_ln1545_239_fu_7946_p2;
wire   [7:0] xor_ln1545_236_fu_7930_p2;
wire   [7:0] xor_ln1545_233_fu_7914_p2;
wire   [7:0] xor_ln1545_230_fu_7898_p2;
wire   [7:0] xor_ln1545_227_fu_7882_p2;
wire   [7:0] xor_ln1545_224_fu_7866_p2;
wire   [7:0] xor_ln1545_221_fu_7850_p2;
wire   [7:0] xor_ln1545_218_fu_7834_p2;
wire   [7:0] xor_ln1545_215_fu_7818_p2;
wire   [7:0] xor_ln1545_212_fu_7802_p2;
wire   [7:0] xor_ln1545_209_fu_7786_p2;
wire   [7:0] xor_ln1545_206_fu_7770_p2;
wire   [7:0] xor_ln1545_203_fu_7754_p2;
wire   [7:0] xor_ln1545_200_fu_7738_p2;
wire   [7:0] xor_ln1545_197_fu_7722_p2;
wire   [127:0] p_Result_5_fu_7968_p17;
wire   [127:0] state_V_24_fu_8004_p2;
wire   [7:0] trunc_ln708_5_fu_8009_p1;
wire   [7:0] tmp_158_fu_8018_p4;
wire   [7:0] tmp_159_fu_8033_p4;
wire   [7:0] tmp_160_fu_8048_p4;
wire   [7:0] tmp_161_fu_8063_p4;
wire   [7:0] tmp_162_fu_8078_p4;
wire   [7:0] tmp_163_fu_8093_p4;
wire   [7:0] tmp_164_fu_8108_p4;
wire   [7:0] tmp_165_fu_8123_p4;
wire   [7:0] tmp_166_fu_8138_p4;
wire   [7:0] tmp_167_fu_8153_p4;
wire   [7:0] tmp_168_fu_8168_p4;
wire   [7:0] tmp_169_fu_8183_p4;
wire   [7:0] tmp_170_fu_8198_p4;
wire   [7:0] tmp_171_fu_8213_p4;
wire   [7:0] tmp_172_fu_8228_p4;
wire   [7:0] tmp_174_fu_8341_p4;
wire   [7:0] trunc_ln674_80_fu_8323_p1;
wire   [7:0] xor_ln1545_246_fu_8551_p2;
wire   [7:0] xor_ln1545_244_fu_8547_p2;
wire   [7:0] trunc_ln674_81_fu_8337_p1;
wire   [7:0] tmp_175_fu_8355_p4;
wire   [7:0] xor_ln1545_249_fu_8567_p2;
wire   [7:0] xor_ln1545_247_fu_8563_p2;
wire   [7:0] trunc_ln674_82_fu_8351_p1;
wire   [7:0] tmp_176_fu_8369_p4;
wire   [7:0] xor_ln1545_252_fu_8583_p2;
wire   [7:0] xor_ln1545_250_fu_8579_p2;
wire   [7:0] tmp_173_fu_8327_p4;
wire   [7:0] trunc_ln674_83_fu_8365_p1;
wire   [7:0] xor_ln1545_255_fu_8599_p2;
wire   [7:0] xor_ln1545_253_fu_8595_p2;
wire   [7:0] tmp_178_fu_8397_p4;
wire   [7:0] trunc_ln674_84_fu_8379_p1;
wire   [7:0] xor_ln1545_258_fu_8615_p2;
wire   [7:0] xor_ln1545_256_fu_8611_p2;
wire   [7:0] trunc_ln674_85_fu_8393_p1;
wire   [7:0] tmp_179_fu_8411_p4;
wire   [7:0] xor_ln1545_261_fu_8631_p2;
wire   [7:0] xor_ln1545_259_fu_8627_p2;
wire   [7:0] trunc_ln674_86_fu_8407_p1;
wire   [7:0] tmp_180_fu_8425_p4;
wire   [7:0] xor_ln1545_264_fu_8647_p2;
wire   [7:0] xor_ln1545_262_fu_8643_p2;
wire   [7:0] tmp_177_fu_8383_p4;
wire   [7:0] trunc_ln674_87_fu_8421_p1;
wire   [7:0] xor_ln1545_267_fu_8663_p2;
wire   [7:0] xor_ln1545_265_fu_8659_p2;
wire   [7:0] tmp_182_fu_8453_p4;
wire   [7:0] trunc_ln674_88_fu_8435_p1;
wire   [7:0] xor_ln1545_270_fu_8679_p2;
wire   [7:0] xor_ln1545_268_fu_8675_p2;
wire   [7:0] trunc_ln674_89_fu_8449_p1;
wire   [7:0] tmp_183_fu_8467_p4;
wire   [7:0] xor_ln1545_273_fu_8695_p2;
wire   [7:0] xor_ln1545_271_fu_8691_p2;
wire   [7:0] trunc_ln674_90_fu_8463_p1;
wire   [7:0] tmp_184_fu_8481_p4;
wire   [7:0] xor_ln1545_276_fu_8711_p2;
wire   [7:0] xor_ln1545_274_fu_8707_p2;
wire   [7:0] tmp_181_fu_8439_p4;
wire   [7:0] trunc_ln674_91_fu_8477_p1;
wire   [7:0] xor_ln1545_279_fu_8727_p2;
wire   [7:0] xor_ln1545_277_fu_8723_p2;
wire   [7:0] tmp_186_fu_8509_p4;
wire   [7:0] trunc_ln674_92_fu_8491_p1;
wire   [7:0] xor_ln1545_282_fu_8743_p2;
wire   [7:0] xor_ln1545_280_fu_8739_p2;
wire   [7:0] trunc_ln674_93_fu_8505_p1;
wire   [7:0] tmp_187_fu_8523_p4;
wire   [7:0] xor_ln1545_285_fu_8759_p2;
wire   [7:0] xor_ln1545_283_fu_8755_p2;
wire   [7:0] trunc_ln674_94_fu_8519_p1;
wire   [7:0] tmp_188_fu_8537_p4;
wire   [7:0] xor_ln1545_288_fu_8775_p2;
wire   [7:0] xor_ln1545_286_fu_8771_p2;
wire   [7:0] tmp_185_fu_8495_p4;
wire   [7:0] trunc_ln674_95_fu_8533_p1;
wire   [7:0] xor_ln1545_291_fu_8791_p2;
wire   [7:0] xor_ln1545_289_fu_8787_p2;
wire   [7:0] xor_ln1545_290_fu_8797_p2;
wire   [7:0] xor_ln1545_287_fu_8781_p2;
wire   [7:0] xor_ln1545_284_fu_8765_p2;
wire   [7:0] xor_ln1545_281_fu_8749_p2;
wire   [7:0] xor_ln1545_278_fu_8733_p2;
wire   [7:0] xor_ln1545_275_fu_8717_p2;
wire   [7:0] xor_ln1545_272_fu_8701_p2;
wire   [7:0] xor_ln1545_269_fu_8685_p2;
wire   [7:0] xor_ln1545_266_fu_8669_p2;
wire   [7:0] xor_ln1545_263_fu_8653_p2;
wire   [7:0] xor_ln1545_260_fu_8637_p2;
wire   [7:0] xor_ln1545_257_fu_8621_p2;
wire   [7:0] xor_ln1545_254_fu_8605_p2;
wire   [7:0] xor_ln1545_251_fu_8589_p2;
wire   [7:0] xor_ln1545_248_fu_8573_p2;
wire   [7:0] xor_ln1545_245_fu_8557_p2;
wire   [127:0] p_Result_6_fu_8803_p17;
wire   [127:0] state_V_25_fu_8839_p2;
wire   [7:0] trunc_ln708_6_fu_8844_p1;
wire   [7:0] tmp_189_fu_8853_p4;
wire   [7:0] tmp_190_fu_8868_p4;
wire   [7:0] tmp_191_fu_8883_p4;
wire   [7:0] tmp_192_fu_8898_p4;
wire   [7:0] tmp_193_fu_8913_p4;
wire   [7:0] tmp_194_fu_8928_p4;
wire   [7:0] tmp_195_fu_8943_p4;
wire   [7:0] tmp_196_fu_8958_p4;
wire   [7:0] tmp_197_fu_8973_p4;
wire   [7:0] tmp_198_fu_8988_p4;
wire   [7:0] tmp_199_fu_9003_p4;
wire   [7:0] tmp_200_fu_9018_p4;
wire   [7:0] tmp_201_fu_9033_p4;
wire   [7:0] tmp_202_fu_9048_p4;
wire   [7:0] tmp_203_fu_9063_p4;
wire   [7:0] tmp_205_fu_9176_p4;
wire   [7:0] trunc_ln674_96_fu_9158_p1;
wire   [7:0] xor_ln1545_294_fu_9386_p2;
wire   [7:0] xor_ln1545_292_fu_9382_p2;
wire   [7:0] trunc_ln674_97_fu_9172_p1;
wire   [7:0] tmp_206_fu_9190_p4;
wire   [7:0] xor_ln1545_297_fu_9402_p2;
wire   [7:0] xor_ln1545_295_fu_9398_p2;
wire   [7:0] trunc_ln674_98_fu_9186_p1;
wire   [7:0] tmp_207_fu_9204_p4;
wire   [7:0] xor_ln1545_300_fu_9418_p2;
wire   [7:0] xor_ln1545_298_fu_9414_p2;
wire   [7:0] tmp_204_fu_9162_p4;
wire   [7:0] trunc_ln674_99_fu_9200_p1;
wire   [7:0] xor_ln1545_303_fu_9434_p2;
wire   [7:0] xor_ln1545_301_fu_9430_p2;
wire   [7:0] tmp_209_fu_9232_p4;
wire   [7:0] trunc_ln674_100_fu_9214_p1;
wire   [7:0] xor_ln1545_306_fu_9450_p2;
wire   [7:0] xor_ln1545_304_fu_9446_p2;
wire   [7:0] trunc_ln674_101_fu_9228_p1;
wire   [7:0] tmp_210_fu_9246_p4;
wire   [7:0] xor_ln1545_309_fu_9466_p2;
wire   [7:0] xor_ln1545_307_fu_9462_p2;
wire   [7:0] trunc_ln674_102_fu_9242_p1;
wire   [7:0] tmp_211_fu_9260_p4;
wire   [7:0] xor_ln1545_312_fu_9482_p2;
wire   [7:0] xor_ln1545_310_fu_9478_p2;
wire   [7:0] tmp_208_fu_9218_p4;
wire   [7:0] trunc_ln674_103_fu_9256_p1;
wire   [7:0] xor_ln1545_315_fu_9498_p2;
wire   [7:0] xor_ln1545_313_fu_9494_p2;
wire   [7:0] tmp_213_fu_9288_p4;
wire   [7:0] trunc_ln674_104_fu_9270_p1;
wire   [7:0] xor_ln1545_318_fu_9514_p2;
wire   [7:0] xor_ln1545_316_fu_9510_p2;
wire   [7:0] trunc_ln674_105_fu_9284_p1;
wire   [7:0] tmp_214_fu_9302_p4;
wire   [7:0] xor_ln1545_321_fu_9530_p2;
wire   [7:0] xor_ln1545_319_fu_9526_p2;
wire   [7:0] trunc_ln674_106_fu_9298_p1;
wire   [7:0] tmp_215_fu_9316_p4;
wire   [7:0] xor_ln1545_324_fu_9546_p2;
wire   [7:0] xor_ln1545_322_fu_9542_p2;
wire   [7:0] tmp_212_fu_9274_p4;
wire   [7:0] trunc_ln674_107_fu_9312_p1;
wire   [7:0] xor_ln1545_327_fu_9562_p2;
wire   [7:0] xor_ln1545_325_fu_9558_p2;
wire   [7:0] tmp_217_fu_9344_p4;
wire   [7:0] trunc_ln674_108_fu_9326_p1;
wire   [7:0] xor_ln1545_330_fu_9578_p2;
wire   [7:0] xor_ln1545_328_fu_9574_p2;
wire   [7:0] trunc_ln674_109_fu_9340_p1;
wire   [7:0] tmp_218_fu_9358_p4;
wire   [7:0] xor_ln1545_333_fu_9594_p2;
wire   [7:0] xor_ln1545_331_fu_9590_p2;
wire   [7:0] trunc_ln674_110_fu_9354_p1;
wire   [7:0] tmp_219_fu_9372_p4;
wire   [7:0] xor_ln1545_336_fu_9610_p2;
wire   [7:0] xor_ln1545_334_fu_9606_p2;
wire   [7:0] tmp_216_fu_9330_p4;
wire   [7:0] trunc_ln674_111_fu_9368_p1;
wire   [7:0] xor_ln1545_339_fu_9626_p2;
wire   [7:0] xor_ln1545_337_fu_9622_p2;
wire   [7:0] xor_ln1545_338_fu_9632_p2;
wire   [7:0] xor_ln1545_335_fu_9616_p2;
wire   [7:0] xor_ln1545_332_fu_9600_p2;
wire   [7:0] xor_ln1545_329_fu_9584_p2;
wire   [7:0] xor_ln1545_326_fu_9568_p2;
wire   [7:0] xor_ln1545_323_fu_9552_p2;
wire   [7:0] xor_ln1545_320_fu_9536_p2;
wire   [7:0] xor_ln1545_317_fu_9520_p2;
wire   [7:0] xor_ln1545_314_fu_9504_p2;
wire   [7:0] xor_ln1545_311_fu_9488_p2;
wire   [7:0] xor_ln1545_308_fu_9472_p2;
wire   [7:0] xor_ln1545_305_fu_9456_p2;
wire   [7:0] xor_ln1545_302_fu_9440_p2;
wire   [7:0] xor_ln1545_299_fu_9424_p2;
wire   [7:0] xor_ln1545_296_fu_9408_p2;
wire   [7:0] xor_ln1545_293_fu_9392_p2;
wire   [127:0] p_Result_7_fu_9638_p17;
wire   [127:0] state_V_fu_9674_p2;
wire   [7:0] trunc_ln708_7_fu_9679_p1;
wire   [7:0] tmp_220_fu_9688_p4;
wire   [7:0] tmp_221_fu_9703_p4;
wire   [7:0] tmp_222_fu_9718_p4;
wire   [7:0] tmp_223_fu_9733_p4;
wire   [7:0] tmp_224_fu_9748_p4;
wire   [7:0] tmp_225_fu_9763_p4;
wire   [7:0] tmp_226_fu_9778_p4;
wire   [7:0] tmp_227_fu_9793_p4;
wire   [7:0] tmp_228_fu_9808_p4;
wire   [7:0] tmp_229_fu_9823_p4;
wire   [7:0] tmp_230_fu_9838_p4;
wire   [7:0] tmp_231_fu_9853_p4;
wire   [7:0] tmp_232_fu_9868_p4;
wire   [7:0] tmp_233_fu_9883_p4;
wire   [7:0] tmp_234_fu_9898_p4;
wire   [7:0] tmp_236_fu_10011_p4;
wire   [7:0] trunc_ln674_112_fu_9993_p1;
wire   [7:0] xor_ln1545_342_fu_10221_p2;
wire   [7:0] xor_ln1545_340_fu_10217_p2;
wire   [7:0] trunc_ln674_113_fu_10007_p1;
wire   [7:0] tmp_237_fu_10025_p4;
wire   [7:0] xor_ln1545_345_fu_10237_p2;
wire   [7:0] xor_ln1545_343_fu_10233_p2;
wire   [7:0] trunc_ln674_114_fu_10021_p1;
wire   [7:0] tmp_238_fu_10039_p4;
wire   [7:0] xor_ln1545_348_fu_10253_p2;
wire   [7:0] xor_ln1545_346_fu_10249_p2;
wire   [7:0] tmp_235_fu_9997_p4;
wire   [7:0] trunc_ln674_115_fu_10035_p1;
wire   [7:0] xor_ln1545_351_fu_10269_p2;
wire   [7:0] xor_ln1545_349_fu_10265_p2;
wire   [7:0] tmp_240_fu_10067_p4;
wire   [7:0] trunc_ln674_116_fu_10049_p1;
wire   [7:0] xor_ln1545_354_fu_10285_p2;
wire   [7:0] xor_ln1545_352_fu_10281_p2;
wire   [7:0] trunc_ln674_117_fu_10063_p1;
wire   [7:0] tmp_241_fu_10081_p4;
wire   [7:0] xor_ln1545_357_fu_10301_p2;
wire   [7:0] xor_ln1545_355_fu_10297_p2;
wire   [7:0] trunc_ln674_118_fu_10077_p1;
wire   [7:0] tmp_242_fu_10095_p4;
wire   [7:0] xor_ln1545_360_fu_10317_p2;
wire   [7:0] xor_ln1545_358_fu_10313_p2;
wire   [7:0] tmp_239_fu_10053_p4;
wire   [7:0] trunc_ln674_119_fu_10091_p1;
wire   [7:0] xor_ln1545_363_fu_10333_p2;
wire   [7:0] xor_ln1545_361_fu_10329_p2;
wire   [7:0] tmp_244_fu_10123_p4;
wire   [7:0] trunc_ln674_120_fu_10105_p1;
wire   [7:0] xor_ln1545_366_fu_10349_p2;
wire   [7:0] xor_ln1545_364_fu_10345_p2;
wire   [7:0] trunc_ln674_121_fu_10119_p1;
wire   [7:0] tmp_245_fu_10137_p4;
wire   [7:0] xor_ln1545_369_fu_10365_p2;
wire   [7:0] xor_ln1545_367_fu_10361_p2;
wire   [7:0] trunc_ln674_122_fu_10133_p1;
wire   [7:0] tmp_246_fu_10151_p4;
wire   [7:0] xor_ln1545_372_fu_10381_p2;
wire   [7:0] xor_ln1545_370_fu_10377_p2;
wire   [7:0] tmp_243_fu_10109_p4;
wire   [7:0] trunc_ln674_123_fu_10147_p1;
wire   [7:0] xor_ln1545_375_fu_10397_p2;
wire   [7:0] xor_ln1545_373_fu_10393_p2;
wire   [7:0] tmp_248_fu_10179_p4;
wire   [7:0] trunc_ln674_124_fu_10161_p1;
wire   [7:0] xor_ln1545_378_fu_10413_p2;
wire   [7:0] xor_ln1545_376_fu_10409_p2;
wire   [7:0] trunc_ln674_125_fu_10175_p1;
wire   [7:0] tmp_249_fu_10193_p4;
wire   [7:0] xor_ln1545_381_fu_10429_p2;
wire   [7:0] xor_ln1545_379_fu_10425_p2;
wire   [7:0] trunc_ln674_126_fu_10189_p1;
wire   [7:0] tmp_250_fu_10207_p4;
wire   [7:0] xor_ln1545_384_fu_10445_p2;
wire   [7:0] xor_ln1545_382_fu_10441_p2;
wire   [7:0] tmp_247_fu_10165_p4;
wire   [7:0] trunc_ln674_127_fu_10203_p1;
wire   [7:0] xor_ln1545_387_fu_10461_p2;
wire   [7:0] xor_ln1545_385_fu_10457_p2;
wire   [7:0] xor_ln1545_386_fu_10467_p2;
wire   [7:0] xor_ln1545_383_fu_10451_p2;
wire   [7:0] xor_ln1545_380_fu_10435_p2;
wire   [7:0] xor_ln1545_377_fu_10419_p2;
wire   [7:0] xor_ln1545_374_fu_10403_p2;
wire   [7:0] xor_ln1545_371_fu_10387_p2;
wire   [7:0] xor_ln1545_368_fu_10371_p2;
wire   [7:0] xor_ln1545_365_fu_10355_p2;
wire   [7:0] xor_ln1545_362_fu_10339_p2;
wire   [7:0] xor_ln1545_359_fu_10323_p2;
wire   [7:0] xor_ln1545_356_fu_10307_p2;
wire   [7:0] xor_ln1545_353_fu_10291_p2;
wire   [7:0] xor_ln1545_350_fu_10275_p2;
wire   [7:0] xor_ln1545_347_fu_10259_p2;
wire   [7:0] xor_ln1545_344_fu_10243_p2;
wire   [7:0] xor_ln1545_341_fu_10227_p2;
wire   [127:0] p_Result_8_fu_10473_p17;
wire   [127:0] state_V_26_fu_10509_p2;
wire   [7:0] trunc_ln708_8_fu_10514_p1;
wire   [7:0] tmp_251_fu_10523_p4;
wire   [7:0] tmp_252_fu_10538_p4;
wire   [7:0] tmp_253_fu_10553_p4;
wire   [7:0] tmp_254_fu_10568_p4;
wire   [7:0] tmp_255_fu_10583_p4;
wire   [7:0] tmp_256_fu_10598_p4;
wire   [7:0] tmp_257_fu_10613_p4;
wire   [7:0] tmp_258_fu_10628_p4;
wire   [7:0] tmp_259_fu_10643_p4;
wire   [7:0] tmp_260_fu_10658_p4;
wire   [7:0] tmp_261_fu_10673_p4;
wire   [7:0] tmp_262_fu_10688_p4;
wire   [7:0] tmp_263_fu_10703_p4;
wire   [7:0] tmp_264_fu_10718_p4;
wire   [7:0] tmp_265_fu_10733_p4;
wire   [7:0] tmp_267_fu_10846_p4;
wire   [7:0] trunc_ln674_128_fu_10828_p1;
wire   [7:0] xor_ln1545_390_fu_11056_p2;
wire   [7:0] xor_ln1545_388_fu_11052_p2;
wire   [7:0] trunc_ln674_129_fu_10842_p1;
wire   [7:0] tmp_268_fu_10860_p4;
wire   [7:0] xor_ln1545_393_fu_11072_p2;
wire   [7:0] xor_ln1545_391_fu_11068_p2;
wire   [7:0] trunc_ln674_130_fu_10856_p1;
wire   [7:0] tmp_269_fu_10874_p4;
wire   [7:0] xor_ln1545_396_fu_11088_p2;
wire   [7:0] xor_ln1545_394_fu_11084_p2;
wire   [7:0] tmp_266_fu_10832_p4;
wire   [7:0] trunc_ln674_131_fu_10870_p1;
wire   [7:0] xor_ln1545_399_fu_11104_p2;
wire   [7:0] xor_ln1545_397_fu_11100_p2;
wire   [7:0] tmp_271_fu_10902_p4;
wire   [7:0] trunc_ln674_132_fu_10884_p1;
wire   [7:0] xor_ln1545_402_fu_11120_p2;
wire   [7:0] xor_ln1545_400_fu_11116_p2;
wire   [7:0] trunc_ln674_133_fu_10898_p1;
wire   [7:0] tmp_272_fu_10916_p4;
wire   [7:0] xor_ln1545_405_fu_11136_p2;
wire   [7:0] xor_ln1545_403_fu_11132_p2;
wire   [7:0] trunc_ln674_134_fu_10912_p1;
wire   [7:0] tmp_273_fu_10930_p4;
wire   [7:0] xor_ln1545_408_fu_11152_p2;
wire   [7:0] xor_ln1545_406_fu_11148_p2;
wire   [7:0] tmp_270_fu_10888_p4;
wire   [7:0] trunc_ln674_135_fu_10926_p1;
wire   [7:0] xor_ln1545_411_fu_11168_p2;
wire   [7:0] xor_ln1545_409_fu_11164_p2;
wire   [7:0] tmp_275_fu_10958_p4;
wire   [7:0] trunc_ln674_136_fu_10940_p1;
wire   [7:0] xor_ln1545_414_fu_11184_p2;
wire   [7:0] xor_ln1545_412_fu_11180_p2;
wire   [7:0] trunc_ln674_137_fu_10954_p1;
wire   [7:0] tmp_276_fu_10972_p4;
wire   [7:0] xor_ln1545_417_fu_11200_p2;
wire   [7:0] xor_ln1545_415_fu_11196_p2;
wire   [7:0] trunc_ln674_138_fu_10968_p1;
wire   [7:0] tmp_277_fu_10986_p4;
wire   [7:0] xor_ln1545_420_fu_11216_p2;
wire   [7:0] xor_ln1545_418_fu_11212_p2;
wire   [7:0] tmp_274_fu_10944_p4;
wire   [7:0] trunc_ln674_139_fu_10982_p1;
wire   [7:0] xor_ln1545_423_fu_11232_p2;
wire   [7:0] xor_ln1545_421_fu_11228_p2;
wire   [7:0] tmp_279_fu_11014_p4;
wire   [7:0] trunc_ln674_140_fu_10996_p1;
wire   [7:0] xor_ln1545_426_fu_11248_p2;
wire   [7:0] xor_ln1545_424_fu_11244_p2;
wire   [7:0] trunc_ln674_141_fu_11010_p1;
wire   [7:0] tmp_280_fu_11028_p4;
wire   [7:0] xor_ln1545_429_fu_11264_p2;
wire   [7:0] xor_ln1545_427_fu_11260_p2;
wire   [7:0] trunc_ln674_142_fu_11024_p1;
wire   [7:0] tmp_281_fu_11042_p4;
wire   [7:0] xor_ln1545_432_fu_11280_p2;
wire   [7:0] xor_ln1545_430_fu_11276_p2;
wire   [7:0] tmp_278_fu_11000_p4;
wire   [7:0] trunc_ln674_143_fu_11038_p1;
wire   [7:0] xor_ln1545_435_fu_11296_p2;
wire   [7:0] xor_ln1545_433_fu_11292_p2;
wire   [7:0] xor_ln1545_434_fu_11302_p2;
wire   [7:0] xor_ln1545_431_fu_11286_p2;
wire   [7:0] xor_ln1545_428_fu_11270_p2;
wire   [7:0] xor_ln1545_425_fu_11254_p2;
wire   [7:0] xor_ln1545_422_fu_11238_p2;
wire   [7:0] xor_ln1545_419_fu_11222_p2;
wire   [7:0] xor_ln1545_416_fu_11206_p2;
wire   [7:0] xor_ln1545_413_fu_11190_p2;
wire   [7:0] xor_ln1545_410_fu_11174_p2;
wire   [7:0] xor_ln1545_407_fu_11158_p2;
wire   [7:0] xor_ln1545_404_fu_11142_p2;
wire   [7:0] xor_ln1545_401_fu_11126_p2;
wire   [7:0] xor_ln1545_398_fu_11110_p2;
wire   [7:0] xor_ln1545_395_fu_11094_p2;
wire   [7:0] xor_ln1545_392_fu_11078_p2;
wire   [7:0] xor_ln1545_389_fu_11062_p2;
wire   [127:0] p_Result_9_fu_11308_p17;
wire   [127:0] state_V_27_fu_11344_p2;
wire   [7:0] trunc_ln708_9_fu_11349_p1;
wire   [7:0] tmp_282_fu_11358_p4;
wire   [7:0] tmp_283_fu_11373_p4;
wire   [7:0] tmp_284_fu_11388_p4;
wire   [7:0] tmp_285_fu_11403_p4;
wire   [7:0] tmp_286_fu_11418_p4;
wire   [7:0] tmp_287_fu_11433_p4;
wire   [7:0] tmp_288_fu_11448_p4;
wire   [7:0] tmp_289_fu_11463_p4;
wire   [7:0] tmp_290_fu_11478_p4;
wire   [7:0] tmp_291_fu_11493_p4;
wire   [7:0] tmp_292_fu_11508_p4;
wire   [7:0] tmp_293_fu_11523_p4;
wire   [7:0] tmp_294_fu_11538_p4;
wire   [7:0] tmp_295_fu_11553_p4;
wire   [7:0] tmp_296_fu_11568_p4;
wire   [127:0] p_Result_10_fu_11583_p17;
reg   [0:0] ap_NS_fsm;
reg    ap_idle_pp0_0to18;
reg    ap_reset_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 1'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter5 = 1'b0;
#0 ap_enable_reg_pp0_iter6 = 1'b0;
#0 ap_enable_reg_pp0_iter7 = 1'b0;
#0 ap_enable_reg_pp0_iter8 = 1'b0;
#0 ap_enable_reg_pp0_iter9 = 1'b0;
#0 ap_enable_reg_pp0_iter10 = 1'b0;
#0 ap_enable_reg_pp0_iter11 = 1'b0;
#0 ap_enable_reg_pp0_iter12 = 1'b0;
#0 ap_enable_reg_pp0_iter13 = 1'b0;
#0 ap_enable_reg_pp0_iter14 = 1'b0;
#0 ap_enable_reg_pp0_iter15 = 1'b0;
#0 ap_enable_reg_pp0_iter16 = 1'b0;
#0 ap_enable_reg_pp0_iter17 = 1'b0;
#0 ap_enable_reg_pp0_iter18 = 1'b0;
#0 ap_enable_reg_pp0_iter19 = 1'b0;
end

testEnc_process_r_cipher_0_ssbox_ROM_NP_LUTRAM_1R #(
    .DataWidth( 8 ),
    .AddressRange( 256 ),
    .AddressWidth( 8 ))
cipher_0_ssbox_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(cipher_0_ssbox_address0),
    .ce0(cipher_0_ssbox_ce0),
    .q0(cipher_0_ssbox_q0),
    .address1(cipher_0_ssbox_address1),
    .ce1(cipher_0_ssbox_ce1),
    .q1(cipher_0_ssbox_q1),
    .address2(cipher_0_ssbox_address2),
    .ce2(cipher_0_ssbox_ce2),
    .q2(cipher_0_ssbox_q2),
    .address3(cipher_0_ssbox_address3),
    .ce3(cipher_0_ssbox_ce3),
    .q3(cipher_0_ssbox_q3),
    .address4(cipher_0_ssbox_address4),
    .ce4(cipher_0_ssbox_ce4),
    .q4(cipher_0_ssbox_q4),
    .address5(cipher_0_ssbox_address5),
    .ce5(cipher_0_ssbox_ce5),
    .q5(cipher_0_ssbox_q5),
    .address6(cipher_0_ssbox_address6),
    .ce6(cipher_0_ssbox_ce6),
    .q6(cipher_0_ssbox_q6),
    .address7(cipher_0_ssbox_address7),
    .ce7(cipher_0_ssbox_ce7),
    .q7(cipher_0_ssbox_q7),
    .address8(cipher_0_ssbox_address8),
    .ce8(cipher_0_ssbox_ce8),
    .q8(cipher_0_ssbox_q8),
    .address9(cipher_0_ssbox_address9),
    .ce9(cipher_0_ssbox_ce9),
    .q9(cipher_0_ssbox_q9),
    .address10(cipher_0_ssbox_address10),
    .ce10(cipher_0_ssbox_ce10),
    .q10(cipher_0_ssbox_q10),
    .address11(cipher_0_ssbox_address11),
    .ce11(cipher_0_ssbox_ce11),
    .q11(cipher_0_ssbox_q11),
    .address12(cipher_0_ssbox_address12),
    .ce12(cipher_0_ssbox_ce12),
    .q12(cipher_0_ssbox_q12),
    .address13(cipher_0_ssbox_address13),
    .ce13(cipher_0_ssbox_ce13),
    .q13(cipher_0_ssbox_q13),
    .address14(cipher_0_ssbox_address14),
    .ce14(cipher_0_ssbox_ce14),
    .q14(cipher_0_ssbox_q14),
    .address15(cipher_0_ssbox_address15),
    .ce15(cipher_0_ssbox_ce15),
    .q15(cipher_0_ssbox_q15),
    .address16(cipher_0_ssbox_address16),
    .ce16(cipher_0_ssbox_ce16),
    .q16(cipher_0_ssbox_q16),
    .address17(cipher_0_ssbox_address17),
    .ce17(cipher_0_ssbox_ce17),
    .q17(cipher_0_ssbox_q17),
    .address18(cipher_0_ssbox_address18),
    .ce18(cipher_0_ssbox_ce18),
    .q18(cipher_0_ssbox_q18),
    .address19(cipher_0_ssbox_address19),
    .ce19(cipher_0_ssbox_ce19),
    .q19(cipher_0_ssbox_q19),
    .address20(cipher_0_ssbox_address20),
    .ce20(cipher_0_ssbox_ce20),
    .q20(cipher_0_ssbox_q20),
    .address21(cipher_0_ssbox_address21),
    .ce21(cipher_0_ssbox_ce21),
    .q21(cipher_0_ssbox_q21),
    .address22(cipher_0_ssbox_address22),
    .ce22(cipher_0_ssbox_ce22),
    .q22(cipher_0_ssbox_q22),
    .address23(cipher_0_ssbox_address23),
    .ce23(cipher_0_ssbox_ce23),
    .q23(cipher_0_ssbox_q23),
    .address24(cipher_0_ssbox_address24),
    .ce24(cipher_0_ssbox_ce24),
    .q24(cipher_0_ssbox_q24),
    .address25(cipher_0_ssbox_address25),
    .ce25(cipher_0_ssbox_ce25),
    .q25(cipher_0_ssbox_q25),
    .address26(cipher_0_ssbox_address26),
    .ce26(cipher_0_ssbox_ce26),
    .q26(cipher_0_ssbox_q26),
    .address27(cipher_0_ssbox_address27),
    .ce27(cipher_0_ssbox_ce27),
    .q27(cipher_0_ssbox_q27),
    .address28(cipher_0_ssbox_address28),
    .ce28(cipher_0_ssbox_ce28),
    .q28(cipher_0_ssbox_q28),
    .address29(cipher_0_ssbox_address29),
    .ce29(cipher_0_ssbox_ce29),
    .q29(cipher_0_ssbox_q29),
    .address30(cipher_0_ssbox_address30),
    .ce30(cipher_0_ssbox_ce30),
    .q30(cipher_0_ssbox_q30),
    .address31(cipher_0_ssbox_address31),
    .ce31(cipher_0_ssbox_ce31),
    .q31(cipher_0_ssbox_q31),
    .address32(cipher_0_ssbox_address32),
    .ce32(cipher_0_ssbox_ce32),
    .q32(cipher_0_ssbox_q32),
    .address33(cipher_0_ssbox_address33),
    .ce33(cipher_0_ssbox_ce33),
    .q33(cipher_0_ssbox_q33),
    .address34(cipher_0_ssbox_address34),
    .ce34(cipher_0_ssbox_ce34),
    .q34(cipher_0_ssbox_q34),
    .address35(cipher_0_ssbox_address35),
    .ce35(cipher_0_ssbox_ce35),
    .q35(cipher_0_ssbox_q35),
    .address36(cipher_0_ssbox_address36),
    .ce36(cipher_0_ssbox_ce36),
    .q36(cipher_0_ssbox_q36),
    .address37(cipher_0_ssbox_address37),
    .ce37(cipher_0_ssbox_ce37),
    .q37(cipher_0_ssbox_q37),
    .address38(cipher_0_ssbox_address38),
    .ce38(cipher_0_ssbox_ce38),
    .q38(cipher_0_ssbox_q38),
    .address39(cipher_0_ssbox_address39),
    .ce39(cipher_0_ssbox_ce39),
    .q39(cipher_0_ssbox_q39),
    .address40(cipher_0_ssbox_address40),
    .ce40(cipher_0_ssbox_ce40),
    .q40(cipher_0_ssbox_q40),
    .address41(cipher_0_ssbox_address41),
    .ce41(cipher_0_ssbox_ce41),
    .q41(cipher_0_ssbox_q41),
    .address42(cipher_0_ssbox_address42),
    .ce42(cipher_0_ssbox_ce42),
    .q42(cipher_0_ssbox_q42),
    .address43(cipher_0_ssbox_address43),
    .ce43(cipher_0_ssbox_ce43),
    .q43(cipher_0_ssbox_q43),
    .address44(cipher_0_ssbox_address44),
    .ce44(cipher_0_ssbox_ce44),
    .q44(cipher_0_ssbox_q44),
    .address45(cipher_0_ssbox_address45),
    .ce45(cipher_0_ssbox_ce45),
    .q45(cipher_0_ssbox_q45),
    .address46(cipher_0_ssbox_address46),
    .ce46(cipher_0_ssbox_ce46),
    .q46(cipher_0_ssbox_q46),
    .address47(cipher_0_ssbox_address47),
    .ce47(cipher_0_ssbox_ce47),
    .q47(cipher_0_ssbox_q47),
    .address48(cipher_0_ssbox_address48),
    .ce48(cipher_0_ssbox_ce48),
    .q48(cipher_0_ssbox_q48),
    .address49(cipher_0_ssbox_address49),
    .ce49(cipher_0_ssbox_ce49),
    .q49(cipher_0_ssbox_q49),
    .address50(cipher_0_ssbox_address50),
    .ce50(cipher_0_ssbox_ce50),
    .q50(cipher_0_ssbox_q50),
    .address51(cipher_0_ssbox_address51),
    .ce51(cipher_0_ssbox_ce51),
    .q51(cipher_0_ssbox_q51),
    .address52(cipher_0_ssbox_address52),
    .ce52(cipher_0_ssbox_ce52),
    .q52(cipher_0_ssbox_q52),
    .address53(cipher_0_ssbox_address53),
    .ce53(cipher_0_ssbox_ce53),
    .q53(cipher_0_ssbox_q53),
    .address54(cipher_0_ssbox_address54),
    .ce54(cipher_0_ssbox_ce54),
    .q54(cipher_0_ssbox_q54),
    .address55(cipher_0_ssbox_address55),
    .ce55(cipher_0_ssbox_ce55),
    .q55(cipher_0_ssbox_q55),
    .address56(cipher_0_ssbox_address56),
    .ce56(cipher_0_ssbox_ce56),
    .q56(cipher_0_ssbox_q56),
    .address57(cipher_0_ssbox_address57),
    .ce57(cipher_0_ssbox_ce57),
    .q57(cipher_0_ssbox_q57),
    .address58(cipher_0_ssbox_address58),
    .ce58(cipher_0_ssbox_ce58),
    .q58(cipher_0_ssbox_q58),
    .address59(cipher_0_ssbox_address59),
    .ce59(cipher_0_ssbox_ce59),
    .q59(cipher_0_ssbox_q59),
    .address60(cipher_0_ssbox_address60),
    .ce60(cipher_0_ssbox_ce60),
    .q60(cipher_0_ssbox_q60),
    .address61(cipher_0_ssbox_address61),
    .ce61(cipher_0_ssbox_ce61),
    .q61(cipher_0_ssbox_q61),
    .address62(cipher_0_ssbox_address62),
    .ce62(cipher_0_ssbox_ce62),
    .q62(cipher_0_ssbox_q62),
    .address63(cipher_0_ssbox_address63),
    .ce63(cipher_0_ssbox_ce63),
    .q63(cipher_0_ssbox_q63),
    .address64(cipher_0_ssbox_address64),
    .ce64(cipher_0_ssbox_ce64),
    .q64(cipher_0_ssbox_q64),
    .address65(cipher_0_ssbox_address65),
    .ce65(cipher_0_ssbox_ce65),
    .q65(cipher_0_ssbox_q65),
    .address66(cipher_0_ssbox_address66),
    .ce66(cipher_0_ssbox_ce66),
    .q66(cipher_0_ssbox_q66),
    .address67(cipher_0_ssbox_address67),
    .ce67(cipher_0_ssbox_ce67),
    .q67(cipher_0_ssbox_q67),
    .address68(cipher_0_ssbox_address68),
    .ce68(cipher_0_ssbox_ce68),
    .q68(cipher_0_ssbox_q68),
    .address69(cipher_0_ssbox_address69),
    .ce69(cipher_0_ssbox_ce69),
    .q69(cipher_0_ssbox_q69),
    .address70(cipher_0_ssbox_address70),
    .ce70(cipher_0_ssbox_ce70),
    .q70(cipher_0_ssbox_q70),
    .address71(cipher_0_ssbox_address71),
    .ce71(cipher_0_ssbox_ce71),
    .q71(cipher_0_ssbox_q71),
    .address72(cipher_0_ssbox_address72),
    .ce72(cipher_0_ssbox_ce72),
    .q72(cipher_0_ssbox_q72),
    .address73(cipher_0_ssbox_address73),
    .ce73(cipher_0_ssbox_ce73),
    .q73(cipher_0_ssbox_q73),
    .address74(cipher_0_ssbox_address74),
    .ce74(cipher_0_ssbox_ce74),
    .q74(cipher_0_ssbox_q74),
    .address75(cipher_0_ssbox_address75),
    .ce75(cipher_0_ssbox_ce75),
    .q75(cipher_0_ssbox_q75),
    .address76(cipher_0_ssbox_address76),
    .ce76(cipher_0_ssbox_ce76),
    .q76(cipher_0_ssbox_q76),
    .address77(cipher_0_ssbox_address77),
    .ce77(cipher_0_ssbox_ce77),
    .q77(cipher_0_ssbox_q77),
    .address78(cipher_0_ssbox_address78),
    .ce78(cipher_0_ssbox_ce78),
    .q78(cipher_0_ssbox_q78),
    .address79(cipher_0_ssbox_address79),
    .ce79(cipher_0_ssbox_ce79),
    .q79(cipher_0_ssbox_q79),
    .address80(cipher_0_ssbox_address80),
    .ce80(cipher_0_ssbox_ce80),
    .q80(cipher_0_ssbox_q80),
    .address81(cipher_0_ssbox_address81),
    .ce81(cipher_0_ssbox_ce81),
    .q81(cipher_0_ssbox_q81),
    .address82(cipher_0_ssbox_address82),
    .ce82(cipher_0_ssbox_ce82),
    .q82(cipher_0_ssbox_q82),
    .address83(cipher_0_ssbox_address83),
    .ce83(cipher_0_ssbox_ce83),
    .q83(cipher_0_ssbox_q83),
    .address84(cipher_0_ssbox_address84),
    .ce84(cipher_0_ssbox_ce84),
    .q84(cipher_0_ssbox_q84),
    .address85(cipher_0_ssbox_address85),
    .ce85(cipher_0_ssbox_ce85),
    .q85(cipher_0_ssbox_q85),
    .address86(cipher_0_ssbox_address86),
    .ce86(cipher_0_ssbox_ce86),
    .q86(cipher_0_ssbox_q86),
    .address87(cipher_0_ssbox_address87),
    .ce87(cipher_0_ssbox_ce87),
    .q87(cipher_0_ssbox_q87),
    .address88(cipher_0_ssbox_address88),
    .ce88(cipher_0_ssbox_ce88),
    .q88(cipher_0_ssbox_q88),
    .address89(cipher_0_ssbox_address89),
    .ce89(cipher_0_ssbox_ce89),
    .q89(cipher_0_ssbox_q89),
    .address90(cipher_0_ssbox_address90),
    .ce90(cipher_0_ssbox_ce90),
    .q90(cipher_0_ssbox_q90),
    .address91(cipher_0_ssbox_address91),
    .ce91(cipher_0_ssbox_ce91),
    .q91(cipher_0_ssbox_q91),
    .address92(cipher_0_ssbox_address92),
    .ce92(cipher_0_ssbox_ce92),
    .q92(cipher_0_ssbox_q92),
    .address93(cipher_0_ssbox_address93),
    .ce93(cipher_0_ssbox_ce93),
    .q93(cipher_0_ssbox_q93),
    .address94(cipher_0_ssbox_address94),
    .ce94(cipher_0_ssbox_ce94),
    .q94(cipher_0_ssbox_q94),
    .address95(cipher_0_ssbox_address95),
    .ce95(cipher_0_ssbox_ce95),
    .q95(cipher_0_ssbox_q95),
    .address96(cipher_0_ssbox_address96),
    .ce96(cipher_0_ssbox_ce96),
    .q96(cipher_0_ssbox_q96),
    .address97(cipher_0_ssbox_address97),
    .ce97(cipher_0_ssbox_ce97),
    .q97(cipher_0_ssbox_q97),
    .address98(cipher_0_ssbox_address98),
    .ce98(cipher_0_ssbox_ce98),
    .q98(cipher_0_ssbox_q98),
    .address99(cipher_0_ssbox_address99),
    .ce99(cipher_0_ssbox_ce99),
    .q99(cipher_0_ssbox_q99),
    .address100(cipher_0_ssbox_address100),
    .ce100(cipher_0_ssbox_ce100),
    .q100(cipher_0_ssbox_q100),
    .address101(cipher_0_ssbox_address101),
    .ce101(cipher_0_ssbox_ce101),
    .q101(cipher_0_ssbox_q101),
    .address102(cipher_0_ssbox_address102),
    .ce102(cipher_0_ssbox_ce102),
    .q102(cipher_0_ssbox_q102),
    .address103(cipher_0_ssbox_address103),
    .ce103(cipher_0_ssbox_ce103),
    .q103(cipher_0_ssbox_q103),
    .address104(cipher_0_ssbox_address104),
    .ce104(cipher_0_ssbox_ce104),
    .q104(cipher_0_ssbox_q104),
    .address105(cipher_0_ssbox_address105),
    .ce105(cipher_0_ssbox_ce105),
    .q105(cipher_0_ssbox_q105),
    .address106(cipher_0_ssbox_address106),
    .ce106(cipher_0_ssbox_ce106),
    .q106(cipher_0_ssbox_q106),
    .address107(cipher_0_ssbox_address107),
    .ce107(cipher_0_ssbox_ce107),
    .q107(cipher_0_ssbox_q107),
    .address108(cipher_0_ssbox_address108),
    .ce108(cipher_0_ssbox_ce108),
    .q108(cipher_0_ssbox_q108),
    .address109(cipher_0_ssbox_address109),
    .ce109(cipher_0_ssbox_ce109),
    .q109(cipher_0_ssbox_q109),
    .address110(cipher_0_ssbox_address110),
    .ce110(cipher_0_ssbox_ce110),
    .q110(cipher_0_ssbox_q110),
    .address111(cipher_0_ssbox_address111),
    .ce111(cipher_0_ssbox_ce111),
    .q111(cipher_0_ssbox_q111),
    .address112(cipher_0_ssbox_address112),
    .ce112(cipher_0_ssbox_ce112),
    .q112(cipher_0_ssbox_q112),
    .address113(cipher_0_ssbox_address113),
    .ce113(cipher_0_ssbox_ce113),
    .q113(cipher_0_ssbox_q113),
    .address114(cipher_0_ssbox_address114),
    .ce114(cipher_0_ssbox_ce114),
    .q114(cipher_0_ssbox_q114),
    .address115(cipher_0_ssbox_address115),
    .ce115(cipher_0_ssbox_ce115),
    .q115(cipher_0_ssbox_q115),
    .address116(cipher_0_ssbox_address116),
    .ce116(cipher_0_ssbox_ce116),
    .q116(cipher_0_ssbox_q116),
    .address117(cipher_0_ssbox_address117),
    .ce117(cipher_0_ssbox_ce117),
    .q117(cipher_0_ssbox_q117),
    .address118(cipher_0_ssbox_address118),
    .ce118(cipher_0_ssbox_ce118),
    .q118(cipher_0_ssbox_q118),
    .address119(cipher_0_ssbox_address119),
    .ce119(cipher_0_ssbox_ce119),
    .q119(cipher_0_ssbox_q119),
    .address120(cipher_0_ssbox_address120),
    .ce120(cipher_0_ssbox_ce120),
    .q120(cipher_0_ssbox_q120),
    .address121(cipher_0_ssbox_address121),
    .ce121(cipher_0_ssbox_ce121),
    .q121(cipher_0_ssbox_q121),
    .address122(cipher_0_ssbox_address122),
    .ce122(cipher_0_ssbox_ce122),
    .q122(cipher_0_ssbox_q122),
    .address123(cipher_0_ssbox_address123),
    .ce123(cipher_0_ssbox_ce123),
    .q123(cipher_0_ssbox_q123),
    .address124(cipher_0_ssbox_address124),
    .ce124(cipher_0_ssbox_ce124),
    .q124(cipher_0_ssbox_q124),
    .address125(cipher_0_ssbox_address125),
    .ce125(cipher_0_ssbox_ce125),
    .q125(cipher_0_ssbox_q125),
    .address126(cipher_0_ssbox_address126),
    .ce126(cipher_0_ssbox_ce126),
    .q126(cipher_0_ssbox_q126),
    .address127(cipher_0_ssbox_address127),
    .ce127(cipher_0_ssbox_ce127),
    .q127(cipher_0_ssbox_q127),
    .address128(cipher_0_ssbox_address128),
    .ce128(cipher_0_ssbox_ce128),
    .q128(cipher_0_ssbox_q128),
    .address129(cipher_0_ssbox_address129),
    .ce129(cipher_0_ssbox_ce129),
    .q129(cipher_0_ssbox_q129),
    .address130(cipher_0_ssbox_address130),
    .ce130(cipher_0_ssbox_ce130),
    .q130(cipher_0_ssbox_q130),
    .address131(cipher_0_ssbox_address131),
    .ce131(cipher_0_ssbox_ce131),
    .q131(cipher_0_ssbox_q131),
    .address132(cipher_0_ssbox_address132),
    .ce132(cipher_0_ssbox_ce132),
    .q132(cipher_0_ssbox_q132),
    .address133(cipher_0_ssbox_address133),
    .ce133(cipher_0_ssbox_ce133),
    .q133(cipher_0_ssbox_q133),
    .address134(cipher_0_ssbox_address134),
    .ce134(cipher_0_ssbox_ce134),
    .q134(cipher_0_ssbox_q134),
    .address135(cipher_0_ssbox_address135),
    .ce135(cipher_0_ssbox_ce135),
    .q135(cipher_0_ssbox_q135),
    .address136(cipher_0_ssbox_address136),
    .ce136(cipher_0_ssbox_ce136),
    .q136(cipher_0_ssbox_q136),
    .address137(cipher_0_ssbox_address137),
    .ce137(cipher_0_ssbox_ce137),
    .q137(cipher_0_ssbox_q137),
    .address138(cipher_0_ssbox_address138),
    .ce138(cipher_0_ssbox_ce138),
    .q138(cipher_0_ssbox_q138),
    .address139(cipher_0_ssbox_address139),
    .ce139(cipher_0_ssbox_ce139),
    .q139(cipher_0_ssbox_q139),
    .address140(cipher_0_ssbox_address140),
    .ce140(cipher_0_ssbox_ce140),
    .q140(cipher_0_ssbox_q140),
    .address141(cipher_0_ssbox_address141),
    .ce141(cipher_0_ssbox_ce141),
    .q141(cipher_0_ssbox_q141),
    .address142(cipher_0_ssbox_address142),
    .ce142(cipher_0_ssbox_ce142),
    .q142(cipher_0_ssbox_q142),
    .address143(cipher_0_ssbox_address143),
    .ce143(cipher_0_ssbox_ce143),
    .q143(cipher_0_ssbox_q143),
    .address144(cipher_0_ssbox_address144),
    .ce144(cipher_0_ssbox_ce144),
    .q144(cipher_0_ssbox_q144),
    .address145(cipher_0_ssbox_address145),
    .ce145(cipher_0_ssbox_ce145),
    .q145(cipher_0_ssbox_q145),
    .address146(cipher_0_ssbox_address146),
    .ce146(cipher_0_ssbox_ce146),
    .q146(cipher_0_ssbox_q146),
    .address147(cipher_0_ssbox_address147),
    .ce147(cipher_0_ssbox_ce147),
    .q147(cipher_0_ssbox_q147),
    .address148(cipher_0_ssbox_address148),
    .ce148(cipher_0_ssbox_ce148),
    .q148(cipher_0_ssbox_q148),
    .address149(cipher_0_ssbox_address149),
    .ce149(cipher_0_ssbox_ce149),
    .q149(cipher_0_ssbox_q149),
    .address150(cipher_0_ssbox_address150),
    .ce150(cipher_0_ssbox_ce150),
    .q150(cipher_0_ssbox_q150),
    .address151(cipher_0_ssbox_address151),
    .ce151(cipher_0_ssbox_ce151),
    .q151(cipher_0_ssbox_q151),
    .address152(cipher_0_ssbox_address152),
    .ce152(cipher_0_ssbox_ce152),
    .q152(cipher_0_ssbox_q152),
    .address153(cipher_0_ssbox_address153),
    .ce153(cipher_0_ssbox_ce153),
    .q153(cipher_0_ssbox_q153),
    .address154(cipher_0_ssbox_address154),
    .ce154(cipher_0_ssbox_ce154),
    .q154(cipher_0_ssbox_q154),
    .address155(cipher_0_ssbox_address155),
    .ce155(cipher_0_ssbox_ce155),
    .q155(cipher_0_ssbox_q155),
    .address156(cipher_0_ssbox_address156),
    .ce156(cipher_0_ssbox_ce156),
    .q156(cipher_0_ssbox_q156),
    .address157(cipher_0_ssbox_address157),
    .ce157(cipher_0_ssbox_ce157),
    .q157(cipher_0_ssbox_q157),
    .address158(cipher_0_ssbox_address158),
    .ce158(cipher_0_ssbox_ce158),
    .q158(cipher_0_ssbox_q158),
    .address159(cipher_0_ssbox_address159),
    .ce159(cipher_0_ssbox_ce159),
    .q159(cipher_0_ssbox_q159)
);

testEnc_process_r_cipher_0_p16box_ROM_NP_LUTRAM_1R #(
    .DataWidth( 16 ),
    .AddressRange( 256 ),
    .AddressWidth( 8 ))
cipher_0_p16box_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(cipher_0_p16box_address0),
    .ce0(cipher_0_p16box_ce0),
    .q0(cipher_0_p16box_q0),
    .address1(cipher_0_p16box_address1),
    .ce1(cipher_0_p16box_ce1),
    .q1(cipher_0_p16box_q1),
    .address2(cipher_0_p16box_address2),
    .ce2(cipher_0_p16box_ce2),
    .q2(cipher_0_p16box_q2),
    .address3(cipher_0_p16box_address3),
    .ce3(cipher_0_p16box_ce3),
    .q3(cipher_0_p16box_q3),
    .address4(cipher_0_p16box_address4),
    .ce4(cipher_0_p16box_ce4),
    .q4(cipher_0_p16box_q4),
    .address5(cipher_0_p16box_address5),
    .ce5(cipher_0_p16box_ce5),
    .q5(cipher_0_p16box_q5),
    .address6(cipher_0_p16box_address6),
    .ce6(cipher_0_p16box_ce6),
    .q6(cipher_0_p16box_q6),
    .address7(cipher_0_p16box_address7),
    .ce7(cipher_0_p16box_ce7),
    .q7(cipher_0_p16box_q7),
    .address8(cipher_0_p16box_address8),
    .ce8(cipher_0_p16box_ce8),
    .q8(cipher_0_p16box_q8),
    .address9(cipher_0_p16box_address9),
    .ce9(cipher_0_p16box_ce9),
    .q9(cipher_0_p16box_q9),
    .address10(cipher_0_p16box_address10),
    .ce10(cipher_0_p16box_ce10),
    .q10(cipher_0_p16box_q10),
    .address11(cipher_0_p16box_address11),
    .ce11(cipher_0_p16box_ce11),
    .q11(cipher_0_p16box_q11),
    .address12(cipher_0_p16box_address12),
    .ce12(cipher_0_p16box_ce12),
    .q12(cipher_0_p16box_q12),
    .address13(cipher_0_p16box_address13),
    .ce13(cipher_0_p16box_ce13),
    .q13(cipher_0_p16box_q13),
    .address14(cipher_0_p16box_address14),
    .ce14(cipher_0_p16box_ce14),
    .q14(cipher_0_p16box_q14),
    .address15(cipher_0_p16box_address15),
    .ce15(cipher_0_p16box_ce15),
    .q15(cipher_0_p16box_q15),
    .address16(cipher_0_p16box_address16),
    .ce16(cipher_0_p16box_ce16),
    .q16(cipher_0_p16box_q16),
    .address17(cipher_0_p16box_address17),
    .ce17(cipher_0_p16box_ce17),
    .q17(cipher_0_p16box_q17),
    .address18(cipher_0_p16box_address18),
    .ce18(cipher_0_p16box_ce18),
    .q18(cipher_0_p16box_q18),
    .address19(cipher_0_p16box_address19),
    .ce19(cipher_0_p16box_ce19),
    .q19(cipher_0_p16box_q19),
    .address20(cipher_0_p16box_address20),
    .ce20(cipher_0_p16box_ce20),
    .q20(cipher_0_p16box_q20),
    .address21(cipher_0_p16box_address21),
    .ce21(cipher_0_p16box_ce21),
    .q21(cipher_0_p16box_q21),
    .address22(cipher_0_p16box_address22),
    .ce22(cipher_0_p16box_ce22),
    .q22(cipher_0_p16box_q22),
    .address23(cipher_0_p16box_address23),
    .ce23(cipher_0_p16box_ce23),
    .q23(cipher_0_p16box_q23),
    .address24(cipher_0_p16box_address24),
    .ce24(cipher_0_p16box_ce24),
    .q24(cipher_0_p16box_q24),
    .address25(cipher_0_p16box_address25),
    .ce25(cipher_0_p16box_ce25),
    .q25(cipher_0_p16box_q25),
    .address26(cipher_0_p16box_address26),
    .ce26(cipher_0_p16box_ce26),
    .q26(cipher_0_p16box_q26),
    .address27(cipher_0_p16box_address27),
    .ce27(cipher_0_p16box_ce27),
    .q27(cipher_0_p16box_q27),
    .address28(cipher_0_p16box_address28),
    .ce28(cipher_0_p16box_ce28),
    .q28(cipher_0_p16box_q28),
    .address29(cipher_0_p16box_address29),
    .ce29(cipher_0_p16box_ce29),
    .q29(cipher_0_p16box_q29),
    .address30(cipher_0_p16box_address30),
    .ce30(cipher_0_p16box_ce30),
    .q30(cipher_0_p16box_q30),
    .address31(cipher_0_p16box_address31),
    .ce31(cipher_0_p16box_ce31),
    .q31(cipher_0_p16box_q31),
    .address32(cipher_0_p16box_address32),
    .ce32(cipher_0_p16box_ce32),
    .q32(cipher_0_p16box_q32),
    .address33(cipher_0_p16box_address33),
    .ce33(cipher_0_p16box_ce33),
    .q33(cipher_0_p16box_q33),
    .address34(cipher_0_p16box_address34),
    .ce34(cipher_0_p16box_ce34),
    .q34(cipher_0_p16box_q34),
    .address35(cipher_0_p16box_address35),
    .ce35(cipher_0_p16box_ce35),
    .q35(cipher_0_p16box_q35),
    .address36(cipher_0_p16box_address36),
    .ce36(cipher_0_p16box_ce36),
    .q36(cipher_0_p16box_q36),
    .address37(cipher_0_p16box_address37),
    .ce37(cipher_0_p16box_ce37),
    .q37(cipher_0_p16box_q37),
    .address38(cipher_0_p16box_address38),
    .ce38(cipher_0_p16box_ce38),
    .q38(cipher_0_p16box_q38),
    .address39(cipher_0_p16box_address39),
    .ce39(cipher_0_p16box_ce39),
    .q39(cipher_0_p16box_q39),
    .address40(cipher_0_p16box_address40),
    .ce40(cipher_0_p16box_ce40),
    .q40(cipher_0_p16box_q40),
    .address41(cipher_0_p16box_address41),
    .ce41(cipher_0_p16box_ce41),
    .q41(cipher_0_p16box_q41),
    .address42(cipher_0_p16box_address42),
    .ce42(cipher_0_p16box_ce42),
    .q42(cipher_0_p16box_q42),
    .address43(cipher_0_p16box_address43),
    .ce43(cipher_0_p16box_ce43),
    .q43(cipher_0_p16box_q43),
    .address44(cipher_0_p16box_address44),
    .ce44(cipher_0_p16box_ce44),
    .q44(cipher_0_p16box_q44),
    .address45(cipher_0_p16box_address45),
    .ce45(cipher_0_p16box_ce45),
    .q45(cipher_0_p16box_q45),
    .address46(cipher_0_p16box_address46),
    .ce46(cipher_0_p16box_ce46),
    .q46(cipher_0_p16box_q46),
    .address47(cipher_0_p16box_address47),
    .ce47(cipher_0_p16box_ce47),
    .q47(cipher_0_p16box_q47),
    .address48(cipher_0_p16box_address48),
    .ce48(cipher_0_p16box_ce48),
    .q48(cipher_0_p16box_q48),
    .address49(cipher_0_p16box_address49),
    .ce49(cipher_0_p16box_ce49),
    .q49(cipher_0_p16box_q49),
    .address50(cipher_0_p16box_address50),
    .ce50(cipher_0_p16box_ce50),
    .q50(cipher_0_p16box_q50),
    .address51(cipher_0_p16box_address51),
    .ce51(cipher_0_p16box_ce51),
    .q51(cipher_0_p16box_q51),
    .address52(cipher_0_p16box_address52),
    .ce52(cipher_0_p16box_ce52),
    .q52(cipher_0_p16box_q52),
    .address53(cipher_0_p16box_address53),
    .ce53(cipher_0_p16box_ce53),
    .q53(cipher_0_p16box_q53),
    .address54(cipher_0_p16box_address54),
    .ce54(cipher_0_p16box_ce54),
    .q54(cipher_0_p16box_q54),
    .address55(cipher_0_p16box_address55),
    .ce55(cipher_0_p16box_ce55),
    .q55(cipher_0_p16box_q55),
    .address56(cipher_0_p16box_address56),
    .ce56(cipher_0_p16box_ce56),
    .q56(cipher_0_p16box_q56),
    .address57(cipher_0_p16box_address57),
    .ce57(cipher_0_p16box_ce57),
    .q57(cipher_0_p16box_q57),
    .address58(cipher_0_p16box_address58),
    .ce58(cipher_0_p16box_ce58),
    .q58(cipher_0_p16box_q58),
    .address59(cipher_0_p16box_address59),
    .ce59(cipher_0_p16box_ce59),
    .q59(cipher_0_p16box_q59),
    .address60(cipher_0_p16box_address60),
    .ce60(cipher_0_p16box_ce60),
    .q60(cipher_0_p16box_q60),
    .address61(cipher_0_p16box_address61),
    .ce61(cipher_0_p16box_ce61),
    .q61(cipher_0_p16box_q61),
    .address62(cipher_0_p16box_address62),
    .ce62(cipher_0_p16box_ce62),
    .q62(cipher_0_p16box_q62),
    .address63(cipher_0_p16box_address63),
    .ce63(cipher_0_p16box_ce63),
    .q63(cipher_0_p16box_q63),
    .address64(cipher_0_p16box_address64),
    .ce64(cipher_0_p16box_ce64),
    .q64(cipher_0_p16box_q64),
    .address65(cipher_0_p16box_address65),
    .ce65(cipher_0_p16box_ce65),
    .q65(cipher_0_p16box_q65),
    .address66(cipher_0_p16box_address66),
    .ce66(cipher_0_p16box_ce66),
    .q66(cipher_0_p16box_q66),
    .address67(cipher_0_p16box_address67),
    .ce67(cipher_0_p16box_ce67),
    .q67(cipher_0_p16box_q67),
    .address68(cipher_0_p16box_address68),
    .ce68(cipher_0_p16box_ce68),
    .q68(cipher_0_p16box_q68),
    .address69(cipher_0_p16box_address69),
    .ce69(cipher_0_p16box_ce69),
    .q69(cipher_0_p16box_q69),
    .address70(cipher_0_p16box_address70),
    .ce70(cipher_0_p16box_ce70),
    .q70(cipher_0_p16box_q70),
    .address71(cipher_0_p16box_address71),
    .ce71(cipher_0_p16box_ce71),
    .q71(cipher_0_p16box_q71),
    .address72(cipher_0_p16box_address72),
    .ce72(cipher_0_p16box_ce72),
    .q72(cipher_0_p16box_q72),
    .address73(cipher_0_p16box_address73),
    .ce73(cipher_0_p16box_ce73),
    .q73(cipher_0_p16box_q73),
    .address74(cipher_0_p16box_address74),
    .ce74(cipher_0_p16box_ce74),
    .q74(cipher_0_p16box_q74),
    .address75(cipher_0_p16box_address75),
    .ce75(cipher_0_p16box_ce75),
    .q75(cipher_0_p16box_q75),
    .address76(cipher_0_p16box_address76),
    .ce76(cipher_0_p16box_ce76),
    .q76(cipher_0_p16box_q76),
    .address77(cipher_0_p16box_address77),
    .ce77(cipher_0_p16box_ce77),
    .q77(cipher_0_p16box_q77),
    .address78(cipher_0_p16box_address78),
    .ce78(cipher_0_p16box_ce78),
    .q78(cipher_0_p16box_q78),
    .address79(cipher_0_p16box_address79),
    .ce79(cipher_0_p16box_ce79),
    .q79(cipher_0_p16box_q79),
    .address80(cipher_0_p16box_address80),
    .ce80(cipher_0_p16box_ce80),
    .q80(cipher_0_p16box_q80),
    .address81(cipher_0_p16box_address81),
    .ce81(cipher_0_p16box_ce81),
    .q81(cipher_0_p16box_q81),
    .address82(cipher_0_p16box_address82),
    .ce82(cipher_0_p16box_ce82),
    .q82(cipher_0_p16box_q82),
    .address83(cipher_0_p16box_address83),
    .ce83(cipher_0_p16box_ce83),
    .q83(cipher_0_p16box_q83),
    .address84(cipher_0_p16box_address84),
    .ce84(cipher_0_p16box_ce84),
    .q84(cipher_0_p16box_q84),
    .address85(cipher_0_p16box_address85),
    .ce85(cipher_0_p16box_ce85),
    .q85(cipher_0_p16box_q85),
    .address86(cipher_0_p16box_address86),
    .ce86(cipher_0_p16box_ce86),
    .q86(cipher_0_p16box_q86),
    .address87(cipher_0_p16box_address87),
    .ce87(cipher_0_p16box_ce87),
    .q87(cipher_0_p16box_q87),
    .address88(cipher_0_p16box_address88),
    .ce88(cipher_0_p16box_ce88),
    .q88(cipher_0_p16box_q88),
    .address89(cipher_0_p16box_address89),
    .ce89(cipher_0_p16box_ce89),
    .q89(cipher_0_p16box_q89),
    .address90(cipher_0_p16box_address90),
    .ce90(cipher_0_p16box_ce90),
    .q90(cipher_0_p16box_q90),
    .address91(cipher_0_p16box_address91),
    .ce91(cipher_0_p16box_ce91),
    .q91(cipher_0_p16box_q91),
    .address92(cipher_0_p16box_address92),
    .ce92(cipher_0_p16box_ce92),
    .q92(cipher_0_p16box_q92),
    .address93(cipher_0_p16box_address93),
    .ce93(cipher_0_p16box_ce93),
    .q93(cipher_0_p16box_q93),
    .address94(cipher_0_p16box_address94),
    .ce94(cipher_0_p16box_ce94),
    .q94(cipher_0_p16box_q94),
    .address95(cipher_0_p16box_address95),
    .ce95(cipher_0_p16box_ce95),
    .q95(cipher_0_p16box_q95),
    .address96(cipher_0_p16box_address96),
    .ce96(cipher_0_p16box_ce96),
    .q96(cipher_0_p16box_q96),
    .address97(cipher_0_p16box_address97),
    .ce97(cipher_0_p16box_ce97),
    .q97(cipher_0_p16box_q97),
    .address98(cipher_0_p16box_address98),
    .ce98(cipher_0_p16box_ce98),
    .q98(cipher_0_p16box_q98),
    .address99(cipher_0_p16box_address99),
    .ce99(cipher_0_p16box_ce99),
    .q99(cipher_0_p16box_q99),
    .address100(cipher_0_p16box_address100),
    .ce100(cipher_0_p16box_ce100),
    .q100(cipher_0_p16box_q100),
    .address101(cipher_0_p16box_address101),
    .ce101(cipher_0_p16box_ce101),
    .q101(cipher_0_p16box_q101),
    .address102(cipher_0_p16box_address102),
    .ce102(cipher_0_p16box_ce102),
    .q102(cipher_0_p16box_q102),
    .address103(cipher_0_p16box_address103),
    .ce103(cipher_0_p16box_ce103),
    .q103(cipher_0_p16box_q103),
    .address104(cipher_0_p16box_address104),
    .ce104(cipher_0_p16box_ce104),
    .q104(cipher_0_p16box_q104),
    .address105(cipher_0_p16box_address105),
    .ce105(cipher_0_p16box_ce105),
    .q105(cipher_0_p16box_q105),
    .address106(cipher_0_p16box_address106),
    .ce106(cipher_0_p16box_ce106),
    .q106(cipher_0_p16box_q106),
    .address107(cipher_0_p16box_address107),
    .ce107(cipher_0_p16box_ce107),
    .q107(cipher_0_p16box_q107),
    .address108(cipher_0_p16box_address108),
    .ce108(cipher_0_p16box_ce108),
    .q108(cipher_0_p16box_q108),
    .address109(cipher_0_p16box_address109),
    .ce109(cipher_0_p16box_ce109),
    .q109(cipher_0_p16box_q109),
    .address110(cipher_0_p16box_address110),
    .ce110(cipher_0_p16box_ce110),
    .q110(cipher_0_p16box_q110),
    .address111(cipher_0_p16box_address111),
    .ce111(cipher_0_p16box_ce111),
    .q111(cipher_0_p16box_q111),
    .address112(cipher_0_p16box_address112),
    .ce112(cipher_0_p16box_ce112),
    .q112(cipher_0_p16box_q112),
    .address113(cipher_0_p16box_address113),
    .ce113(cipher_0_p16box_ce113),
    .q113(cipher_0_p16box_q113),
    .address114(cipher_0_p16box_address114),
    .ce114(cipher_0_p16box_ce114),
    .q114(cipher_0_p16box_q114),
    .address115(cipher_0_p16box_address115),
    .ce115(cipher_0_p16box_ce115),
    .q115(cipher_0_p16box_q115),
    .address116(cipher_0_p16box_address116),
    .ce116(cipher_0_p16box_ce116),
    .q116(cipher_0_p16box_q116),
    .address117(cipher_0_p16box_address117),
    .ce117(cipher_0_p16box_ce117),
    .q117(cipher_0_p16box_q117),
    .address118(cipher_0_p16box_address118),
    .ce118(cipher_0_p16box_ce118),
    .q118(cipher_0_p16box_q118),
    .address119(cipher_0_p16box_address119),
    .ce119(cipher_0_p16box_ce119),
    .q119(cipher_0_p16box_q119),
    .address120(cipher_0_p16box_address120),
    .ce120(cipher_0_p16box_ce120),
    .q120(cipher_0_p16box_q120),
    .address121(cipher_0_p16box_address121),
    .ce121(cipher_0_p16box_ce121),
    .q121(cipher_0_p16box_q121),
    .address122(cipher_0_p16box_address122),
    .ce122(cipher_0_p16box_ce122),
    .q122(cipher_0_p16box_q122),
    .address123(cipher_0_p16box_address123),
    .ce123(cipher_0_p16box_ce123),
    .q123(cipher_0_p16box_q123),
    .address124(cipher_0_p16box_address124),
    .ce124(cipher_0_p16box_ce124),
    .q124(cipher_0_p16box_q124),
    .address125(cipher_0_p16box_address125),
    .ce125(cipher_0_p16box_ce125),
    .q125(cipher_0_p16box_q125),
    .address126(cipher_0_p16box_address126),
    .ce126(cipher_0_p16box_ce126),
    .q126(cipher_0_p16box_q126),
    .address127(cipher_0_p16box_address127),
    .ce127(cipher_0_p16box_ce127),
    .q127(cipher_0_p16box_q127),
    .address128(cipher_0_p16box_address128),
    .ce128(cipher_0_p16box_ce128),
    .q128(cipher_0_p16box_q128),
    .address129(cipher_0_p16box_address129),
    .ce129(cipher_0_p16box_ce129),
    .q129(cipher_0_p16box_q129),
    .address130(cipher_0_p16box_address130),
    .ce130(cipher_0_p16box_ce130),
    .q130(cipher_0_p16box_q130),
    .address131(cipher_0_p16box_address131),
    .ce131(cipher_0_p16box_ce131),
    .q131(cipher_0_p16box_q131),
    .address132(cipher_0_p16box_address132),
    .ce132(cipher_0_p16box_ce132),
    .q132(cipher_0_p16box_q132),
    .address133(cipher_0_p16box_address133),
    .ce133(cipher_0_p16box_ce133),
    .q133(cipher_0_p16box_q133),
    .address134(cipher_0_p16box_address134),
    .ce134(cipher_0_p16box_ce134),
    .q134(cipher_0_p16box_q134),
    .address135(cipher_0_p16box_address135),
    .ce135(cipher_0_p16box_ce135),
    .q135(cipher_0_p16box_q135),
    .address136(cipher_0_p16box_address136),
    .ce136(cipher_0_p16box_ce136),
    .q136(cipher_0_p16box_q136),
    .address137(cipher_0_p16box_address137),
    .ce137(cipher_0_p16box_ce137),
    .q137(cipher_0_p16box_q137),
    .address138(cipher_0_p16box_address138),
    .ce138(cipher_0_p16box_ce138),
    .q138(cipher_0_p16box_q138),
    .address139(cipher_0_p16box_address139),
    .ce139(cipher_0_p16box_ce139),
    .q139(cipher_0_p16box_q139),
    .address140(cipher_0_p16box_address140),
    .ce140(cipher_0_p16box_ce140),
    .q140(cipher_0_p16box_q140),
    .address141(cipher_0_p16box_address141),
    .ce141(cipher_0_p16box_ce141),
    .q141(cipher_0_p16box_q141),
    .address142(cipher_0_p16box_address142),
    .ce142(cipher_0_p16box_ce142),
    .q142(cipher_0_p16box_q142),
    .address143(cipher_0_p16box_address143),
    .ce143(cipher_0_p16box_ce143),
    .q143(cipher_0_p16box_q143)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_enable_reg_pp0_iter1 <= ap_start;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter10 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter10 <= ap_enable_reg_pp0_iter9;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter11 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter11 <= ap_enable_reg_pp0_iter10;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter12 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter12 <= ap_enable_reg_pp0_iter11;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter13 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter13 <= ap_enable_reg_pp0_iter12;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter14 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter14 <= ap_enable_reg_pp0_iter13;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter15 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter15 <= ap_enable_reg_pp0_iter14;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter16 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter16 <= ap_enable_reg_pp0_iter15;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter17 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter17 <= ap_enable_reg_pp0_iter16;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter18 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter18 <= ap_enable_reg_pp0_iter17;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter19 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter19 <= ap_enable_reg_pp0_iter18;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter5 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter6 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter7 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter8 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter8 <= ap_enable_reg_pp0_iter7;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter9 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter9 <= ap_enable_reg_pp0_iter8;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        p_read_10_reg_11669 <= p_read1;
        p_read_10_reg_11669_pp0_iter1_reg <= p_read_10_reg_11669;
        p_read_1_reg_11624 <= p_read10;
        p_read_1_reg_11624_pp0_iter1_reg <= p_read_1_reg_11624;
        p_read_2_reg_11629 <= p_read9;
        p_read_2_reg_11629_pp0_iter1_reg <= p_read_2_reg_11629;
        p_read_3_reg_11634 <= p_read8;
        p_read_3_reg_11634_pp0_iter1_reg <= p_read_3_reg_11634;
        p_read_4_reg_11639 <= p_read7;
        p_read_4_reg_11639_pp0_iter1_reg <= p_read_4_reg_11639;
        p_read_5_reg_11644 <= p_read6;
        p_read_5_reg_11644_pp0_iter1_reg <= p_read_5_reg_11644;
        p_read_6_reg_11649 <= p_read5;
        p_read_6_reg_11649_pp0_iter1_reg <= p_read_6_reg_11649;
        p_read_7_reg_11654 <= p_read4;
        p_read_7_reg_11654_pp0_iter1_reg <= p_read_7_reg_11654;
        p_read_8_reg_11659 <= p_read3;
        p_read_8_reg_11659_pp0_iter1_reg <= p_read_8_reg_11659;
        p_read_9_reg_11664 <= p_read2;
        p_read_9_reg_11664_pp0_iter1_reg <= p_read_9_reg_11664;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        p_read_1_reg_11624_pp0_iter10_reg <= p_read_1_reg_11624_pp0_iter9_reg;
        p_read_1_reg_11624_pp0_iter11_reg <= p_read_1_reg_11624_pp0_iter10_reg;
        p_read_1_reg_11624_pp0_iter12_reg <= p_read_1_reg_11624_pp0_iter11_reg;
        p_read_1_reg_11624_pp0_iter13_reg <= p_read_1_reg_11624_pp0_iter12_reg;
        p_read_1_reg_11624_pp0_iter14_reg <= p_read_1_reg_11624_pp0_iter13_reg;
        p_read_1_reg_11624_pp0_iter15_reg <= p_read_1_reg_11624_pp0_iter14_reg;
        p_read_1_reg_11624_pp0_iter16_reg <= p_read_1_reg_11624_pp0_iter15_reg;
        p_read_1_reg_11624_pp0_iter17_reg <= p_read_1_reg_11624_pp0_iter16_reg;
        p_read_1_reg_11624_pp0_iter18_reg <= p_read_1_reg_11624_pp0_iter17_reg;
        p_read_1_reg_11624_pp0_iter2_reg <= p_read_1_reg_11624_pp0_iter1_reg;
        p_read_1_reg_11624_pp0_iter3_reg <= p_read_1_reg_11624_pp0_iter2_reg;
        p_read_1_reg_11624_pp0_iter4_reg <= p_read_1_reg_11624_pp0_iter3_reg;
        p_read_1_reg_11624_pp0_iter5_reg <= p_read_1_reg_11624_pp0_iter4_reg;
        p_read_1_reg_11624_pp0_iter6_reg <= p_read_1_reg_11624_pp0_iter5_reg;
        p_read_1_reg_11624_pp0_iter7_reg <= p_read_1_reg_11624_pp0_iter6_reg;
        p_read_1_reg_11624_pp0_iter8_reg <= p_read_1_reg_11624_pp0_iter7_reg;
        p_read_1_reg_11624_pp0_iter9_reg <= p_read_1_reg_11624_pp0_iter8_reg;
        p_read_2_reg_11629_pp0_iter10_reg <= p_read_2_reg_11629_pp0_iter9_reg;
        p_read_2_reg_11629_pp0_iter11_reg <= p_read_2_reg_11629_pp0_iter10_reg;
        p_read_2_reg_11629_pp0_iter12_reg <= p_read_2_reg_11629_pp0_iter11_reg;
        p_read_2_reg_11629_pp0_iter13_reg <= p_read_2_reg_11629_pp0_iter12_reg;
        p_read_2_reg_11629_pp0_iter14_reg <= p_read_2_reg_11629_pp0_iter13_reg;
        p_read_2_reg_11629_pp0_iter15_reg <= p_read_2_reg_11629_pp0_iter14_reg;
        p_read_2_reg_11629_pp0_iter16_reg <= p_read_2_reg_11629_pp0_iter15_reg;
        p_read_2_reg_11629_pp0_iter17_reg <= p_read_2_reg_11629_pp0_iter16_reg;
        p_read_2_reg_11629_pp0_iter2_reg <= p_read_2_reg_11629_pp0_iter1_reg;
        p_read_2_reg_11629_pp0_iter3_reg <= p_read_2_reg_11629_pp0_iter2_reg;
        p_read_2_reg_11629_pp0_iter4_reg <= p_read_2_reg_11629_pp0_iter3_reg;
        p_read_2_reg_11629_pp0_iter5_reg <= p_read_2_reg_11629_pp0_iter4_reg;
        p_read_2_reg_11629_pp0_iter6_reg <= p_read_2_reg_11629_pp0_iter5_reg;
        p_read_2_reg_11629_pp0_iter7_reg <= p_read_2_reg_11629_pp0_iter6_reg;
        p_read_2_reg_11629_pp0_iter8_reg <= p_read_2_reg_11629_pp0_iter7_reg;
        p_read_2_reg_11629_pp0_iter9_reg <= p_read_2_reg_11629_pp0_iter8_reg;
        p_read_3_reg_11634_pp0_iter10_reg <= p_read_3_reg_11634_pp0_iter9_reg;
        p_read_3_reg_11634_pp0_iter11_reg <= p_read_3_reg_11634_pp0_iter10_reg;
        p_read_3_reg_11634_pp0_iter12_reg <= p_read_3_reg_11634_pp0_iter11_reg;
        p_read_3_reg_11634_pp0_iter13_reg <= p_read_3_reg_11634_pp0_iter12_reg;
        p_read_3_reg_11634_pp0_iter14_reg <= p_read_3_reg_11634_pp0_iter13_reg;
        p_read_3_reg_11634_pp0_iter15_reg <= p_read_3_reg_11634_pp0_iter14_reg;
        p_read_3_reg_11634_pp0_iter2_reg <= p_read_3_reg_11634_pp0_iter1_reg;
        p_read_3_reg_11634_pp0_iter3_reg <= p_read_3_reg_11634_pp0_iter2_reg;
        p_read_3_reg_11634_pp0_iter4_reg <= p_read_3_reg_11634_pp0_iter3_reg;
        p_read_3_reg_11634_pp0_iter5_reg <= p_read_3_reg_11634_pp0_iter4_reg;
        p_read_3_reg_11634_pp0_iter6_reg <= p_read_3_reg_11634_pp0_iter5_reg;
        p_read_3_reg_11634_pp0_iter7_reg <= p_read_3_reg_11634_pp0_iter6_reg;
        p_read_3_reg_11634_pp0_iter8_reg <= p_read_3_reg_11634_pp0_iter7_reg;
        p_read_3_reg_11634_pp0_iter9_reg <= p_read_3_reg_11634_pp0_iter8_reg;
        p_read_4_reg_11639_pp0_iter10_reg <= p_read_4_reg_11639_pp0_iter9_reg;
        p_read_4_reg_11639_pp0_iter11_reg <= p_read_4_reg_11639_pp0_iter10_reg;
        p_read_4_reg_11639_pp0_iter12_reg <= p_read_4_reg_11639_pp0_iter11_reg;
        p_read_4_reg_11639_pp0_iter13_reg <= p_read_4_reg_11639_pp0_iter12_reg;
        p_read_4_reg_11639_pp0_iter2_reg <= p_read_4_reg_11639_pp0_iter1_reg;
        p_read_4_reg_11639_pp0_iter3_reg <= p_read_4_reg_11639_pp0_iter2_reg;
        p_read_4_reg_11639_pp0_iter4_reg <= p_read_4_reg_11639_pp0_iter3_reg;
        p_read_4_reg_11639_pp0_iter5_reg <= p_read_4_reg_11639_pp0_iter4_reg;
        p_read_4_reg_11639_pp0_iter6_reg <= p_read_4_reg_11639_pp0_iter5_reg;
        p_read_4_reg_11639_pp0_iter7_reg <= p_read_4_reg_11639_pp0_iter6_reg;
        p_read_4_reg_11639_pp0_iter8_reg <= p_read_4_reg_11639_pp0_iter7_reg;
        p_read_4_reg_11639_pp0_iter9_reg <= p_read_4_reg_11639_pp0_iter8_reg;
        p_read_5_reg_11644_pp0_iter10_reg <= p_read_5_reg_11644_pp0_iter9_reg;
        p_read_5_reg_11644_pp0_iter11_reg <= p_read_5_reg_11644_pp0_iter10_reg;
        p_read_5_reg_11644_pp0_iter2_reg <= p_read_5_reg_11644_pp0_iter1_reg;
        p_read_5_reg_11644_pp0_iter3_reg <= p_read_5_reg_11644_pp0_iter2_reg;
        p_read_5_reg_11644_pp0_iter4_reg <= p_read_5_reg_11644_pp0_iter3_reg;
        p_read_5_reg_11644_pp0_iter5_reg <= p_read_5_reg_11644_pp0_iter4_reg;
        p_read_5_reg_11644_pp0_iter6_reg <= p_read_5_reg_11644_pp0_iter5_reg;
        p_read_5_reg_11644_pp0_iter7_reg <= p_read_5_reg_11644_pp0_iter6_reg;
        p_read_5_reg_11644_pp0_iter8_reg <= p_read_5_reg_11644_pp0_iter7_reg;
        p_read_5_reg_11644_pp0_iter9_reg <= p_read_5_reg_11644_pp0_iter8_reg;
        p_read_6_reg_11649_pp0_iter2_reg <= p_read_6_reg_11649_pp0_iter1_reg;
        p_read_6_reg_11649_pp0_iter3_reg <= p_read_6_reg_11649_pp0_iter2_reg;
        p_read_6_reg_11649_pp0_iter4_reg <= p_read_6_reg_11649_pp0_iter3_reg;
        p_read_6_reg_11649_pp0_iter5_reg <= p_read_6_reg_11649_pp0_iter4_reg;
        p_read_6_reg_11649_pp0_iter6_reg <= p_read_6_reg_11649_pp0_iter5_reg;
        p_read_6_reg_11649_pp0_iter7_reg <= p_read_6_reg_11649_pp0_iter6_reg;
        p_read_6_reg_11649_pp0_iter8_reg <= p_read_6_reg_11649_pp0_iter7_reg;
        p_read_6_reg_11649_pp0_iter9_reg <= p_read_6_reg_11649_pp0_iter8_reg;
        p_read_7_reg_11654_pp0_iter2_reg <= p_read_7_reg_11654_pp0_iter1_reg;
        p_read_7_reg_11654_pp0_iter3_reg <= p_read_7_reg_11654_pp0_iter2_reg;
        p_read_7_reg_11654_pp0_iter4_reg <= p_read_7_reg_11654_pp0_iter3_reg;
        p_read_7_reg_11654_pp0_iter5_reg <= p_read_7_reg_11654_pp0_iter4_reg;
        p_read_7_reg_11654_pp0_iter6_reg <= p_read_7_reg_11654_pp0_iter5_reg;
        p_read_7_reg_11654_pp0_iter7_reg <= p_read_7_reg_11654_pp0_iter6_reg;
        p_read_8_reg_11659_pp0_iter2_reg <= p_read_8_reg_11659_pp0_iter1_reg;
        p_read_8_reg_11659_pp0_iter3_reg <= p_read_8_reg_11659_pp0_iter2_reg;
        p_read_8_reg_11659_pp0_iter4_reg <= p_read_8_reg_11659_pp0_iter3_reg;
        p_read_8_reg_11659_pp0_iter5_reg <= p_read_8_reg_11659_pp0_iter4_reg;
        p_read_9_reg_11664_pp0_iter2_reg <= p_read_9_reg_11664_pp0_iter1_reg;
        p_read_9_reg_11664_pp0_iter3_reg <= p_read_9_reg_11664_pp0_iter2_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        tmp_1_V_10_reg_11760 <= cipher_0_ssbox_q158;
        tmp_2_1_V_10_reg_11766 <= cipher_0_ssbox_q157;
        tmp_2_2_V_10_reg_11790 <= cipher_0_ssbox_q153;
        tmp_3_V_10_reg_11844 <= cipher_0_ssbox_q144;
        tmp_V_11_reg_11796 <= cipher_0_ssbox_q152;
        tmp_V_12_reg_11826 <= cipher_0_ssbox_q147;
        tmp_V_15_reg_11820 <= cipher_0_ssbox_q148;
        tmp_V_1_reg_11784 <= cipher_0_ssbox_q154;
        tmp_V_2_reg_11814 <= cipher_0_ssbox_q149;
        tmp_V_4_reg_11778 <= cipher_0_ssbox_q155;
        tmp_V_5_reg_11808 <= cipher_0_ssbox_q150;
        tmp_V_6_reg_11838 <= cipher_0_ssbox_q145;
        tmp_V_7_reg_11772 <= cipher_0_ssbox_q156;
        tmp_V_8_reg_11802 <= cipher_0_ssbox_q151;
        tmp_V_9_reg_11832 <= cipher_0_ssbox_q146;
        tmp_V_reg_11754 <= cipher_0_ssbox_q159;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        tmp_1_V_11_reg_12016 <= cipher_0_ssbox_q142;
        tmp_2_1_V_11_reg_12022 <= cipher_0_ssbox_q141;
        tmp_2_2_V_11_reg_12046 <= cipher_0_ssbox_q137;
        tmp_3_V_11_reg_12100 <= cipher_0_ssbox_q128;
        tmp_V_16_reg_12010 <= cipher_0_ssbox_q143;
        tmp_V_17_reg_12040 <= cipher_0_ssbox_q138;
        tmp_V_18_reg_12070 <= cipher_0_ssbox_q133;
        tmp_V_20_reg_12034 <= cipher_0_ssbox_q139;
        tmp_V_21_reg_12064 <= cipher_0_ssbox_q134;
        tmp_V_22_reg_12094 <= cipher_0_ssbox_q129;
        tmp_V_23_reg_12028 <= cipher_0_ssbox_q140;
        tmp_V_24_reg_12058 <= cipher_0_ssbox_q135;
        tmp_V_25_reg_12088 <= cipher_0_ssbox_q130;
        tmp_V_27_reg_12052 <= cipher_0_ssbox_q136;
        tmp_V_28_reg_12082 <= cipher_0_ssbox_q131;
        tmp_V_31_reg_12076 <= cipher_0_ssbox_q132;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        tmp_1_V_12_reg_12272 <= cipher_0_ssbox_q126;
        tmp_2_1_V_12_reg_12278 <= cipher_0_ssbox_q125;
        tmp_2_2_V_12_reg_12302 <= cipher_0_ssbox_q121;
        tmp_3_V_12_reg_12356 <= cipher_0_ssbox_q112;
        tmp_V_32_reg_12266 <= cipher_0_ssbox_q127;
        tmp_V_33_reg_12296 <= cipher_0_ssbox_q122;
        tmp_V_34_reg_12326 <= cipher_0_ssbox_q117;
        tmp_V_36_reg_12290 <= cipher_0_ssbox_q123;
        tmp_V_37_reg_12320 <= cipher_0_ssbox_q118;
        tmp_V_38_reg_12350 <= cipher_0_ssbox_q113;
        tmp_V_39_reg_12284 <= cipher_0_ssbox_q124;
        tmp_V_40_reg_12314 <= cipher_0_ssbox_q119;
        tmp_V_41_reg_12344 <= cipher_0_ssbox_q114;
        tmp_V_43_reg_12308 <= cipher_0_ssbox_q120;
        tmp_V_44_reg_12338 <= cipher_0_ssbox_q115;
        tmp_V_47_reg_12332 <= cipher_0_ssbox_q116;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        tmp_1_V_13_reg_12528 <= cipher_0_ssbox_q110;
        tmp_2_1_V_13_reg_12534 <= cipher_0_ssbox_q109;
        tmp_2_2_V_13_reg_12558 <= cipher_0_ssbox_q105;
        tmp_3_V_13_reg_12612 <= cipher_0_ssbox_q96;
        tmp_V_48_reg_12522 <= cipher_0_ssbox_q111;
        tmp_V_49_reg_12552 <= cipher_0_ssbox_q106;
        tmp_V_50_reg_12582 <= cipher_0_ssbox_q101;
        tmp_V_52_reg_12546 <= cipher_0_ssbox_q107;
        tmp_V_53_reg_12576 <= cipher_0_ssbox_q102;
        tmp_V_54_reg_12606 <= cipher_0_ssbox_q97;
        tmp_V_55_reg_12540 <= cipher_0_ssbox_q108;
        tmp_V_56_reg_12570 <= cipher_0_ssbox_q103;
        tmp_V_57_reg_12600 <= cipher_0_ssbox_q98;
        tmp_V_59_reg_12564 <= cipher_0_ssbox_q104;
        tmp_V_60_reg_12594 <= cipher_0_ssbox_q99;
        tmp_V_63_reg_12588 <= cipher_0_ssbox_q100;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        tmp_1_V_14_reg_12784 <= cipher_0_ssbox_q94;
        tmp_2_1_V_14_reg_12790 <= cipher_0_ssbox_q93;
        tmp_2_2_V_14_reg_12814 <= cipher_0_ssbox_q89;
        tmp_3_V_14_reg_12868 <= cipher_0_ssbox_q80;
        tmp_V_64_reg_12778 <= cipher_0_ssbox_q95;
        tmp_V_65_reg_12808 <= cipher_0_ssbox_q90;
        tmp_V_66_reg_12838 <= cipher_0_ssbox_q85;
        tmp_V_68_reg_12802 <= cipher_0_ssbox_q91;
        tmp_V_69_reg_12832 <= cipher_0_ssbox_q86;
        tmp_V_70_reg_12862 <= cipher_0_ssbox_q81;
        tmp_V_71_reg_12796 <= cipher_0_ssbox_q92;
        tmp_V_72_reg_12826 <= cipher_0_ssbox_q87;
        tmp_V_73_reg_12856 <= cipher_0_ssbox_q82;
        tmp_V_75_reg_12820 <= cipher_0_ssbox_q88;
        tmp_V_76_reg_12850 <= cipher_0_ssbox_q83;
        tmp_V_79_reg_12844 <= cipher_0_ssbox_q84;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        tmp_1_V_15_reg_13040 <= cipher_0_ssbox_q78;
        tmp_2_1_V_15_reg_13046 <= cipher_0_ssbox_q77;
        tmp_2_2_V_15_reg_13070 <= cipher_0_ssbox_q73;
        tmp_3_V_15_reg_13124 <= cipher_0_ssbox_q64;
        tmp_V_80_reg_13034 <= cipher_0_ssbox_q79;
        tmp_V_81_reg_13064 <= cipher_0_ssbox_q74;
        tmp_V_82_reg_13094 <= cipher_0_ssbox_q69;
        tmp_V_84_reg_13058 <= cipher_0_ssbox_q75;
        tmp_V_85_reg_13088 <= cipher_0_ssbox_q70;
        tmp_V_86_reg_13118 <= cipher_0_ssbox_q65;
        tmp_V_87_reg_13052 <= cipher_0_ssbox_q76;
        tmp_V_88_reg_13082 <= cipher_0_ssbox_q71;
        tmp_V_89_reg_13112 <= cipher_0_ssbox_q66;
        tmp_V_91_reg_13076 <= cipher_0_ssbox_q72;
        tmp_V_92_reg_13106 <= cipher_0_ssbox_q67;
        tmp_V_95_reg_13100 <= cipher_0_ssbox_q68;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        tmp_1_V_16_reg_13296 <= cipher_0_ssbox_q62;
        tmp_2_1_V_16_reg_13302 <= cipher_0_ssbox_q61;
        tmp_2_2_V_16_reg_13326 <= cipher_0_ssbox_q57;
        tmp_3_V_16_reg_13380 <= cipher_0_ssbox_q48;
        tmp_V_100_reg_13314 <= cipher_0_ssbox_q59;
        tmp_V_101_reg_13344 <= cipher_0_ssbox_q54;
        tmp_V_102_reg_13374 <= cipher_0_ssbox_q49;
        tmp_V_103_reg_13308 <= cipher_0_ssbox_q60;
        tmp_V_104_reg_13338 <= cipher_0_ssbox_q55;
        tmp_V_105_reg_13368 <= cipher_0_ssbox_q50;
        tmp_V_107_reg_13332 <= cipher_0_ssbox_q56;
        tmp_V_108_reg_13362 <= cipher_0_ssbox_q51;
        tmp_V_111_reg_13356 <= cipher_0_ssbox_q52;
        tmp_V_96_reg_13290 <= cipher_0_ssbox_q63;
        tmp_V_97_reg_13320 <= cipher_0_ssbox_q58;
        tmp_V_98_reg_13350 <= cipher_0_ssbox_q53;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        tmp_1_V_17_reg_13552 <= cipher_0_ssbox_q46;
        tmp_2_1_V_17_reg_13558 <= cipher_0_ssbox_q45;
        tmp_2_2_V_17_reg_13582 <= cipher_0_ssbox_q41;
        tmp_3_V_17_reg_13636 <= cipher_0_ssbox_q32;
        tmp_V_112_reg_13546 <= cipher_0_ssbox_q47;
        tmp_V_113_reg_13576 <= cipher_0_ssbox_q42;
        tmp_V_114_reg_13606 <= cipher_0_ssbox_q37;
        tmp_V_116_reg_13570 <= cipher_0_ssbox_q43;
        tmp_V_117_reg_13600 <= cipher_0_ssbox_q38;
        tmp_V_118_reg_13630 <= cipher_0_ssbox_q33;
        tmp_V_119_reg_13564 <= cipher_0_ssbox_q44;
        tmp_V_120_reg_13594 <= cipher_0_ssbox_q39;
        tmp_V_121_reg_13624 <= cipher_0_ssbox_q34;
        tmp_V_123_reg_13588 <= cipher_0_ssbox_q40;
        tmp_V_124_reg_13618 <= cipher_0_ssbox_q35;
        tmp_V_127_reg_13612 <= cipher_0_ssbox_q36;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        tmp_1_V_18_reg_13808 <= cipher_0_ssbox_q30;
        tmp_2_1_V_18_reg_13814 <= cipher_0_ssbox_q29;
        tmp_2_2_V_18_reg_13838 <= cipher_0_ssbox_q25;
        tmp_3_V_18_reg_13892 <= cipher_0_ssbox_q16;
        tmp_V_128_reg_13802 <= cipher_0_ssbox_q31;
        tmp_V_129_reg_13832 <= cipher_0_ssbox_q26;
        tmp_V_130_reg_13862 <= cipher_0_ssbox_q21;
        tmp_V_132_reg_13826 <= cipher_0_ssbox_q27;
        tmp_V_133_reg_13856 <= cipher_0_ssbox_q22;
        tmp_V_134_reg_13886 <= cipher_0_ssbox_q17;
        tmp_V_135_reg_13820 <= cipher_0_ssbox_q28;
        tmp_V_136_reg_13850 <= cipher_0_ssbox_q23;
        tmp_V_137_reg_13880 <= cipher_0_ssbox_q18;
        tmp_V_139_reg_13844 <= cipher_0_ssbox_q24;
        tmp_V_140_reg_13874 <= cipher_0_ssbox_q19;
        tmp_V_143_reg_13868 <= cipher_0_ssbox_q20;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_idle_pp0 == 1'b1) & (ap_start == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b0) & (ap_enable_reg_pp0_iter18 == 1'b0) & (ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b0) & (ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0_0to18 = 1'b1;
    end else begin
        ap_idle_pp0_0to18 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((ap_idle_pp0_0to18 == 1'b1) & (ap_start == 1'b0))) begin
        ap_reset_idle_pp0 = 1'b1;
    end else begin
        ap_reset_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce0 = 1'b1;
    end else begin
        cipher_0_p16box_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce1 = 1'b1;
    end else begin
        cipher_0_p16box_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce10 = 1'b1;
    end else begin
        cipher_0_p16box_ce10 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce100 = 1'b1;
    end else begin
        cipher_0_p16box_ce100 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce101 = 1'b1;
    end else begin
        cipher_0_p16box_ce101 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce102 = 1'b1;
    end else begin
        cipher_0_p16box_ce102 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce103 = 1'b1;
    end else begin
        cipher_0_p16box_ce103 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce104 = 1'b1;
    end else begin
        cipher_0_p16box_ce104 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce105 = 1'b1;
    end else begin
        cipher_0_p16box_ce105 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce106 = 1'b1;
    end else begin
        cipher_0_p16box_ce106 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce107 = 1'b1;
    end else begin
        cipher_0_p16box_ce107 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce108 = 1'b1;
    end else begin
        cipher_0_p16box_ce108 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce109 = 1'b1;
    end else begin
        cipher_0_p16box_ce109 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce11 = 1'b1;
    end else begin
        cipher_0_p16box_ce11 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce110 = 1'b1;
    end else begin
        cipher_0_p16box_ce110 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce111 = 1'b1;
    end else begin
        cipher_0_p16box_ce111 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce112 = 1'b1;
    end else begin
        cipher_0_p16box_ce112 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce113 = 1'b1;
    end else begin
        cipher_0_p16box_ce113 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce114 = 1'b1;
    end else begin
        cipher_0_p16box_ce114 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce115 = 1'b1;
    end else begin
        cipher_0_p16box_ce115 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce116 = 1'b1;
    end else begin
        cipher_0_p16box_ce116 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce117 = 1'b1;
    end else begin
        cipher_0_p16box_ce117 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce118 = 1'b1;
    end else begin
        cipher_0_p16box_ce118 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce119 = 1'b1;
    end else begin
        cipher_0_p16box_ce119 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce12 = 1'b1;
    end else begin
        cipher_0_p16box_ce12 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce120 = 1'b1;
    end else begin
        cipher_0_p16box_ce120 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce121 = 1'b1;
    end else begin
        cipher_0_p16box_ce121 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce122 = 1'b1;
    end else begin
        cipher_0_p16box_ce122 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce123 = 1'b1;
    end else begin
        cipher_0_p16box_ce123 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce124 = 1'b1;
    end else begin
        cipher_0_p16box_ce124 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce125 = 1'b1;
    end else begin
        cipher_0_p16box_ce125 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce126 = 1'b1;
    end else begin
        cipher_0_p16box_ce126 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce127 = 1'b1;
    end else begin
        cipher_0_p16box_ce127 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce128 = 1'b1;
    end else begin
        cipher_0_p16box_ce128 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce129 = 1'b1;
    end else begin
        cipher_0_p16box_ce129 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce13 = 1'b1;
    end else begin
        cipher_0_p16box_ce13 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce130 = 1'b1;
    end else begin
        cipher_0_p16box_ce130 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce131 = 1'b1;
    end else begin
        cipher_0_p16box_ce131 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce132 = 1'b1;
    end else begin
        cipher_0_p16box_ce132 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce133 = 1'b1;
    end else begin
        cipher_0_p16box_ce133 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce134 = 1'b1;
    end else begin
        cipher_0_p16box_ce134 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce135 = 1'b1;
    end else begin
        cipher_0_p16box_ce135 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce136 = 1'b1;
    end else begin
        cipher_0_p16box_ce136 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce137 = 1'b1;
    end else begin
        cipher_0_p16box_ce137 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce138 = 1'b1;
    end else begin
        cipher_0_p16box_ce138 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce139 = 1'b1;
    end else begin
        cipher_0_p16box_ce139 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce14 = 1'b1;
    end else begin
        cipher_0_p16box_ce14 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce140 = 1'b1;
    end else begin
        cipher_0_p16box_ce140 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce141 = 1'b1;
    end else begin
        cipher_0_p16box_ce141 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce142 = 1'b1;
    end else begin
        cipher_0_p16box_ce142 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce143 = 1'b1;
    end else begin
        cipher_0_p16box_ce143 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce15 = 1'b1;
    end else begin
        cipher_0_p16box_ce15 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce16 = 1'b1;
    end else begin
        cipher_0_p16box_ce16 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce17 = 1'b1;
    end else begin
        cipher_0_p16box_ce17 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce18 = 1'b1;
    end else begin
        cipher_0_p16box_ce18 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce19 = 1'b1;
    end else begin
        cipher_0_p16box_ce19 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce2 = 1'b1;
    end else begin
        cipher_0_p16box_ce2 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce20 = 1'b1;
    end else begin
        cipher_0_p16box_ce20 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce21 = 1'b1;
    end else begin
        cipher_0_p16box_ce21 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce22 = 1'b1;
    end else begin
        cipher_0_p16box_ce22 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce23 = 1'b1;
    end else begin
        cipher_0_p16box_ce23 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce24 = 1'b1;
    end else begin
        cipher_0_p16box_ce24 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce25 = 1'b1;
    end else begin
        cipher_0_p16box_ce25 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce26 = 1'b1;
    end else begin
        cipher_0_p16box_ce26 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce27 = 1'b1;
    end else begin
        cipher_0_p16box_ce27 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce28 = 1'b1;
    end else begin
        cipher_0_p16box_ce28 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce29 = 1'b1;
    end else begin
        cipher_0_p16box_ce29 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce3 = 1'b1;
    end else begin
        cipher_0_p16box_ce3 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce30 = 1'b1;
    end else begin
        cipher_0_p16box_ce30 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce31 = 1'b1;
    end else begin
        cipher_0_p16box_ce31 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce32 = 1'b1;
    end else begin
        cipher_0_p16box_ce32 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce33 = 1'b1;
    end else begin
        cipher_0_p16box_ce33 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce34 = 1'b1;
    end else begin
        cipher_0_p16box_ce34 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce35 = 1'b1;
    end else begin
        cipher_0_p16box_ce35 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce36 = 1'b1;
    end else begin
        cipher_0_p16box_ce36 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce37 = 1'b1;
    end else begin
        cipher_0_p16box_ce37 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce38 = 1'b1;
    end else begin
        cipher_0_p16box_ce38 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce39 = 1'b1;
    end else begin
        cipher_0_p16box_ce39 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce4 = 1'b1;
    end else begin
        cipher_0_p16box_ce4 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce40 = 1'b1;
    end else begin
        cipher_0_p16box_ce40 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce41 = 1'b1;
    end else begin
        cipher_0_p16box_ce41 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce42 = 1'b1;
    end else begin
        cipher_0_p16box_ce42 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce43 = 1'b1;
    end else begin
        cipher_0_p16box_ce43 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce44 = 1'b1;
    end else begin
        cipher_0_p16box_ce44 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce45 = 1'b1;
    end else begin
        cipher_0_p16box_ce45 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce46 = 1'b1;
    end else begin
        cipher_0_p16box_ce46 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce47 = 1'b1;
    end else begin
        cipher_0_p16box_ce47 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce48 = 1'b1;
    end else begin
        cipher_0_p16box_ce48 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce49 = 1'b1;
    end else begin
        cipher_0_p16box_ce49 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce5 = 1'b1;
    end else begin
        cipher_0_p16box_ce5 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce50 = 1'b1;
    end else begin
        cipher_0_p16box_ce50 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce51 = 1'b1;
    end else begin
        cipher_0_p16box_ce51 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce52 = 1'b1;
    end else begin
        cipher_0_p16box_ce52 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce53 = 1'b1;
    end else begin
        cipher_0_p16box_ce53 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce54 = 1'b1;
    end else begin
        cipher_0_p16box_ce54 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce55 = 1'b1;
    end else begin
        cipher_0_p16box_ce55 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce56 = 1'b1;
    end else begin
        cipher_0_p16box_ce56 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce57 = 1'b1;
    end else begin
        cipher_0_p16box_ce57 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce58 = 1'b1;
    end else begin
        cipher_0_p16box_ce58 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce59 = 1'b1;
    end else begin
        cipher_0_p16box_ce59 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce6 = 1'b1;
    end else begin
        cipher_0_p16box_ce6 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce60 = 1'b1;
    end else begin
        cipher_0_p16box_ce60 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce61 = 1'b1;
    end else begin
        cipher_0_p16box_ce61 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce62 = 1'b1;
    end else begin
        cipher_0_p16box_ce62 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce63 = 1'b1;
    end else begin
        cipher_0_p16box_ce63 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce64 = 1'b1;
    end else begin
        cipher_0_p16box_ce64 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce65 = 1'b1;
    end else begin
        cipher_0_p16box_ce65 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce66 = 1'b1;
    end else begin
        cipher_0_p16box_ce66 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce67 = 1'b1;
    end else begin
        cipher_0_p16box_ce67 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce68 = 1'b1;
    end else begin
        cipher_0_p16box_ce68 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce69 = 1'b1;
    end else begin
        cipher_0_p16box_ce69 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce7 = 1'b1;
    end else begin
        cipher_0_p16box_ce7 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce70 = 1'b1;
    end else begin
        cipher_0_p16box_ce70 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce71 = 1'b1;
    end else begin
        cipher_0_p16box_ce71 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce72 = 1'b1;
    end else begin
        cipher_0_p16box_ce72 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce73 = 1'b1;
    end else begin
        cipher_0_p16box_ce73 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce74 = 1'b1;
    end else begin
        cipher_0_p16box_ce74 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce75 = 1'b1;
    end else begin
        cipher_0_p16box_ce75 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce76 = 1'b1;
    end else begin
        cipher_0_p16box_ce76 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce77 = 1'b1;
    end else begin
        cipher_0_p16box_ce77 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce78 = 1'b1;
    end else begin
        cipher_0_p16box_ce78 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce79 = 1'b1;
    end else begin
        cipher_0_p16box_ce79 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce8 = 1'b1;
    end else begin
        cipher_0_p16box_ce8 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce80 = 1'b1;
    end else begin
        cipher_0_p16box_ce80 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce81 = 1'b1;
    end else begin
        cipher_0_p16box_ce81 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce82 = 1'b1;
    end else begin
        cipher_0_p16box_ce82 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce83 = 1'b1;
    end else begin
        cipher_0_p16box_ce83 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce84 = 1'b1;
    end else begin
        cipher_0_p16box_ce84 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce85 = 1'b1;
    end else begin
        cipher_0_p16box_ce85 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce86 = 1'b1;
    end else begin
        cipher_0_p16box_ce86 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce87 = 1'b1;
    end else begin
        cipher_0_p16box_ce87 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce88 = 1'b1;
    end else begin
        cipher_0_p16box_ce88 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce89 = 1'b1;
    end else begin
        cipher_0_p16box_ce89 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce9 = 1'b1;
    end else begin
        cipher_0_p16box_ce9 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce90 = 1'b1;
    end else begin
        cipher_0_p16box_ce90 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce91 = 1'b1;
    end else begin
        cipher_0_p16box_ce91 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce92 = 1'b1;
    end else begin
        cipher_0_p16box_ce92 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce93 = 1'b1;
    end else begin
        cipher_0_p16box_ce93 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce94 = 1'b1;
    end else begin
        cipher_0_p16box_ce94 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce95 = 1'b1;
    end else begin
        cipher_0_p16box_ce95 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce96 = 1'b1;
    end else begin
        cipher_0_p16box_ce96 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce97 = 1'b1;
    end else begin
        cipher_0_p16box_ce97 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce98 = 1'b1;
    end else begin
        cipher_0_p16box_ce98 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_p16box_ce99 = 1'b1;
    end else begin
        cipher_0_p16box_ce99 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce0 = 1'b1;
    end else begin
        cipher_0_ssbox_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce1 = 1'b1;
    end else begin
        cipher_0_ssbox_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce10 = 1'b1;
    end else begin
        cipher_0_ssbox_ce10 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce100 = 1'b1;
    end else begin
        cipher_0_ssbox_ce100 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce101 = 1'b1;
    end else begin
        cipher_0_ssbox_ce101 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce102 = 1'b1;
    end else begin
        cipher_0_ssbox_ce102 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce103 = 1'b1;
    end else begin
        cipher_0_ssbox_ce103 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce104 = 1'b1;
    end else begin
        cipher_0_ssbox_ce104 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce105 = 1'b1;
    end else begin
        cipher_0_ssbox_ce105 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce106 = 1'b1;
    end else begin
        cipher_0_ssbox_ce106 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce107 = 1'b1;
    end else begin
        cipher_0_ssbox_ce107 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce108 = 1'b1;
    end else begin
        cipher_0_ssbox_ce108 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce109 = 1'b1;
    end else begin
        cipher_0_ssbox_ce109 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce11 = 1'b1;
    end else begin
        cipher_0_ssbox_ce11 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce110 = 1'b1;
    end else begin
        cipher_0_ssbox_ce110 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce111 = 1'b1;
    end else begin
        cipher_0_ssbox_ce111 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce112 = 1'b1;
    end else begin
        cipher_0_ssbox_ce112 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce113 = 1'b1;
    end else begin
        cipher_0_ssbox_ce113 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce114 = 1'b1;
    end else begin
        cipher_0_ssbox_ce114 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce115 = 1'b1;
    end else begin
        cipher_0_ssbox_ce115 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce116 = 1'b1;
    end else begin
        cipher_0_ssbox_ce116 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce117 = 1'b1;
    end else begin
        cipher_0_ssbox_ce117 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce118 = 1'b1;
    end else begin
        cipher_0_ssbox_ce118 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce119 = 1'b1;
    end else begin
        cipher_0_ssbox_ce119 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce12 = 1'b1;
    end else begin
        cipher_0_ssbox_ce12 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce120 = 1'b1;
    end else begin
        cipher_0_ssbox_ce120 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce121 = 1'b1;
    end else begin
        cipher_0_ssbox_ce121 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce122 = 1'b1;
    end else begin
        cipher_0_ssbox_ce122 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce123 = 1'b1;
    end else begin
        cipher_0_ssbox_ce123 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce124 = 1'b1;
    end else begin
        cipher_0_ssbox_ce124 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce125 = 1'b1;
    end else begin
        cipher_0_ssbox_ce125 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce126 = 1'b1;
    end else begin
        cipher_0_ssbox_ce126 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce127 = 1'b1;
    end else begin
        cipher_0_ssbox_ce127 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce128 = 1'b1;
    end else begin
        cipher_0_ssbox_ce128 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce129 = 1'b1;
    end else begin
        cipher_0_ssbox_ce129 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce13 = 1'b1;
    end else begin
        cipher_0_ssbox_ce13 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce130 = 1'b1;
    end else begin
        cipher_0_ssbox_ce130 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce131 = 1'b1;
    end else begin
        cipher_0_ssbox_ce131 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce132 = 1'b1;
    end else begin
        cipher_0_ssbox_ce132 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce133 = 1'b1;
    end else begin
        cipher_0_ssbox_ce133 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce134 = 1'b1;
    end else begin
        cipher_0_ssbox_ce134 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce135 = 1'b1;
    end else begin
        cipher_0_ssbox_ce135 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce136 = 1'b1;
    end else begin
        cipher_0_ssbox_ce136 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce137 = 1'b1;
    end else begin
        cipher_0_ssbox_ce137 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce138 = 1'b1;
    end else begin
        cipher_0_ssbox_ce138 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce139 = 1'b1;
    end else begin
        cipher_0_ssbox_ce139 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce14 = 1'b1;
    end else begin
        cipher_0_ssbox_ce14 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce140 = 1'b1;
    end else begin
        cipher_0_ssbox_ce140 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce141 = 1'b1;
    end else begin
        cipher_0_ssbox_ce141 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce142 = 1'b1;
    end else begin
        cipher_0_ssbox_ce142 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce143 = 1'b1;
    end else begin
        cipher_0_ssbox_ce143 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce144 = 1'b1;
    end else begin
        cipher_0_ssbox_ce144 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce145 = 1'b1;
    end else begin
        cipher_0_ssbox_ce145 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce146 = 1'b1;
    end else begin
        cipher_0_ssbox_ce146 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce147 = 1'b1;
    end else begin
        cipher_0_ssbox_ce147 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce148 = 1'b1;
    end else begin
        cipher_0_ssbox_ce148 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce149 = 1'b1;
    end else begin
        cipher_0_ssbox_ce149 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce15 = 1'b1;
    end else begin
        cipher_0_ssbox_ce15 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce150 = 1'b1;
    end else begin
        cipher_0_ssbox_ce150 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce151 = 1'b1;
    end else begin
        cipher_0_ssbox_ce151 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce152 = 1'b1;
    end else begin
        cipher_0_ssbox_ce152 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce153 = 1'b1;
    end else begin
        cipher_0_ssbox_ce153 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce154 = 1'b1;
    end else begin
        cipher_0_ssbox_ce154 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce155 = 1'b1;
    end else begin
        cipher_0_ssbox_ce155 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce156 = 1'b1;
    end else begin
        cipher_0_ssbox_ce156 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce157 = 1'b1;
    end else begin
        cipher_0_ssbox_ce157 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce158 = 1'b1;
    end else begin
        cipher_0_ssbox_ce158 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce159 = 1'b1;
    end else begin
        cipher_0_ssbox_ce159 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce16 = 1'b1;
    end else begin
        cipher_0_ssbox_ce16 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce17 = 1'b1;
    end else begin
        cipher_0_ssbox_ce17 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce18 = 1'b1;
    end else begin
        cipher_0_ssbox_ce18 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce19 = 1'b1;
    end else begin
        cipher_0_ssbox_ce19 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce2 = 1'b1;
    end else begin
        cipher_0_ssbox_ce2 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce20 = 1'b1;
    end else begin
        cipher_0_ssbox_ce20 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce21 = 1'b1;
    end else begin
        cipher_0_ssbox_ce21 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce22 = 1'b1;
    end else begin
        cipher_0_ssbox_ce22 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce23 = 1'b1;
    end else begin
        cipher_0_ssbox_ce23 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce24 = 1'b1;
    end else begin
        cipher_0_ssbox_ce24 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce25 = 1'b1;
    end else begin
        cipher_0_ssbox_ce25 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce26 = 1'b1;
    end else begin
        cipher_0_ssbox_ce26 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce27 = 1'b1;
    end else begin
        cipher_0_ssbox_ce27 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce28 = 1'b1;
    end else begin
        cipher_0_ssbox_ce28 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce29 = 1'b1;
    end else begin
        cipher_0_ssbox_ce29 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce3 = 1'b1;
    end else begin
        cipher_0_ssbox_ce3 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce30 = 1'b1;
    end else begin
        cipher_0_ssbox_ce30 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce31 = 1'b1;
    end else begin
        cipher_0_ssbox_ce31 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce32 = 1'b1;
    end else begin
        cipher_0_ssbox_ce32 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce33 = 1'b1;
    end else begin
        cipher_0_ssbox_ce33 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce34 = 1'b1;
    end else begin
        cipher_0_ssbox_ce34 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce35 = 1'b1;
    end else begin
        cipher_0_ssbox_ce35 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce36 = 1'b1;
    end else begin
        cipher_0_ssbox_ce36 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce37 = 1'b1;
    end else begin
        cipher_0_ssbox_ce37 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce38 = 1'b1;
    end else begin
        cipher_0_ssbox_ce38 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce39 = 1'b1;
    end else begin
        cipher_0_ssbox_ce39 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce4 = 1'b1;
    end else begin
        cipher_0_ssbox_ce4 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce40 = 1'b1;
    end else begin
        cipher_0_ssbox_ce40 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce41 = 1'b1;
    end else begin
        cipher_0_ssbox_ce41 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce42 = 1'b1;
    end else begin
        cipher_0_ssbox_ce42 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce43 = 1'b1;
    end else begin
        cipher_0_ssbox_ce43 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce44 = 1'b1;
    end else begin
        cipher_0_ssbox_ce44 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce45 = 1'b1;
    end else begin
        cipher_0_ssbox_ce45 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce46 = 1'b1;
    end else begin
        cipher_0_ssbox_ce46 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce47 = 1'b1;
    end else begin
        cipher_0_ssbox_ce47 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce48 = 1'b1;
    end else begin
        cipher_0_ssbox_ce48 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce49 = 1'b1;
    end else begin
        cipher_0_ssbox_ce49 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce5 = 1'b1;
    end else begin
        cipher_0_ssbox_ce5 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce50 = 1'b1;
    end else begin
        cipher_0_ssbox_ce50 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce51 = 1'b1;
    end else begin
        cipher_0_ssbox_ce51 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce52 = 1'b1;
    end else begin
        cipher_0_ssbox_ce52 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce53 = 1'b1;
    end else begin
        cipher_0_ssbox_ce53 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce54 = 1'b1;
    end else begin
        cipher_0_ssbox_ce54 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce55 = 1'b1;
    end else begin
        cipher_0_ssbox_ce55 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce56 = 1'b1;
    end else begin
        cipher_0_ssbox_ce56 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce57 = 1'b1;
    end else begin
        cipher_0_ssbox_ce57 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce58 = 1'b1;
    end else begin
        cipher_0_ssbox_ce58 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce59 = 1'b1;
    end else begin
        cipher_0_ssbox_ce59 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce6 = 1'b1;
    end else begin
        cipher_0_ssbox_ce6 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce60 = 1'b1;
    end else begin
        cipher_0_ssbox_ce60 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce61 = 1'b1;
    end else begin
        cipher_0_ssbox_ce61 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce62 = 1'b1;
    end else begin
        cipher_0_ssbox_ce62 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce63 = 1'b1;
    end else begin
        cipher_0_ssbox_ce63 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce64 = 1'b1;
    end else begin
        cipher_0_ssbox_ce64 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce65 = 1'b1;
    end else begin
        cipher_0_ssbox_ce65 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce66 = 1'b1;
    end else begin
        cipher_0_ssbox_ce66 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce67 = 1'b1;
    end else begin
        cipher_0_ssbox_ce67 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce68 = 1'b1;
    end else begin
        cipher_0_ssbox_ce68 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce69 = 1'b1;
    end else begin
        cipher_0_ssbox_ce69 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce7 = 1'b1;
    end else begin
        cipher_0_ssbox_ce7 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce70 = 1'b1;
    end else begin
        cipher_0_ssbox_ce70 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce71 = 1'b1;
    end else begin
        cipher_0_ssbox_ce71 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce72 = 1'b1;
    end else begin
        cipher_0_ssbox_ce72 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce73 = 1'b1;
    end else begin
        cipher_0_ssbox_ce73 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce74 = 1'b1;
    end else begin
        cipher_0_ssbox_ce74 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce75 = 1'b1;
    end else begin
        cipher_0_ssbox_ce75 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce76 = 1'b1;
    end else begin
        cipher_0_ssbox_ce76 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce77 = 1'b1;
    end else begin
        cipher_0_ssbox_ce77 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce78 = 1'b1;
    end else begin
        cipher_0_ssbox_ce78 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce79 = 1'b1;
    end else begin
        cipher_0_ssbox_ce79 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce8 = 1'b1;
    end else begin
        cipher_0_ssbox_ce8 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce80 = 1'b1;
    end else begin
        cipher_0_ssbox_ce80 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce81 = 1'b1;
    end else begin
        cipher_0_ssbox_ce81 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce82 = 1'b1;
    end else begin
        cipher_0_ssbox_ce82 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce83 = 1'b1;
    end else begin
        cipher_0_ssbox_ce83 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce84 = 1'b1;
    end else begin
        cipher_0_ssbox_ce84 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce85 = 1'b1;
    end else begin
        cipher_0_ssbox_ce85 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce86 = 1'b1;
    end else begin
        cipher_0_ssbox_ce86 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce87 = 1'b1;
    end else begin
        cipher_0_ssbox_ce87 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce88 = 1'b1;
    end else begin
        cipher_0_ssbox_ce88 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce89 = 1'b1;
    end else begin
        cipher_0_ssbox_ce89 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce9 = 1'b1;
    end else begin
        cipher_0_ssbox_ce9 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce90 = 1'b1;
    end else begin
        cipher_0_ssbox_ce90 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce91 = 1'b1;
    end else begin
        cipher_0_ssbox_ce91 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce92 = 1'b1;
    end else begin
        cipher_0_ssbox_ce92 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce93 = 1'b1;
    end else begin
        cipher_0_ssbox_ce93 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce94 = 1'b1;
    end else begin
        cipher_0_ssbox_ce94 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce95 = 1'b1;
    end else begin
        cipher_0_ssbox_ce95 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce96 = 1'b1;
    end else begin
        cipher_0_ssbox_ce96 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce97 = 1'b1;
    end else begin
        cipher_0_ssbox_ce97 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce98 = 1'b1;
    end else begin
        cipher_0_ssbox_ce98 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        cipher_0_ssbox_ce99 = 1'b1;
    end else begin
        cipher_0_ssbox_ce99 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_state10_pp0_stage0_iter9 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage0_iter10 = ~(1'b1 == 1'b1);

assign ap_block_state12_pp0_stage0_iter11 = ~(1'b1 == 1'b1);

assign ap_block_state13_pp0_stage0_iter12 = ~(1'b1 == 1'b1);

assign ap_block_state14_pp0_stage0_iter13 = ~(1'b1 == 1'b1);

assign ap_block_state15_pp0_stage0_iter14 = ~(1'b1 == 1'b1);

assign ap_block_state16_pp0_stage0_iter15 = ~(1'b1 == 1'b1);

assign ap_block_state17_pp0_stage0_iter16 = ~(1'b1 == 1'b1);

assign ap_block_state18_pp0_stage0_iter17 = ~(1'b1 == 1'b1);

assign ap_block_state19_pp0_stage0_iter18 = ~(1'b1 == 1'b1);

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state20_pp0_stage0_iter19 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter8 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_enable_reg_pp0_iter0 = ap_start;

assign ap_return = (p_read_1_reg_11624_pp0_iter18_reg ^ p_Result_10_fu_11583_p17);

assign cipher_0_p16box_address0 = zext_ln587_143_fu_10823_p1;

assign cipher_0_p16box_address1 = zext_ln587_142_fu_10818_p1;

assign cipher_0_p16box_address10 = zext_ln587_133_fu_10773_p1;

assign cipher_0_p16box_address100 = zext_ln587_43_fu_5793_p1;

assign cipher_0_p16box_address101 = zext_ln587_42_fu_5788_p1;

assign cipher_0_p16box_address102 = zext_ln587_41_fu_5783_p1;

assign cipher_0_p16box_address103 = zext_ln587_40_fu_5778_p1;

assign cipher_0_p16box_address104 = zext_ln587_39_fu_5773_p1;

assign cipher_0_p16box_address105 = zext_ln587_38_fu_5768_p1;

assign cipher_0_p16box_address106 = zext_ln587_37_fu_5763_p1;

assign cipher_0_p16box_address107 = zext_ln587_36_fu_5758_p1;

assign cipher_0_p16box_address108 = zext_ln587_35_fu_5753_p1;

assign cipher_0_p16box_address109 = zext_ln587_34_fu_5748_p1;

assign cipher_0_p16box_address11 = zext_ln587_132_fu_10768_p1;

assign cipher_0_p16box_address110 = zext_ln587_33_fu_5743_p1;

assign cipher_0_p16box_address111 = zext_ln587_32_fu_5738_p1;

assign cipher_0_p16box_address112 = zext_ln587_31_fu_4978_p1;

assign cipher_0_p16box_address113 = zext_ln587_30_fu_4973_p1;

assign cipher_0_p16box_address114 = zext_ln587_29_fu_4968_p1;

assign cipher_0_p16box_address115 = zext_ln587_28_fu_4963_p1;

assign cipher_0_p16box_address116 = zext_ln587_27_fu_4958_p1;

assign cipher_0_p16box_address117 = zext_ln587_26_fu_4953_p1;

assign cipher_0_p16box_address118 = zext_ln587_25_fu_4948_p1;

assign cipher_0_p16box_address119 = zext_ln587_24_fu_4943_p1;

assign cipher_0_p16box_address12 = zext_ln587_131_fu_10763_p1;

assign cipher_0_p16box_address120 = zext_ln587_23_fu_4938_p1;

assign cipher_0_p16box_address121 = zext_ln587_22_fu_4933_p1;

assign cipher_0_p16box_address122 = zext_ln587_21_fu_4928_p1;

assign cipher_0_p16box_address123 = zext_ln587_20_fu_4923_p1;

assign cipher_0_p16box_address124 = zext_ln587_19_fu_4918_p1;

assign cipher_0_p16box_address125 = zext_ln587_18_fu_4913_p1;

assign cipher_0_p16box_address126 = zext_ln587_17_fu_4908_p1;

assign cipher_0_p16box_address127 = zext_ln587_16_fu_4903_p1;

assign cipher_0_p16box_address128 = zext_ln587_15_fu_4143_p1;

assign cipher_0_p16box_address129 = zext_ln587_14_fu_4138_p1;

assign cipher_0_p16box_address13 = zext_ln587_130_fu_10758_p1;

assign cipher_0_p16box_address130 = zext_ln587_13_fu_4133_p1;

assign cipher_0_p16box_address131 = zext_ln587_12_fu_4128_p1;

assign cipher_0_p16box_address132 = zext_ln587_11_fu_4123_p1;

assign cipher_0_p16box_address133 = zext_ln587_10_fu_4118_p1;

assign cipher_0_p16box_address134 = zext_ln587_9_fu_4113_p1;

assign cipher_0_p16box_address135 = zext_ln587_8_fu_4108_p1;

assign cipher_0_p16box_address136 = zext_ln587_7_fu_4103_p1;

assign cipher_0_p16box_address137 = zext_ln587_6_fu_4098_p1;

assign cipher_0_p16box_address138 = zext_ln587_5_fu_4093_p1;

assign cipher_0_p16box_address139 = zext_ln587_4_fu_4088_p1;

assign cipher_0_p16box_address14 = zext_ln587_129_fu_10753_p1;

assign cipher_0_p16box_address140 = zext_ln587_3_fu_4083_p1;

assign cipher_0_p16box_address141 = zext_ln587_2_fu_4078_p1;

assign cipher_0_p16box_address142 = zext_ln587_1_fu_4073_p1;

assign cipher_0_p16box_address143 = zext_ln587_fu_4068_p1;

assign cipher_0_p16box_address15 = zext_ln587_128_fu_10748_p1;

assign cipher_0_p16box_address16 = zext_ln587_127_fu_9988_p1;

assign cipher_0_p16box_address17 = zext_ln587_126_fu_9983_p1;

assign cipher_0_p16box_address18 = zext_ln587_125_fu_9978_p1;

assign cipher_0_p16box_address19 = zext_ln587_124_fu_9973_p1;

assign cipher_0_p16box_address2 = zext_ln587_141_fu_10813_p1;

assign cipher_0_p16box_address20 = zext_ln587_123_fu_9968_p1;

assign cipher_0_p16box_address21 = zext_ln587_122_fu_9963_p1;

assign cipher_0_p16box_address22 = zext_ln587_121_fu_9958_p1;

assign cipher_0_p16box_address23 = zext_ln587_120_fu_9953_p1;

assign cipher_0_p16box_address24 = zext_ln587_119_fu_9948_p1;

assign cipher_0_p16box_address25 = zext_ln587_118_fu_9943_p1;

assign cipher_0_p16box_address26 = zext_ln587_117_fu_9938_p1;

assign cipher_0_p16box_address27 = zext_ln587_116_fu_9933_p1;

assign cipher_0_p16box_address28 = zext_ln587_115_fu_9928_p1;

assign cipher_0_p16box_address29 = zext_ln587_114_fu_9923_p1;

assign cipher_0_p16box_address3 = zext_ln587_140_fu_10808_p1;

assign cipher_0_p16box_address30 = zext_ln587_113_fu_9918_p1;

assign cipher_0_p16box_address31 = zext_ln587_112_fu_9913_p1;

assign cipher_0_p16box_address32 = zext_ln587_111_fu_9153_p1;

assign cipher_0_p16box_address33 = zext_ln587_110_fu_9148_p1;

assign cipher_0_p16box_address34 = zext_ln587_109_fu_9143_p1;

assign cipher_0_p16box_address35 = zext_ln587_108_fu_9138_p1;

assign cipher_0_p16box_address36 = zext_ln587_107_fu_9133_p1;

assign cipher_0_p16box_address37 = zext_ln587_106_fu_9128_p1;

assign cipher_0_p16box_address38 = zext_ln587_105_fu_9123_p1;

assign cipher_0_p16box_address39 = zext_ln587_104_fu_9118_p1;

assign cipher_0_p16box_address4 = zext_ln587_139_fu_10803_p1;

assign cipher_0_p16box_address40 = zext_ln587_103_fu_9113_p1;

assign cipher_0_p16box_address41 = zext_ln587_102_fu_9108_p1;

assign cipher_0_p16box_address42 = zext_ln587_101_fu_9103_p1;

assign cipher_0_p16box_address43 = zext_ln587_100_fu_9098_p1;

assign cipher_0_p16box_address44 = zext_ln587_99_fu_9093_p1;

assign cipher_0_p16box_address45 = zext_ln587_98_fu_9088_p1;

assign cipher_0_p16box_address46 = zext_ln587_97_fu_9083_p1;

assign cipher_0_p16box_address47 = zext_ln587_96_fu_9078_p1;

assign cipher_0_p16box_address48 = zext_ln587_95_fu_8318_p1;

assign cipher_0_p16box_address49 = zext_ln587_94_fu_8313_p1;

assign cipher_0_p16box_address5 = zext_ln587_138_fu_10798_p1;

assign cipher_0_p16box_address50 = zext_ln587_93_fu_8308_p1;

assign cipher_0_p16box_address51 = zext_ln587_92_fu_8303_p1;

assign cipher_0_p16box_address52 = zext_ln587_91_fu_8298_p1;

assign cipher_0_p16box_address53 = zext_ln587_90_fu_8293_p1;

assign cipher_0_p16box_address54 = zext_ln587_89_fu_8288_p1;

assign cipher_0_p16box_address55 = zext_ln587_88_fu_8283_p1;

assign cipher_0_p16box_address56 = zext_ln587_87_fu_8278_p1;

assign cipher_0_p16box_address57 = zext_ln587_86_fu_8273_p1;

assign cipher_0_p16box_address58 = zext_ln587_85_fu_8268_p1;

assign cipher_0_p16box_address59 = zext_ln587_84_fu_8263_p1;

assign cipher_0_p16box_address6 = zext_ln587_137_fu_10793_p1;

assign cipher_0_p16box_address60 = zext_ln587_83_fu_8258_p1;

assign cipher_0_p16box_address61 = zext_ln587_82_fu_8253_p1;

assign cipher_0_p16box_address62 = zext_ln587_81_fu_8248_p1;

assign cipher_0_p16box_address63 = zext_ln587_80_fu_8243_p1;

assign cipher_0_p16box_address64 = zext_ln587_79_fu_7483_p1;

assign cipher_0_p16box_address65 = zext_ln587_78_fu_7478_p1;

assign cipher_0_p16box_address66 = zext_ln587_77_fu_7473_p1;

assign cipher_0_p16box_address67 = zext_ln587_76_fu_7468_p1;

assign cipher_0_p16box_address68 = zext_ln587_75_fu_7463_p1;

assign cipher_0_p16box_address69 = zext_ln587_74_fu_7458_p1;

assign cipher_0_p16box_address7 = zext_ln587_136_fu_10788_p1;

assign cipher_0_p16box_address70 = zext_ln587_73_fu_7453_p1;

assign cipher_0_p16box_address71 = zext_ln587_72_fu_7448_p1;

assign cipher_0_p16box_address72 = zext_ln587_71_fu_7443_p1;

assign cipher_0_p16box_address73 = zext_ln587_70_fu_7438_p1;

assign cipher_0_p16box_address74 = zext_ln587_69_fu_7433_p1;

assign cipher_0_p16box_address75 = zext_ln587_68_fu_7428_p1;

assign cipher_0_p16box_address76 = zext_ln587_67_fu_7423_p1;

assign cipher_0_p16box_address77 = zext_ln587_66_fu_7418_p1;

assign cipher_0_p16box_address78 = zext_ln587_65_fu_7413_p1;

assign cipher_0_p16box_address79 = zext_ln587_64_fu_7408_p1;

assign cipher_0_p16box_address8 = zext_ln587_135_fu_10783_p1;

assign cipher_0_p16box_address80 = zext_ln587_63_fu_6648_p1;

assign cipher_0_p16box_address81 = zext_ln587_62_fu_6643_p1;

assign cipher_0_p16box_address82 = zext_ln587_61_fu_6638_p1;

assign cipher_0_p16box_address83 = zext_ln587_60_fu_6633_p1;

assign cipher_0_p16box_address84 = zext_ln587_59_fu_6628_p1;

assign cipher_0_p16box_address85 = zext_ln587_58_fu_6623_p1;

assign cipher_0_p16box_address86 = zext_ln587_57_fu_6618_p1;

assign cipher_0_p16box_address87 = zext_ln587_56_fu_6613_p1;

assign cipher_0_p16box_address88 = zext_ln587_55_fu_6608_p1;

assign cipher_0_p16box_address89 = zext_ln587_54_fu_6603_p1;

assign cipher_0_p16box_address9 = zext_ln587_134_fu_10778_p1;

assign cipher_0_p16box_address90 = zext_ln587_53_fu_6598_p1;

assign cipher_0_p16box_address91 = zext_ln587_52_fu_6593_p1;

assign cipher_0_p16box_address92 = zext_ln587_51_fu_6588_p1;

assign cipher_0_p16box_address93 = zext_ln587_50_fu_6583_p1;

assign cipher_0_p16box_address94 = zext_ln587_49_fu_6578_p1;

assign cipher_0_p16box_address95 = zext_ln587_48_fu_6573_p1;

assign cipher_0_p16box_address96 = zext_ln587_47_fu_5813_p1;

assign cipher_0_p16box_address97 = zext_ln587_46_fu_5808_p1;

assign cipher_0_p16box_address98 = zext_ln587_45_fu_5803_p1;

assign cipher_0_p16box_address99 = zext_ln587_44_fu_5798_p1;

assign cipher_0_ssbox_address0 = zext_ln708_162_fu_11578_p1;

assign cipher_0_ssbox_address1 = zext_ln708_161_fu_11563_p1;

assign cipher_0_ssbox_address10 = zext_ln708_152_fu_11428_p1;

assign cipher_0_ssbox_address100 = zext_ln708_62_fu_6508_p1;

assign cipher_0_ssbox_address101 = zext_ln708_61_fu_6493_p1;

assign cipher_0_ssbox_address102 = zext_ln708_60_fu_6478_p1;

assign cipher_0_ssbox_address103 = zext_ln708_59_fu_6463_p1;

assign cipher_0_ssbox_address104 = zext_ln708_58_fu_6448_p1;

assign cipher_0_ssbox_address105 = zext_ln708_57_fu_6433_p1;

assign cipher_0_ssbox_address106 = zext_ln708_56_fu_6418_p1;

assign cipher_0_ssbox_address107 = zext_ln708_55_fu_6403_p1;

assign cipher_0_ssbox_address108 = zext_ln708_54_fu_6388_p1;

assign cipher_0_ssbox_address109 = zext_ln708_53_fu_6373_p1;

assign cipher_0_ssbox_address11 = zext_ln708_151_fu_11413_p1;

assign cipher_0_ssbox_address110 = zext_ln708_52_fu_6358_p1;

assign cipher_0_ssbox_address111 = zext_ln708_51_fu_6343_p1;

assign cipher_0_ssbox_address112 = zext_ln708_50_fu_5733_p1;

assign cipher_0_ssbox_address113 = zext_ln708_49_fu_5718_p1;

assign cipher_0_ssbox_address114 = zext_ln708_48_fu_5703_p1;

assign cipher_0_ssbox_address115 = zext_ln708_47_fu_5688_p1;

assign cipher_0_ssbox_address116 = zext_ln708_46_fu_5673_p1;

assign cipher_0_ssbox_address117 = zext_ln708_45_fu_5658_p1;

assign cipher_0_ssbox_address118 = zext_ln708_44_fu_5643_p1;

assign cipher_0_ssbox_address119 = zext_ln708_43_fu_5628_p1;

assign cipher_0_ssbox_address12 = zext_ln708_150_fu_11398_p1;

assign cipher_0_ssbox_address120 = zext_ln708_42_fu_5613_p1;

assign cipher_0_ssbox_address121 = zext_ln708_41_fu_5598_p1;

assign cipher_0_ssbox_address122 = zext_ln708_40_fu_5583_p1;

assign cipher_0_ssbox_address123 = zext_ln708_39_fu_5568_p1;

assign cipher_0_ssbox_address124 = zext_ln708_38_fu_5553_p1;

assign cipher_0_ssbox_address125 = zext_ln708_37_fu_5538_p1;

assign cipher_0_ssbox_address126 = zext_ln708_36_fu_5523_p1;

assign cipher_0_ssbox_address127 = zext_ln708_35_fu_5508_p1;

assign cipher_0_ssbox_address128 = zext_ln708_34_fu_4898_p1;

assign cipher_0_ssbox_address129 = zext_ln708_33_fu_4883_p1;

assign cipher_0_ssbox_address13 = zext_ln708_149_fu_11383_p1;

assign cipher_0_ssbox_address130 = zext_ln708_32_fu_4868_p1;

assign cipher_0_ssbox_address131 = zext_ln708_31_fu_4853_p1;

assign cipher_0_ssbox_address132 = zext_ln708_30_fu_4838_p1;

assign cipher_0_ssbox_address133 = zext_ln708_29_fu_4823_p1;

assign cipher_0_ssbox_address134 = zext_ln708_28_fu_4808_p1;

assign cipher_0_ssbox_address135 = zext_ln708_27_fu_4793_p1;

assign cipher_0_ssbox_address136 = zext_ln708_26_fu_4778_p1;

assign cipher_0_ssbox_address137 = zext_ln708_25_fu_4763_p1;

assign cipher_0_ssbox_address138 = zext_ln708_24_fu_4748_p1;

assign cipher_0_ssbox_address139 = zext_ln708_23_fu_4733_p1;

assign cipher_0_ssbox_address14 = zext_ln708_148_fu_11368_p1;

assign cipher_0_ssbox_address140 = zext_ln708_22_fu_4718_p1;

assign cipher_0_ssbox_address141 = zext_ln708_21_fu_4703_p1;

assign cipher_0_ssbox_address142 = zext_ln708_20_fu_4688_p1;

assign cipher_0_ssbox_address143 = zext_ln708_19_fu_4673_p1;

assign cipher_0_ssbox_address144 = zext_ln708_18_fu_4063_p1;

assign cipher_0_ssbox_address145 = zext_ln708_17_fu_4048_p1;

assign cipher_0_ssbox_address146 = zext_ln708_16_fu_4033_p1;

assign cipher_0_ssbox_address147 = zext_ln708_15_fu_4018_p1;

assign cipher_0_ssbox_address148 = zext_ln708_14_fu_4003_p1;

assign cipher_0_ssbox_address149 = zext_ln708_13_fu_3988_p1;

assign cipher_0_ssbox_address15 = zext_ln708_147_fu_11353_p1;

assign cipher_0_ssbox_address150 = zext_ln708_12_fu_3973_p1;

assign cipher_0_ssbox_address151 = zext_ln708_11_fu_3958_p1;

assign cipher_0_ssbox_address152 = zext_ln708_10_fu_3943_p1;

assign cipher_0_ssbox_address153 = zext_ln708_9_fu_3928_p1;

assign cipher_0_ssbox_address154 = zext_ln708_8_fu_3913_p1;

assign cipher_0_ssbox_address155 = zext_ln708_7_fu_3898_p1;

assign cipher_0_ssbox_address156 = zext_ln708_6_fu_3883_p1;

assign cipher_0_ssbox_address157 = zext_ln708_5_fu_3868_p1;

assign cipher_0_ssbox_address158 = zext_ln708_4_fu_3853_p1;

assign cipher_0_ssbox_address159 = zext_ln708_fu_3838_p1;

assign cipher_0_ssbox_address16 = zext_ln708_146_fu_10743_p1;

assign cipher_0_ssbox_address17 = zext_ln708_145_fu_10728_p1;

assign cipher_0_ssbox_address18 = zext_ln708_144_fu_10713_p1;

assign cipher_0_ssbox_address19 = zext_ln708_143_fu_10698_p1;

assign cipher_0_ssbox_address2 = zext_ln708_160_fu_11548_p1;

assign cipher_0_ssbox_address20 = zext_ln708_142_fu_10683_p1;

assign cipher_0_ssbox_address21 = zext_ln708_141_fu_10668_p1;

assign cipher_0_ssbox_address22 = zext_ln708_140_fu_10653_p1;

assign cipher_0_ssbox_address23 = zext_ln708_139_fu_10638_p1;

assign cipher_0_ssbox_address24 = zext_ln708_138_fu_10623_p1;

assign cipher_0_ssbox_address25 = zext_ln708_137_fu_10608_p1;

assign cipher_0_ssbox_address26 = zext_ln708_136_fu_10593_p1;

assign cipher_0_ssbox_address27 = zext_ln708_135_fu_10578_p1;

assign cipher_0_ssbox_address28 = zext_ln708_134_fu_10563_p1;

assign cipher_0_ssbox_address29 = zext_ln708_133_fu_10548_p1;

assign cipher_0_ssbox_address3 = zext_ln708_159_fu_11533_p1;

assign cipher_0_ssbox_address30 = zext_ln708_132_fu_10533_p1;

assign cipher_0_ssbox_address31 = zext_ln708_131_fu_10518_p1;

assign cipher_0_ssbox_address32 = zext_ln708_130_fu_9908_p1;

assign cipher_0_ssbox_address33 = zext_ln708_129_fu_9893_p1;

assign cipher_0_ssbox_address34 = zext_ln708_128_fu_9878_p1;

assign cipher_0_ssbox_address35 = zext_ln708_127_fu_9863_p1;

assign cipher_0_ssbox_address36 = zext_ln708_126_fu_9848_p1;

assign cipher_0_ssbox_address37 = zext_ln708_125_fu_9833_p1;

assign cipher_0_ssbox_address38 = zext_ln708_124_fu_9818_p1;

assign cipher_0_ssbox_address39 = zext_ln708_123_fu_9803_p1;

assign cipher_0_ssbox_address4 = zext_ln708_158_fu_11518_p1;

assign cipher_0_ssbox_address40 = zext_ln708_122_fu_9788_p1;

assign cipher_0_ssbox_address41 = zext_ln708_121_fu_9773_p1;

assign cipher_0_ssbox_address42 = zext_ln708_120_fu_9758_p1;

assign cipher_0_ssbox_address43 = zext_ln708_119_fu_9743_p1;

assign cipher_0_ssbox_address44 = zext_ln708_118_fu_9728_p1;

assign cipher_0_ssbox_address45 = zext_ln708_117_fu_9713_p1;

assign cipher_0_ssbox_address46 = zext_ln708_116_fu_9698_p1;

assign cipher_0_ssbox_address47 = zext_ln708_115_fu_9683_p1;

assign cipher_0_ssbox_address48 = zext_ln708_114_fu_9073_p1;

assign cipher_0_ssbox_address49 = zext_ln708_113_fu_9058_p1;

assign cipher_0_ssbox_address5 = zext_ln708_157_fu_11503_p1;

assign cipher_0_ssbox_address50 = zext_ln708_112_fu_9043_p1;

assign cipher_0_ssbox_address51 = zext_ln708_111_fu_9028_p1;

assign cipher_0_ssbox_address52 = zext_ln708_110_fu_9013_p1;

assign cipher_0_ssbox_address53 = zext_ln708_109_fu_8998_p1;

assign cipher_0_ssbox_address54 = zext_ln708_108_fu_8983_p1;

assign cipher_0_ssbox_address55 = zext_ln708_107_fu_8968_p1;

assign cipher_0_ssbox_address56 = zext_ln708_106_fu_8953_p1;

assign cipher_0_ssbox_address57 = zext_ln708_105_fu_8938_p1;

assign cipher_0_ssbox_address58 = zext_ln708_104_fu_8923_p1;

assign cipher_0_ssbox_address59 = zext_ln708_103_fu_8908_p1;

assign cipher_0_ssbox_address6 = zext_ln708_156_fu_11488_p1;

assign cipher_0_ssbox_address60 = zext_ln708_102_fu_8893_p1;

assign cipher_0_ssbox_address61 = zext_ln708_101_fu_8878_p1;

assign cipher_0_ssbox_address62 = zext_ln708_100_fu_8863_p1;

assign cipher_0_ssbox_address63 = zext_ln708_99_fu_8848_p1;

assign cipher_0_ssbox_address64 = zext_ln708_98_fu_8238_p1;

assign cipher_0_ssbox_address65 = zext_ln708_97_fu_8223_p1;

assign cipher_0_ssbox_address66 = zext_ln708_96_fu_8208_p1;

assign cipher_0_ssbox_address67 = zext_ln708_95_fu_8193_p1;

assign cipher_0_ssbox_address68 = zext_ln708_94_fu_8178_p1;

assign cipher_0_ssbox_address69 = zext_ln708_93_fu_8163_p1;

assign cipher_0_ssbox_address7 = zext_ln708_155_fu_11473_p1;

assign cipher_0_ssbox_address70 = zext_ln708_92_fu_8148_p1;

assign cipher_0_ssbox_address71 = zext_ln708_91_fu_8133_p1;

assign cipher_0_ssbox_address72 = zext_ln708_90_fu_8118_p1;

assign cipher_0_ssbox_address73 = zext_ln708_89_fu_8103_p1;

assign cipher_0_ssbox_address74 = zext_ln708_88_fu_8088_p1;

assign cipher_0_ssbox_address75 = zext_ln708_87_fu_8073_p1;

assign cipher_0_ssbox_address76 = zext_ln708_86_fu_8058_p1;

assign cipher_0_ssbox_address77 = zext_ln708_85_fu_8043_p1;

assign cipher_0_ssbox_address78 = zext_ln708_84_fu_8028_p1;

assign cipher_0_ssbox_address79 = zext_ln708_83_fu_8013_p1;

assign cipher_0_ssbox_address8 = zext_ln708_154_fu_11458_p1;

assign cipher_0_ssbox_address80 = zext_ln708_82_fu_7403_p1;

assign cipher_0_ssbox_address81 = zext_ln708_81_fu_7388_p1;

assign cipher_0_ssbox_address82 = zext_ln708_80_fu_7373_p1;

assign cipher_0_ssbox_address83 = zext_ln708_79_fu_7358_p1;

assign cipher_0_ssbox_address84 = zext_ln708_78_fu_7343_p1;

assign cipher_0_ssbox_address85 = zext_ln708_77_fu_7328_p1;

assign cipher_0_ssbox_address86 = zext_ln708_76_fu_7313_p1;

assign cipher_0_ssbox_address87 = zext_ln708_75_fu_7298_p1;

assign cipher_0_ssbox_address88 = zext_ln708_74_fu_7283_p1;

assign cipher_0_ssbox_address89 = zext_ln708_73_fu_7268_p1;

assign cipher_0_ssbox_address9 = zext_ln708_153_fu_11443_p1;

assign cipher_0_ssbox_address90 = zext_ln708_72_fu_7253_p1;

assign cipher_0_ssbox_address91 = zext_ln708_71_fu_7238_p1;

assign cipher_0_ssbox_address92 = zext_ln708_70_fu_7223_p1;

assign cipher_0_ssbox_address93 = zext_ln708_69_fu_7208_p1;

assign cipher_0_ssbox_address94 = zext_ln708_68_fu_7193_p1;

assign cipher_0_ssbox_address95 = zext_ln708_67_fu_7178_p1;

assign cipher_0_ssbox_address96 = zext_ln708_66_fu_6568_p1;

assign cipher_0_ssbox_address97 = zext_ln708_65_fu_6553_p1;

assign cipher_0_ssbox_address98 = zext_ln708_64_fu_6538_p1;

assign cipher_0_ssbox_address99 = zext_ln708_63_fu_6523_p1;

assign p_Result_10_fu_11583_p17 = {{{{{{{{{{{{{{{{cipher_0_ssbox_q4}, {cipher_0_ssbox_q9}}, {cipher_0_ssbox_q14}}, {cipher_0_ssbox_q3}}, {cipher_0_ssbox_q8}}, {cipher_0_ssbox_q13}}, {cipher_0_ssbox_q2}}, {cipher_0_ssbox_q7}}, {cipher_0_ssbox_q12}}, {cipher_0_ssbox_q1}}, {cipher_0_ssbox_q6}}, {cipher_0_ssbox_q11}}, {cipher_0_ssbox_q0}}, {cipher_0_ssbox_q5}}, {cipher_0_ssbox_q10}}, {cipher_0_ssbox_q15}};

assign p_Result_2_fu_5463_p17 = {{{{{{{{{{{{{{{{xor_ln1545_98_fu_5457_p2}, {xor_ln1545_95_fu_5441_p2}}, {xor_ln1545_92_fu_5425_p2}}, {xor_ln1545_89_fu_5409_p2}}, {xor_ln1545_86_fu_5393_p2}}, {xor_ln1545_83_fu_5377_p2}}, {xor_ln1545_80_fu_5361_p2}}, {xor_ln1545_77_fu_5345_p2}}, {xor_ln1545_74_fu_5329_p2}}, {xor_ln1545_71_fu_5313_p2}}, {xor_ln1545_68_fu_5297_p2}}, {xor_ln1545_65_fu_5281_p2}}, {xor_ln1545_62_fu_5265_p2}}, {xor_ln1545_59_fu_5249_p2}}, {xor_ln1545_56_fu_5233_p2}}, {xor_ln1545_53_fu_5217_p2}};

assign p_Result_3_fu_6298_p17 = {{{{{{{{{{{{{{{{xor_ln1545_146_fu_6292_p2}, {xor_ln1545_143_fu_6276_p2}}, {xor_ln1545_140_fu_6260_p2}}, {xor_ln1545_137_fu_6244_p2}}, {xor_ln1545_134_fu_6228_p2}}, {xor_ln1545_131_fu_6212_p2}}, {xor_ln1545_128_fu_6196_p2}}, {xor_ln1545_125_fu_6180_p2}}, {xor_ln1545_122_fu_6164_p2}}, {xor_ln1545_119_fu_6148_p2}}, {xor_ln1545_116_fu_6132_p2}}, {xor_ln1545_113_fu_6116_p2}}, {xor_ln1545_110_fu_6100_p2}}, {xor_ln1545_107_fu_6084_p2}}, {xor_ln1545_104_fu_6068_p2}}, {xor_ln1545_101_fu_6052_p2}};

assign p_Result_4_fu_7133_p17 = {{{{{{{{{{{{{{{{xor_ln1545_194_fu_7127_p2}, {xor_ln1545_191_fu_7111_p2}}, {xor_ln1545_188_fu_7095_p2}}, {xor_ln1545_185_fu_7079_p2}}, {xor_ln1545_182_fu_7063_p2}}, {xor_ln1545_179_fu_7047_p2}}, {xor_ln1545_176_fu_7031_p2}}, {xor_ln1545_173_fu_7015_p2}}, {xor_ln1545_170_fu_6999_p2}}, {xor_ln1545_167_fu_6983_p2}}, {xor_ln1545_164_fu_6967_p2}}, {xor_ln1545_161_fu_6951_p2}}, {xor_ln1545_158_fu_6935_p2}}, {xor_ln1545_155_fu_6919_p2}}, {xor_ln1545_152_fu_6903_p2}}, {xor_ln1545_149_fu_6887_p2}};

assign p_Result_5_fu_7968_p17 = {{{{{{{{{{{{{{{{xor_ln1545_242_fu_7962_p2}, {xor_ln1545_239_fu_7946_p2}}, {xor_ln1545_236_fu_7930_p2}}, {xor_ln1545_233_fu_7914_p2}}, {xor_ln1545_230_fu_7898_p2}}, {xor_ln1545_227_fu_7882_p2}}, {xor_ln1545_224_fu_7866_p2}}, {xor_ln1545_221_fu_7850_p2}}, {xor_ln1545_218_fu_7834_p2}}, {xor_ln1545_215_fu_7818_p2}}, {xor_ln1545_212_fu_7802_p2}}, {xor_ln1545_209_fu_7786_p2}}, {xor_ln1545_206_fu_7770_p2}}, {xor_ln1545_203_fu_7754_p2}}, {xor_ln1545_200_fu_7738_p2}}, {xor_ln1545_197_fu_7722_p2}};

assign p_Result_6_fu_8803_p17 = {{{{{{{{{{{{{{{{xor_ln1545_290_fu_8797_p2}, {xor_ln1545_287_fu_8781_p2}}, {xor_ln1545_284_fu_8765_p2}}, {xor_ln1545_281_fu_8749_p2}}, {xor_ln1545_278_fu_8733_p2}}, {xor_ln1545_275_fu_8717_p2}}, {xor_ln1545_272_fu_8701_p2}}, {xor_ln1545_269_fu_8685_p2}}, {xor_ln1545_266_fu_8669_p2}}, {xor_ln1545_263_fu_8653_p2}}, {xor_ln1545_260_fu_8637_p2}}, {xor_ln1545_257_fu_8621_p2}}, {xor_ln1545_254_fu_8605_p2}}, {xor_ln1545_251_fu_8589_p2}}, {xor_ln1545_248_fu_8573_p2}}, {xor_ln1545_245_fu_8557_p2}};

assign p_Result_7_fu_9638_p17 = {{{{{{{{{{{{{{{{xor_ln1545_338_fu_9632_p2}, {xor_ln1545_335_fu_9616_p2}}, {xor_ln1545_332_fu_9600_p2}}, {xor_ln1545_329_fu_9584_p2}}, {xor_ln1545_326_fu_9568_p2}}, {xor_ln1545_323_fu_9552_p2}}, {xor_ln1545_320_fu_9536_p2}}, {xor_ln1545_317_fu_9520_p2}}, {xor_ln1545_314_fu_9504_p2}}, {xor_ln1545_311_fu_9488_p2}}, {xor_ln1545_308_fu_9472_p2}}, {xor_ln1545_305_fu_9456_p2}}, {xor_ln1545_302_fu_9440_p2}}, {xor_ln1545_299_fu_9424_p2}}, {xor_ln1545_296_fu_9408_p2}}, {xor_ln1545_293_fu_9392_p2}};

assign p_Result_8_fu_10473_p17 = {{{{{{{{{{{{{{{{xor_ln1545_386_fu_10467_p2}, {xor_ln1545_383_fu_10451_p2}}, {xor_ln1545_380_fu_10435_p2}}, {xor_ln1545_377_fu_10419_p2}}, {xor_ln1545_374_fu_10403_p2}}, {xor_ln1545_371_fu_10387_p2}}, {xor_ln1545_368_fu_10371_p2}}, {xor_ln1545_365_fu_10355_p2}}, {xor_ln1545_362_fu_10339_p2}}, {xor_ln1545_359_fu_10323_p2}}, {xor_ln1545_356_fu_10307_p2}}, {xor_ln1545_353_fu_10291_p2}}, {xor_ln1545_350_fu_10275_p2}}, {xor_ln1545_347_fu_10259_p2}}, {xor_ln1545_344_fu_10243_p2}}, {xor_ln1545_341_fu_10227_p2}};

assign p_Result_9_fu_11308_p17 = {{{{{{{{{{{{{{{{xor_ln1545_434_fu_11302_p2}, {xor_ln1545_431_fu_11286_p2}}, {xor_ln1545_428_fu_11270_p2}}, {xor_ln1545_425_fu_11254_p2}}, {xor_ln1545_422_fu_11238_p2}}, {xor_ln1545_419_fu_11222_p2}}, {xor_ln1545_416_fu_11206_p2}}, {xor_ln1545_413_fu_11190_p2}}, {xor_ln1545_410_fu_11174_p2}}, {xor_ln1545_407_fu_11158_p2}}, {xor_ln1545_404_fu_11142_p2}}, {xor_ln1545_401_fu_11126_p2}}, {xor_ln1545_398_fu_11110_p2}}, {xor_ln1545_395_fu_11094_p2}}, {xor_ln1545_392_fu_11078_p2}}, {xor_ln1545_389_fu_11062_p2}};

assign p_Result_s_fu_4628_p17 = {{{{{{{{{{{{{{{{xor_ln1545_50_fu_4622_p2}, {xor_ln1545_47_fu_4606_p2}}, {xor_ln1545_44_fu_4590_p2}}, {xor_ln1545_41_fu_4574_p2}}, {xor_ln1545_38_fu_4558_p2}}, {xor_ln1545_35_fu_4542_p2}}, {xor_ln1545_32_fu_4526_p2}}, {xor_ln1545_29_fu_4510_p2}}, {xor_ln1545_26_fu_4494_p2}}, {xor_ln1545_23_fu_4478_p2}}, {xor_ln1545_20_fu_4462_p2}}, {xor_ln1545_17_fu_4446_p2}}, {xor_ln1545_14_fu_4430_p2}}, {xor_ln1545_11_fu_4414_p2}}, {xor_ln1545_8_fu_4398_p2}}, {xor_ln1545_5_fu_4382_p2}};

assign ret_V_fu_3828_p2 = (plaintext ^ p_read);

assign state_V_20_fu_4664_p2 = (p_read_10_reg_11669_pp0_iter1_reg ^ p_Result_s_fu_4628_p17);

assign state_V_21_fu_5499_p2 = (p_read_9_reg_11664_pp0_iter3_reg ^ p_Result_2_fu_5463_p17);

assign state_V_22_fu_6334_p2 = (p_read_8_reg_11659_pp0_iter5_reg ^ p_Result_3_fu_6298_p17);

assign state_V_23_fu_7169_p2 = (p_read_7_reg_11654_pp0_iter7_reg ^ p_Result_4_fu_7133_p17);

assign state_V_24_fu_8004_p2 = (p_read_6_reg_11649_pp0_iter9_reg ^ p_Result_5_fu_7968_p17);

assign state_V_25_fu_8839_p2 = (p_read_5_reg_11644_pp0_iter11_reg ^ p_Result_6_fu_8803_p17);

assign state_V_26_fu_10509_p2 = (p_read_3_reg_11634_pp0_iter15_reg ^ p_Result_8_fu_10473_p17);

assign state_V_27_fu_11344_p2 = (p_read_2_reg_11629_pp0_iter17_reg ^ p_Result_9_fu_11308_p17);

assign state_V_fu_9674_p2 = (p_read_4_reg_11639_pp0_iter13_reg ^ p_Result_7_fu_9638_p17);

assign tmp_100_fu_6408_p4 = {{state_V_22_fu_6334_p2[47:40]}};

assign tmp_101_fu_6423_p4 = {{state_V_22_fu_6334_p2[55:48]}};

assign tmp_102_fu_6438_p4 = {{state_V_22_fu_6334_p2[63:56]}};

assign tmp_103_fu_6453_p4 = {{state_V_22_fu_6334_p2[71:64]}};

assign tmp_104_fu_6468_p4 = {{state_V_22_fu_6334_p2[79:72]}};

assign tmp_105_fu_6483_p4 = {{state_V_22_fu_6334_p2[87:80]}};

assign tmp_106_fu_6498_p4 = {{state_V_22_fu_6334_p2[95:88]}};

assign tmp_107_fu_6513_p4 = {{state_V_22_fu_6334_p2[103:96]}};

assign tmp_108_fu_6528_p4 = {{state_V_22_fu_6334_p2[111:104]}};

assign tmp_109_fu_6543_p4 = {{state_V_22_fu_6334_p2[119:112]}};

assign tmp_10_fu_3948_p4 = {{ret_V_fu_3828_p2[71:64]}};

assign tmp_110_fu_6558_p4 = {{state_V_22_fu_6334_p2[127:120]}};

assign tmp_111_fu_6657_p4 = {{cipher_0_p16box_q95[15:8]}};

assign tmp_112_fu_6671_p4 = {{cipher_0_p16box_q94[15:8]}};

assign tmp_113_fu_6685_p4 = {{cipher_0_p16box_q93[15:8]}};

assign tmp_114_fu_6699_p4 = {{cipher_0_p16box_q92[15:8]}};

assign tmp_115_fu_6713_p4 = {{cipher_0_p16box_q91[15:8]}};

assign tmp_116_fu_6727_p4 = {{cipher_0_p16box_q90[15:8]}};

assign tmp_117_fu_6741_p4 = {{cipher_0_p16box_q89[15:8]}};

assign tmp_118_fu_6755_p4 = {{cipher_0_p16box_q88[15:8]}};

assign tmp_119_fu_6769_p4 = {{cipher_0_p16box_q87[15:8]}};

assign tmp_11_fu_3963_p4 = {{ret_V_fu_3828_p2[79:72]}};

assign tmp_120_fu_6783_p4 = {{cipher_0_p16box_q86[15:8]}};

assign tmp_121_fu_6797_p4 = {{cipher_0_p16box_q85[15:8]}};

assign tmp_122_fu_6811_p4 = {{cipher_0_p16box_q84[15:8]}};

assign tmp_123_fu_6825_p4 = {{cipher_0_p16box_q83[15:8]}};

assign tmp_124_fu_6839_p4 = {{cipher_0_p16box_q82[15:8]}};

assign tmp_125_fu_6853_p4 = {{cipher_0_p16box_q81[15:8]}};

assign tmp_126_fu_6867_p4 = {{cipher_0_p16box_q80[15:8]}};

assign tmp_127_fu_7183_p4 = {{state_V_23_fu_7169_p2[15:8]}};

assign tmp_128_fu_7198_p4 = {{state_V_23_fu_7169_p2[23:16]}};

assign tmp_129_fu_7213_p4 = {{state_V_23_fu_7169_p2[31:24]}};

assign tmp_12_fu_3978_p4 = {{ret_V_fu_3828_p2[87:80]}};

assign tmp_130_fu_7228_p4 = {{state_V_23_fu_7169_p2[39:32]}};

assign tmp_131_fu_7243_p4 = {{state_V_23_fu_7169_p2[47:40]}};

assign tmp_132_fu_7258_p4 = {{state_V_23_fu_7169_p2[55:48]}};

assign tmp_133_fu_7273_p4 = {{state_V_23_fu_7169_p2[63:56]}};

assign tmp_134_fu_7288_p4 = {{state_V_23_fu_7169_p2[71:64]}};

assign tmp_135_fu_7303_p4 = {{state_V_23_fu_7169_p2[79:72]}};

assign tmp_136_fu_7318_p4 = {{state_V_23_fu_7169_p2[87:80]}};

assign tmp_137_fu_7333_p4 = {{state_V_23_fu_7169_p2[95:88]}};

assign tmp_138_fu_7348_p4 = {{state_V_23_fu_7169_p2[103:96]}};

assign tmp_139_fu_7363_p4 = {{state_V_23_fu_7169_p2[111:104]}};

assign tmp_13_fu_3993_p4 = {{ret_V_fu_3828_p2[95:88]}};

assign tmp_140_fu_7378_p4 = {{state_V_23_fu_7169_p2[119:112]}};

assign tmp_141_fu_7393_p4 = {{state_V_23_fu_7169_p2[127:120]}};

assign tmp_142_fu_7492_p4 = {{cipher_0_p16box_q79[15:8]}};

assign tmp_143_fu_7506_p4 = {{cipher_0_p16box_q78[15:8]}};

assign tmp_144_fu_7520_p4 = {{cipher_0_p16box_q77[15:8]}};

assign tmp_145_fu_7534_p4 = {{cipher_0_p16box_q76[15:8]}};

assign tmp_146_fu_7548_p4 = {{cipher_0_p16box_q75[15:8]}};

assign tmp_147_fu_7562_p4 = {{cipher_0_p16box_q74[15:8]}};

assign tmp_148_fu_7576_p4 = {{cipher_0_p16box_q73[15:8]}};

assign tmp_149_fu_7590_p4 = {{cipher_0_p16box_q72[15:8]}};

assign tmp_14_fu_4008_p4 = {{ret_V_fu_3828_p2[103:96]}};

assign tmp_150_fu_7604_p4 = {{cipher_0_p16box_q71[15:8]}};

assign tmp_151_fu_7618_p4 = {{cipher_0_p16box_q70[15:8]}};

assign tmp_152_fu_7632_p4 = {{cipher_0_p16box_q69[15:8]}};

assign tmp_153_fu_7646_p4 = {{cipher_0_p16box_q68[15:8]}};

assign tmp_154_fu_7660_p4 = {{cipher_0_p16box_q67[15:8]}};

assign tmp_155_fu_7674_p4 = {{cipher_0_p16box_q66[15:8]}};

assign tmp_156_fu_7688_p4 = {{cipher_0_p16box_q65[15:8]}};

assign tmp_157_fu_7702_p4 = {{cipher_0_p16box_q64[15:8]}};

assign tmp_158_fu_8018_p4 = {{state_V_24_fu_8004_p2[15:8]}};

assign tmp_159_fu_8033_p4 = {{state_V_24_fu_8004_p2[23:16]}};

assign tmp_15_fu_4023_p4 = {{ret_V_fu_3828_p2[111:104]}};

assign tmp_160_fu_8048_p4 = {{state_V_24_fu_8004_p2[31:24]}};

assign tmp_161_fu_8063_p4 = {{state_V_24_fu_8004_p2[39:32]}};

assign tmp_162_fu_8078_p4 = {{state_V_24_fu_8004_p2[47:40]}};

assign tmp_163_fu_8093_p4 = {{state_V_24_fu_8004_p2[55:48]}};

assign tmp_164_fu_8108_p4 = {{state_V_24_fu_8004_p2[63:56]}};

assign tmp_165_fu_8123_p4 = {{state_V_24_fu_8004_p2[71:64]}};

assign tmp_166_fu_8138_p4 = {{state_V_24_fu_8004_p2[79:72]}};

assign tmp_167_fu_8153_p4 = {{state_V_24_fu_8004_p2[87:80]}};

assign tmp_168_fu_8168_p4 = {{state_V_24_fu_8004_p2[95:88]}};

assign tmp_169_fu_8183_p4 = {{state_V_24_fu_8004_p2[103:96]}};

assign tmp_16_fu_4038_p4 = {{ret_V_fu_3828_p2[119:112]}};

assign tmp_170_fu_8198_p4 = {{state_V_24_fu_8004_p2[111:104]}};

assign tmp_171_fu_8213_p4 = {{state_V_24_fu_8004_p2[119:112]}};

assign tmp_172_fu_8228_p4 = {{state_V_24_fu_8004_p2[127:120]}};

assign tmp_173_fu_8327_p4 = {{cipher_0_p16box_q63[15:8]}};

assign tmp_174_fu_8341_p4 = {{cipher_0_p16box_q62[15:8]}};

assign tmp_175_fu_8355_p4 = {{cipher_0_p16box_q61[15:8]}};

assign tmp_176_fu_8369_p4 = {{cipher_0_p16box_q60[15:8]}};

assign tmp_177_fu_8383_p4 = {{cipher_0_p16box_q59[15:8]}};

assign tmp_178_fu_8397_p4 = {{cipher_0_p16box_q58[15:8]}};

assign tmp_179_fu_8411_p4 = {{cipher_0_p16box_q57[15:8]}};

assign tmp_17_fu_4053_p4 = {{ret_V_fu_3828_p2[127:120]}};

assign tmp_180_fu_8425_p4 = {{cipher_0_p16box_q56[15:8]}};

assign tmp_181_fu_8439_p4 = {{cipher_0_p16box_q55[15:8]}};

assign tmp_182_fu_8453_p4 = {{cipher_0_p16box_q54[15:8]}};

assign tmp_183_fu_8467_p4 = {{cipher_0_p16box_q53[15:8]}};

assign tmp_184_fu_8481_p4 = {{cipher_0_p16box_q52[15:8]}};

assign tmp_185_fu_8495_p4 = {{cipher_0_p16box_q51[15:8]}};

assign tmp_186_fu_8509_p4 = {{cipher_0_p16box_q50[15:8]}};

assign tmp_187_fu_8523_p4 = {{cipher_0_p16box_q49[15:8]}};

assign tmp_188_fu_8537_p4 = {{cipher_0_p16box_q48[15:8]}};

assign tmp_189_fu_8853_p4 = {{state_V_25_fu_8839_p2[15:8]}};

assign tmp_18_fu_4152_p4 = {{cipher_0_p16box_q143[15:8]}};

assign tmp_190_fu_8868_p4 = {{state_V_25_fu_8839_p2[23:16]}};

assign tmp_191_fu_8883_p4 = {{state_V_25_fu_8839_p2[31:24]}};

assign tmp_192_fu_8898_p4 = {{state_V_25_fu_8839_p2[39:32]}};

assign tmp_193_fu_8913_p4 = {{state_V_25_fu_8839_p2[47:40]}};

assign tmp_194_fu_8928_p4 = {{state_V_25_fu_8839_p2[55:48]}};

assign tmp_195_fu_8943_p4 = {{state_V_25_fu_8839_p2[63:56]}};

assign tmp_196_fu_8958_p4 = {{state_V_25_fu_8839_p2[71:64]}};

assign tmp_197_fu_8973_p4 = {{state_V_25_fu_8839_p2[79:72]}};

assign tmp_198_fu_8988_p4 = {{state_V_25_fu_8839_p2[87:80]}};

assign tmp_199_fu_9003_p4 = {{state_V_25_fu_8839_p2[95:88]}};

assign tmp_19_fu_4166_p4 = {{cipher_0_p16box_q142[15:8]}};

assign tmp_200_fu_9018_p4 = {{state_V_25_fu_8839_p2[103:96]}};

assign tmp_201_fu_9033_p4 = {{state_V_25_fu_8839_p2[111:104]}};

assign tmp_202_fu_9048_p4 = {{state_V_25_fu_8839_p2[119:112]}};

assign tmp_203_fu_9063_p4 = {{state_V_25_fu_8839_p2[127:120]}};

assign tmp_204_fu_9162_p4 = {{cipher_0_p16box_q47[15:8]}};

assign tmp_205_fu_9176_p4 = {{cipher_0_p16box_q46[15:8]}};

assign tmp_206_fu_9190_p4 = {{cipher_0_p16box_q45[15:8]}};

assign tmp_207_fu_9204_p4 = {{cipher_0_p16box_q44[15:8]}};

assign tmp_208_fu_9218_p4 = {{cipher_0_p16box_q43[15:8]}};

assign tmp_209_fu_9232_p4 = {{cipher_0_p16box_q42[15:8]}};

assign tmp_20_fu_4180_p4 = {{cipher_0_p16box_q141[15:8]}};

assign tmp_210_fu_9246_p4 = {{cipher_0_p16box_q41[15:8]}};

assign tmp_211_fu_9260_p4 = {{cipher_0_p16box_q40[15:8]}};

assign tmp_212_fu_9274_p4 = {{cipher_0_p16box_q39[15:8]}};

assign tmp_213_fu_9288_p4 = {{cipher_0_p16box_q38[15:8]}};

assign tmp_214_fu_9302_p4 = {{cipher_0_p16box_q37[15:8]}};

assign tmp_215_fu_9316_p4 = {{cipher_0_p16box_q36[15:8]}};

assign tmp_216_fu_9330_p4 = {{cipher_0_p16box_q35[15:8]}};

assign tmp_217_fu_9344_p4 = {{cipher_0_p16box_q34[15:8]}};

assign tmp_218_fu_9358_p4 = {{cipher_0_p16box_q33[15:8]}};

assign tmp_219_fu_9372_p4 = {{cipher_0_p16box_q32[15:8]}};

assign tmp_21_fu_4194_p4 = {{cipher_0_p16box_q140[15:8]}};

assign tmp_220_fu_9688_p4 = {{state_V_fu_9674_p2[15:8]}};

assign tmp_221_fu_9703_p4 = {{state_V_fu_9674_p2[23:16]}};

assign tmp_222_fu_9718_p4 = {{state_V_fu_9674_p2[31:24]}};

assign tmp_223_fu_9733_p4 = {{state_V_fu_9674_p2[39:32]}};

assign tmp_224_fu_9748_p4 = {{state_V_fu_9674_p2[47:40]}};

assign tmp_225_fu_9763_p4 = {{state_V_fu_9674_p2[55:48]}};

assign tmp_226_fu_9778_p4 = {{state_V_fu_9674_p2[63:56]}};

assign tmp_227_fu_9793_p4 = {{state_V_fu_9674_p2[71:64]}};

assign tmp_228_fu_9808_p4 = {{state_V_fu_9674_p2[79:72]}};

assign tmp_229_fu_9823_p4 = {{state_V_fu_9674_p2[87:80]}};

assign tmp_22_fu_4208_p4 = {{cipher_0_p16box_q139[15:8]}};

assign tmp_230_fu_9838_p4 = {{state_V_fu_9674_p2[95:88]}};

assign tmp_231_fu_9853_p4 = {{state_V_fu_9674_p2[103:96]}};

assign tmp_232_fu_9868_p4 = {{state_V_fu_9674_p2[111:104]}};

assign tmp_233_fu_9883_p4 = {{state_V_fu_9674_p2[119:112]}};

assign tmp_234_fu_9898_p4 = {{state_V_fu_9674_p2[127:120]}};

assign tmp_235_fu_9997_p4 = {{cipher_0_p16box_q31[15:8]}};

assign tmp_236_fu_10011_p4 = {{cipher_0_p16box_q30[15:8]}};

assign tmp_237_fu_10025_p4 = {{cipher_0_p16box_q29[15:8]}};

assign tmp_238_fu_10039_p4 = {{cipher_0_p16box_q28[15:8]}};

assign tmp_239_fu_10053_p4 = {{cipher_0_p16box_q27[15:8]}};

assign tmp_23_fu_4222_p4 = {{cipher_0_p16box_q138[15:8]}};

assign tmp_240_fu_10067_p4 = {{cipher_0_p16box_q26[15:8]}};

assign tmp_241_fu_10081_p4 = {{cipher_0_p16box_q25[15:8]}};

assign tmp_242_fu_10095_p4 = {{cipher_0_p16box_q24[15:8]}};

assign tmp_243_fu_10109_p4 = {{cipher_0_p16box_q23[15:8]}};

assign tmp_244_fu_10123_p4 = {{cipher_0_p16box_q22[15:8]}};

assign tmp_245_fu_10137_p4 = {{cipher_0_p16box_q21[15:8]}};

assign tmp_246_fu_10151_p4 = {{cipher_0_p16box_q20[15:8]}};

assign tmp_247_fu_10165_p4 = {{cipher_0_p16box_q19[15:8]}};

assign tmp_248_fu_10179_p4 = {{cipher_0_p16box_q18[15:8]}};

assign tmp_249_fu_10193_p4 = {{cipher_0_p16box_q17[15:8]}};

assign tmp_24_fu_4236_p4 = {{cipher_0_p16box_q137[15:8]}};

assign tmp_250_fu_10207_p4 = {{cipher_0_p16box_q16[15:8]}};

assign tmp_251_fu_10523_p4 = {{state_V_26_fu_10509_p2[15:8]}};

assign tmp_252_fu_10538_p4 = {{state_V_26_fu_10509_p2[23:16]}};

assign tmp_253_fu_10553_p4 = {{state_V_26_fu_10509_p2[31:24]}};

assign tmp_254_fu_10568_p4 = {{state_V_26_fu_10509_p2[39:32]}};

assign tmp_255_fu_10583_p4 = {{state_V_26_fu_10509_p2[47:40]}};

assign tmp_256_fu_10598_p4 = {{state_V_26_fu_10509_p2[55:48]}};

assign tmp_257_fu_10613_p4 = {{state_V_26_fu_10509_p2[63:56]}};

assign tmp_258_fu_10628_p4 = {{state_V_26_fu_10509_p2[71:64]}};

assign tmp_259_fu_10643_p4 = {{state_V_26_fu_10509_p2[79:72]}};

assign tmp_25_fu_4250_p4 = {{cipher_0_p16box_q136[15:8]}};

assign tmp_260_fu_10658_p4 = {{state_V_26_fu_10509_p2[87:80]}};

assign tmp_261_fu_10673_p4 = {{state_V_26_fu_10509_p2[95:88]}};

assign tmp_262_fu_10688_p4 = {{state_V_26_fu_10509_p2[103:96]}};

assign tmp_263_fu_10703_p4 = {{state_V_26_fu_10509_p2[111:104]}};

assign tmp_264_fu_10718_p4 = {{state_V_26_fu_10509_p2[119:112]}};

assign tmp_265_fu_10733_p4 = {{state_V_26_fu_10509_p2[127:120]}};

assign tmp_266_fu_10832_p4 = {{cipher_0_p16box_q15[15:8]}};

assign tmp_267_fu_10846_p4 = {{cipher_0_p16box_q14[15:8]}};

assign tmp_268_fu_10860_p4 = {{cipher_0_p16box_q13[15:8]}};

assign tmp_269_fu_10874_p4 = {{cipher_0_p16box_q12[15:8]}};

assign tmp_26_fu_4264_p4 = {{cipher_0_p16box_q135[15:8]}};

assign tmp_270_fu_10888_p4 = {{cipher_0_p16box_q11[15:8]}};

assign tmp_271_fu_10902_p4 = {{cipher_0_p16box_q10[15:8]}};

assign tmp_272_fu_10916_p4 = {{cipher_0_p16box_q9[15:8]}};

assign tmp_273_fu_10930_p4 = {{cipher_0_p16box_q8[15:8]}};

assign tmp_274_fu_10944_p4 = {{cipher_0_p16box_q7[15:8]}};

assign tmp_275_fu_10958_p4 = {{cipher_0_p16box_q6[15:8]}};

assign tmp_276_fu_10972_p4 = {{cipher_0_p16box_q5[15:8]}};

assign tmp_277_fu_10986_p4 = {{cipher_0_p16box_q4[15:8]}};

assign tmp_278_fu_11000_p4 = {{cipher_0_p16box_q3[15:8]}};

assign tmp_279_fu_11014_p4 = {{cipher_0_p16box_q2[15:8]}};

assign tmp_27_fu_4278_p4 = {{cipher_0_p16box_q134[15:8]}};

assign tmp_280_fu_11028_p4 = {{cipher_0_p16box_q1[15:8]}};

assign tmp_281_fu_11042_p4 = {{cipher_0_p16box_q0[15:8]}};

assign tmp_282_fu_11358_p4 = {{state_V_27_fu_11344_p2[15:8]}};

assign tmp_283_fu_11373_p4 = {{state_V_27_fu_11344_p2[23:16]}};

assign tmp_284_fu_11388_p4 = {{state_V_27_fu_11344_p2[31:24]}};

assign tmp_285_fu_11403_p4 = {{state_V_27_fu_11344_p2[39:32]}};

assign tmp_286_fu_11418_p4 = {{state_V_27_fu_11344_p2[47:40]}};

assign tmp_287_fu_11433_p4 = {{state_V_27_fu_11344_p2[55:48]}};

assign tmp_288_fu_11448_p4 = {{state_V_27_fu_11344_p2[63:56]}};

assign tmp_289_fu_11463_p4 = {{state_V_27_fu_11344_p2[71:64]}};

assign tmp_28_fu_4292_p4 = {{cipher_0_p16box_q133[15:8]}};

assign tmp_290_fu_11478_p4 = {{state_V_27_fu_11344_p2[79:72]}};

assign tmp_291_fu_11493_p4 = {{state_V_27_fu_11344_p2[87:80]}};

assign tmp_292_fu_11508_p4 = {{state_V_27_fu_11344_p2[95:88]}};

assign tmp_293_fu_11523_p4 = {{state_V_27_fu_11344_p2[103:96]}};

assign tmp_294_fu_11538_p4 = {{state_V_27_fu_11344_p2[111:104]}};

assign tmp_295_fu_11553_p4 = {{state_V_27_fu_11344_p2[119:112]}};

assign tmp_296_fu_11568_p4 = {{state_V_27_fu_11344_p2[127:120]}};

assign tmp_29_fu_4306_p4 = {{cipher_0_p16box_q132[15:8]}};

assign tmp_30_fu_4320_p4 = {{cipher_0_p16box_q131[15:8]}};

assign tmp_31_fu_4334_p4 = {{cipher_0_p16box_q130[15:8]}};

assign tmp_32_fu_4348_p4 = {{cipher_0_p16box_q129[15:8]}};

assign tmp_33_fu_4362_p4 = {{cipher_0_p16box_q128[15:8]}};

assign tmp_34_fu_4678_p4 = {{state_V_20_fu_4664_p2[15:8]}};

assign tmp_35_fu_4693_p4 = {{state_V_20_fu_4664_p2[23:16]}};

assign tmp_36_fu_4708_p4 = {{state_V_20_fu_4664_p2[31:24]}};

assign tmp_37_fu_4723_p4 = {{state_V_20_fu_4664_p2[39:32]}};

assign tmp_38_fu_4738_p4 = {{state_V_20_fu_4664_p2[47:40]}};

assign tmp_39_fu_4753_p4 = {{state_V_20_fu_4664_p2[55:48]}};

assign tmp_40_fu_4768_p4 = {{state_V_20_fu_4664_p2[63:56]}};

assign tmp_41_fu_4783_p4 = {{state_V_20_fu_4664_p2[71:64]}};

assign tmp_42_fu_4798_p4 = {{state_V_20_fu_4664_p2[79:72]}};

assign tmp_43_fu_4813_p4 = {{state_V_20_fu_4664_p2[87:80]}};

assign tmp_44_fu_4828_p4 = {{state_V_20_fu_4664_p2[95:88]}};

assign tmp_45_fu_4843_p4 = {{state_V_20_fu_4664_p2[103:96]}};

assign tmp_46_fu_4858_p4 = {{state_V_20_fu_4664_p2[111:104]}};

assign tmp_47_fu_4873_p4 = {{state_V_20_fu_4664_p2[119:112]}};

assign tmp_48_fu_4888_p4 = {{state_V_20_fu_4664_p2[127:120]}};

assign tmp_49_fu_4987_p4 = {{cipher_0_p16box_q127[15:8]}};

assign tmp_4_fu_3858_p4 = {{ret_V_fu_3828_p2[23:16]}};

assign tmp_50_fu_5001_p4 = {{cipher_0_p16box_q126[15:8]}};

assign tmp_51_fu_5015_p4 = {{cipher_0_p16box_q125[15:8]}};

assign tmp_52_fu_5029_p4 = {{cipher_0_p16box_q124[15:8]}};

assign tmp_53_fu_5043_p4 = {{cipher_0_p16box_q123[15:8]}};

assign tmp_54_fu_5057_p4 = {{cipher_0_p16box_q122[15:8]}};

assign tmp_55_fu_5071_p4 = {{cipher_0_p16box_q121[15:8]}};

assign tmp_56_fu_5085_p4 = {{cipher_0_p16box_q120[15:8]}};

assign tmp_57_fu_5099_p4 = {{cipher_0_p16box_q119[15:8]}};

assign tmp_58_fu_5113_p4 = {{cipher_0_p16box_q118[15:8]}};

assign tmp_59_fu_5127_p4 = {{cipher_0_p16box_q117[15:8]}};

assign tmp_5_fu_3873_p4 = {{ret_V_fu_3828_p2[31:24]}};

assign tmp_60_fu_5141_p4 = {{cipher_0_p16box_q116[15:8]}};

assign tmp_61_fu_5155_p4 = {{cipher_0_p16box_q115[15:8]}};

assign tmp_62_fu_5169_p4 = {{cipher_0_p16box_q114[15:8]}};

assign tmp_63_fu_5183_p4 = {{cipher_0_p16box_q113[15:8]}};

assign tmp_64_fu_5197_p4 = {{cipher_0_p16box_q112[15:8]}};

assign tmp_65_fu_5513_p4 = {{state_V_21_fu_5499_p2[15:8]}};

assign tmp_66_fu_5528_p4 = {{state_V_21_fu_5499_p2[23:16]}};

assign tmp_67_fu_5543_p4 = {{state_V_21_fu_5499_p2[31:24]}};

assign tmp_68_fu_5558_p4 = {{state_V_21_fu_5499_p2[39:32]}};

assign tmp_69_fu_5573_p4 = {{state_V_21_fu_5499_p2[47:40]}};

assign tmp_6_fu_3888_p4 = {{ret_V_fu_3828_p2[39:32]}};

assign tmp_70_fu_5588_p4 = {{state_V_21_fu_5499_p2[55:48]}};

assign tmp_71_fu_5603_p4 = {{state_V_21_fu_5499_p2[63:56]}};

assign tmp_72_fu_5618_p4 = {{state_V_21_fu_5499_p2[71:64]}};

assign tmp_73_fu_5633_p4 = {{state_V_21_fu_5499_p2[79:72]}};

assign tmp_74_fu_5648_p4 = {{state_V_21_fu_5499_p2[87:80]}};

assign tmp_75_fu_5663_p4 = {{state_V_21_fu_5499_p2[95:88]}};

assign tmp_76_fu_5678_p4 = {{state_V_21_fu_5499_p2[103:96]}};

assign tmp_77_fu_5693_p4 = {{state_V_21_fu_5499_p2[111:104]}};

assign tmp_78_fu_5708_p4 = {{state_V_21_fu_5499_p2[119:112]}};

assign tmp_79_fu_5723_p4 = {{state_V_21_fu_5499_p2[127:120]}};

assign tmp_7_fu_3903_p4 = {{ret_V_fu_3828_p2[47:40]}};

assign tmp_80_fu_5822_p4 = {{cipher_0_p16box_q111[15:8]}};

assign tmp_81_fu_5836_p4 = {{cipher_0_p16box_q110[15:8]}};

assign tmp_82_fu_5850_p4 = {{cipher_0_p16box_q109[15:8]}};

assign tmp_83_fu_5864_p4 = {{cipher_0_p16box_q108[15:8]}};

assign tmp_84_fu_5878_p4 = {{cipher_0_p16box_q107[15:8]}};

assign tmp_85_fu_5892_p4 = {{cipher_0_p16box_q106[15:8]}};

assign tmp_86_fu_5906_p4 = {{cipher_0_p16box_q105[15:8]}};

assign tmp_87_fu_5920_p4 = {{cipher_0_p16box_q104[15:8]}};

assign tmp_88_fu_5934_p4 = {{cipher_0_p16box_q103[15:8]}};

assign tmp_89_fu_5948_p4 = {{cipher_0_p16box_q102[15:8]}};

assign tmp_8_fu_3918_p4 = {{ret_V_fu_3828_p2[55:48]}};

assign tmp_90_fu_5962_p4 = {{cipher_0_p16box_q101[15:8]}};

assign tmp_91_fu_5976_p4 = {{cipher_0_p16box_q100[15:8]}};

assign tmp_92_fu_5990_p4 = {{cipher_0_p16box_q99[15:8]}};

assign tmp_93_fu_6004_p4 = {{cipher_0_p16box_q98[15:8]}};

assign tmp_94_fu_6018_p4 = {{cipher_0_p16box_q97[15:8]}};

assign tmp_95_fu_6032_p4 = {{cipher_0_p16box_q96[15:8]}};

assign tmp_96_fu_6348_p4 = {{state_V_22_fu_6334_p2[15:8]}};

assign tmp_97_fu_6363_p4 = {{state_V_22_fu_6334_p2[23:16]}};

assign tmp_98_fu_6378_p4 = {{state_V_22_fu_6334_p2[31:24]}};

assign tmp_99_fu_6393_p4 = {{state_V_22_fu_6334_p2[39:32]}};

assign tmp_9_fu_3933_p4 = {{ret_V_fu_3828_p2[63:56]}};

assign tmp_s_fu_3843_p4 = {{ret_V_fu_3828_p2[15:8]}};

assign trunc_ln674_100_fu_9214_p1 = cipher_0_p16box_q43[7:0];

assign trunc_ln674_101_fu_9228_p1 = cipher_0_p16box_q42[7:0];

assign trunc_ln674_102_fu_9242_p1 = cipher_0_p16box_q41[7:0];

assign trunc_ln674_103_fu_9256_p1 = cipher_0_p16box_q40[7:0];

assign trunc_ln674_104_fu_9270_p1 = cipher_0_p16box_q39[7:0];

assign trunc_ln674_105_fu_9284_p1 = cipher_0_p16box_q38[7:0];

assign trunc_ln674_106_fu_9298_p1 = cipher_0_p16box_q37[7:0];

assign trunc_ln674_107_fu_9312_p1 = cipher_0_p16box_q36[7:0];

assign trunc_ln674_108_fu_9326_p1 = cipher_0_p16box_q35[7:0];

assign trunc_ln674_109_fu_9340_p1 = cipher_0_p16box_q34[7:0];

assign trunc_ln674_10_fu_4288_p1 = cipher_0_p16box_q133[7:0];

assign trunc_ln674_110_fu_9354_p1 = cipher_0_p16box_q33[7:0];

assign trunc_ln674_111_fu_9368_p1 = cipher_0_p16box_q32[7:0];

assign trunc_ln674_112_fu_9993_p1 = cipher_0_p16box_q31[7:0];

assign trunc_ln674_113_fu_10007_p1 = cipher_0_p16box_q30[7:0];

assign trunc_ln674_114_fu_10021_p1 = cipher_0_p16box_q29[7:0];

assign trunc_ln674_115_fu_10035_p1 = cipher_0_p16box_q28[7:0];

assign trunc_ln674_116_fu_10049_p1 = cipher_0_p16box_q27[7:0];

assign trunc_ln674_117_fu_10063_p1 = cipher_0_p16box_q26[7:0];

assign trunc_ln674_118_fu_10077_p1 = cipher_0_p16box_q25[7:0];

assign trunc_ln674_119_fu_10091_p1 = cipher_0_p16box_q24[7:0];

assign trunc_ln674_11_fu_4302_p1 = cipher_0_p16box_q132[7:0];

assign trunc_ln674_120_fu_10105_p1 = cipher_0_p16box_q23[7:0];

assign trunc_ln674_121_fu_10119_p1 = cipher_0_p16box_q22[7:0];

assign trunc_ln674_122_fu_10133_p1 = cipher_0_p16box_q21[7:0];

assign trunc_ln674_123_fu_10147_p1 = cipher_0_p16box_q20[7:0];

assign trunc_ln674_124_fu_10161_p1 = cipher_0_p16box_q19[7:0];

assign trunc_ln674_125_fu_10175_p1 = cipher_0_p16box_q18[7:0];

assign trunc_ln674_126_fu_10189_p1 = cipher_0_p16box_q17[7:0];

assign trunc_ln674_127_fu_10203_p1 = cipher_0_p16box_q16[7:0];

assign trunc_ln674_128_fu_10828_p1 = cipher_0_p16box_q15[7:0];

assign trunc_ln674_129_fu_10842_p1 = cipher_0_p16box_q14[7:0];

assign trunc_ln674_12_fu_4316_p1 = cipher_0_p16box_q131[7:0];

assign trunc_ln674_130_fu_10856_p1 = cipher_0_p16box_q13[7:0];

assign trunc_ln674_131_fu_10870_p1 = cipher_0_p16box_q12[7:0];

assign trunc_ln674_132_fu_10884_p1 = cipher_0_p16box_q11[7:0];

assign trunc_ln674_133_fu_10898_p1 = cipher_0_p16box_q10[7:0];

assign trunc_ln674_134_fu_10912_p1 = cipher_0_p16box_q9[7:0];

assign trunc_ln674_135_fu_10926_p1 = cipher_0_p16box_q8[7:0];

assign trunc_ln674_136_fu_10940_p1 = cipher_0_p16box_q7[7:0];

assign trunc_ln674_137_fu_10954_p1 = cipher_0_p16box_q6[7:0];

assign trunc_ln674_138_fu_10968_p1 = cipher_0_p16box_q5[7:0];

assign trunc_ln674_139_fu_10982_p1 = cipher_0_p16box_q4[7:0];

assign trunc_ln674_13_fu_4330_p1 = cipher_0_p16box_q130[7:0];

assign trunc_ln674_140_fu_10996_p1 = cipher_0_p16box_q3[7:0];

assign trunc_ln674_141_fu_11010_p1 = cipher_0_p16box_q2[7:0];

assign trunc_ln674_142_fu_11024_p1 = cipher_0_p16box_q1[7:0];

assign trunc_ln674_143_fu_11038_p1 = cipher_0_p16box_q0[7:0];

assign trunc_ln674_14_fu_4344_p1 = cipher_0_p16box_q129[7:0];

assign trunc_ln674_15_fu_4358_p1 = cipher_0_p16box_q128[7:0];

assign trunc_ln674_16_fu_4983_p1 = cipher_0_p16box_q127[7:0];

assign trunc_ln674_17_fu_4997_p1 = cipher_0_p16box_q126[7:0];

assign trunc_ln674_18_fu_5011_p1 = cipher_0_p16box_q125[7:0];

assign trunc_ln674_19_fu_5025_p1 = cipher_0_p16box_q124[7:0];

assign trunc_ln674_1_fu_4162_p1 = cipher_0_p16box_q142[7:0];

assign trunc_ln674_20_fu_5039_p1 = cipher_0_p16box_q123[7:0];

assign trunc_ln674_21_fu_5053_p1 = cipher_0_p16box_q122[7:0];

assign trunc_ln674_22_fu_5067_p1 = cipher_0_p16box_q121[7:0];

assign trunc_ln674_23_fu_5081_p1 = cipher_0_p16box_q120[7:0];

assign trunc_ln674_24_fu_5095_p1 = cipher_0_p16box_q119[7:0];

assign trunc_ln674_25_fu_5109_p1 = cipher_0_p16box_q118[7:0];

assign trunc_ln674_26_fu_5123_p1 = cipher_0_p16box_q117[7:0];

assign trunc_ln674_27_fu_5137_p1 = cipher_0_p16box_q116[7:0];

assign trunc_ln674_28_fu_5151_p1 = cipher_0_p16box_q115[7:0];

assign trunc_ln674_29_fu_5165_p1 = cipher_0_p16box_q114[7:0];

assign trunc_ln674_2_fu_4176_p1 = cipher_0_p16box_q141[7:0];

assign trunc_ln674_30_fu_5179_p1 = cipher_0_p16box_q113[7:0];

assign trunc_ln674_31_fu_5193_p1 = cipher_0_p16box_q112[7:0];

assign trunc_ln674_32_fu_5818_p1 = cipher_0_p16box_q111[7:0];

assign trunc_ln674_33_fu_5832_p1 = cipher_0_p16box_q110[7:0];

assign trunc_ln674_34_fu_5846_p1 = cipher_0_p16box_q109[7:0];

assign trunc_ln674_35_fu_5860_p1 = cipher_0_p16box_q108[7:0];

assign trunc_ln674_36_fu_5874_p1 = cipher_0_p16box_q107[7:0];

assign trunc_ln674_37_fu_5888_p1 = cipher_0_p16box_q106[7:0];

assign trunc_ln674_38_fu_5902_p1 = cipher_0_p16box_q105[7:0];

assign trunc_ln674_39_fu_5916_p1 = cipher_0_p16box_q104[7:0];

assign trunc_ln674_3_fu_4190_p1 = cipher_0_p16box_q140[7:0];

assign trunc_ln674_40_fu_5930_p1 = cipher_0_p16box_q103[7:0];

assign trunc_ln674_41_fu_5944_p1 = cipher_0_p16box_q102[7:0];

assign trunc_ln674_42_fu_5958_p1 = cipher_0_p16box_q101[7:0];

assign trunc_ln674_43_fu_5972_p1 = cipher_0_p16box_q100[7:0];

assign trunc_ln674_44_fu_5986_p1 = cipher_0_p16box_q99[7:0];

assign trunc_ln674_45_fu_6000_p1 = cipher_0_p16box_q98[7:0];

assign trunc_ln674_46_fu_6014_p1 = cipher_0_p16box_q97[7:0];

assign trunc_ln674_47_fu_6028_p1 = cipher_0_p16box_q96[7:0];

assign trunc_ln674_48_fu_6653_p1 = cipher_0_p16box_q95[7:0];

assign trunc_ln674_49_fu_6667_p1 = cipher_0_p16box_q94[7:0];

assign trunc_ln674_4_fu_4204_p1 = cipher_0_p16box_q139[7:0];

assign trunc_ln674_50_fu_6681_p1 = cipher_0_p16box_q93[7:0];

assign trunc_ln674_51_fu_6695_p1 = cipher_0_p16box_q92[7:0];

assign trunc_ln674_52_fu_6709_p1 = cipher_0_p16box_q91[7:0];

assign trunc_ln674_53_fu_6723_p1 = cipher_0_p16box_q90[7:0];

assign trunc_ln674_54_fu_6737_p1 = cipher_0_p16box_q89[7:0];

assign trunc_ln674_55_fu_6751_p1 = cipher_0_p16box_q88[7:0];

assign trunc_ln674_56_fu_6765_p1 = cipher_0_p16box_q87[7:0];

assign trunc_ln674_57_fu_6779_p1 = cipher_0_p16box_q86[7:0];

assign trunc_ln674_58_fu_6793_p1 = cipher_0_p16box_q85[7:0];

assign trunc_ln674_59_fu_6807_p1 = cipher_0_p16box_q84[7:0];

assign trunc_ln674_5_fu_4218_p1 = cipher_0_p16box_q138[7:0];

assign trunc_ln674_60_fu_6821_p1 = cipher_0_p16box_q83[7:0];

assign trunc_ln674_61_fu_6835_p1 = cipher_0_p16box_q82[7:0];

assign trunc_ln674_62_fu_6849_p1 = cipher_0_p16box_q81[7:0];

assign trunc_ln674_63_fu_6863_p1 = cipher_0_p16box_q80[7:0];

assign trunc_ln674_64_fu_7488_p1 = cipher_0_p16box_q79[7:0];

assign trunc_ln674_65_fu_7502_p1 = cipher_0_p16box_q78[7:0];

assign trunc_ln674_66_fu_7516_p1 = cipher_0_p16box_q77[7:0];

assign trunc_ln674_67_fu_7530_p1 = cipher_0_p16box_q76[7:0];

assign trunc_ln674_68_fu_7544_p1 = cipher_0_p16box_q75[7:0];

assign trunc_ln674_69_fu_7558_p1 = cipher_0_p16box_q74[7:0];

assign trunc_ln674_6_fu_4232_p1 = cipher_0_p16box_q137[7:0];

assign trunc_ln674_70_fu_7572_p1 = cipher_0_p16box_q73[7:0];

assign trunc_ln674_71_fu_7586_p1 = cipher_0_p16box_q72[7:0];

assign trunc_ln674_72_fu_7600_p1 = cipher_0_p16box_q71[7:0];

assign trunc_ln674_73_fu_7614_p1 = cipher_0_p16box_q70[7:0];

assign trunc_ln674_74_fu_7628_p1 = cipher_0_p16box_q69[7:0];

assign trunc_ln674_75_fu_7642_p1 = cipher_0_p16box_q68[7:0];

assign trunc_ln674_76_fu_7656_p1 = cipher_0_p16box_q67[7:0];

assign trunc_ln674_77_fu_7670_p1 = cipher_0_p16box_q66[7:0];

assign trunc_ln674_78_fu_7684_p1 = cipher_0_p16box_q65[7:0];

assign trunc_ln674_79_fu_7698_p1 = cipher_0_p16box_q64[7:0];

assign trunc_ln674_7_fu_4246_p1 = cipher_0_p16box_q136[7:0];

assign trunc_ln674_80_fu_8323_p1 = cipher_0_p16box_q63[7:0];

assign trunc_ln674_81_fu_8337_p1 = cipher_0_p16box_q62[7:0];

assign trunc_ln674_82_fu_8351_p1 = cipher_0_p16box_q61[7:0];

assign trunc_ln674_83_fu_8365_p1 = cipher_0_p16box_q60[7:0];

assign trunc_ln674_84_fu_8379_p1 = cipher_0_p16box_q59[7:0];

assign trunc_ln674_85_fu_8393_p1 = cipher_0_p16box_q58[7:0];

assign trunc_ln674_86_fu_8407_p1 = cipher_0_p16box_q57[7:0];

assign trunc_ln674_87_fu_8421_p1 = cipher_0_p16box_q56[7:0];

assign trunc_ln674_88_fu_8435_p1 = cipher_0_p16box_q55[7:0];

assign trunc_ln674_89_fu_8449_p1 = cipher_0_p16box_q54[7:0];

assign trunc_ln674_8_fu_4260_p1 = cipher_0_p16box_q135[7:0];

assign trunc_ln674_90_fu_8463_p1 = cipher_0_p16box_q53[7:0];

assign trunc_ln674_91_fu_8477_p1 = cipher_0_p16box_q52[7:0];

assign trunc_ln674_92_fu_8491_p1 = cipher_0_p16box_q51[7:0];

assign trunc_ln674_93_fu_8505_p1 = cipher_0_p16box_q50[7:0];

assign trunc_ln674_94_fu_8519_p1 = cipher_0_p16box_q49[7:0];

assign trunc_ln674_95_fu_8533_p1 = cipher_0_p16box_q48[7:0];

assign trunc_ln674_96_fu_9158_p1 = cipher_0_p16box_q47[7:0];

assign trunc_ln674_97_fu_9172_p1 = cipher_0_p16box_q46[7:0];

assign trunc_ln674_98_fu_9186_p1 = cipher_0_p16box_q45[7:0];

assign trunc_ln674_99_fu_9200_p1 = cipher_0_p16box_q44[7:0];

assign trunc_ln674_9_fu_4274_p1 = cipher_0_p16box_q134[7:0];

assign trunc_ln674_fu_4148_p1 = cipher_0_p16box_q143[7:0];

assign trunc_ln708_1_fu_4669_p1 = state_V_20_fu_4664_p2[7:0];

assign trunc_ln708_2_fu_5504_p1 = state_V_21_fu_5499_p2[7:0];

assign trunc_ln708_3_fu_6339_p1 = state_V_22_fu_6334_p2[7:0];

assign trunc_ln708_4_fu_7174_p1 = state_V_23_fu_7169_p2[7:0];

assign trunc_ln708_5_fu_8009_p1 = state_V_24_fu_8004_p2[7:0];

assign trunc_ln708_6_fu_8844_p1 = state_V_25_fu_8839_p2[7:0];

assign trunc_ln708_7_fu_9679_p1 = state_V_fu_9674_p2[7:0];

assign trunc_ln708_8_fu_10514_p1 = state_V_26_fu_10509_p2[7:0];

assign trunc_ln708_9_fu_11349_p1 = state_V_27_fu_11344_p2[7:0];

assign trunc_ln708_fu_3834_p1 = ret_V_fu_3828_p2[7:0];

assign xor_ln1545_100_fu_6042_p2 = (tmp_V_34_reg_12326 ^ tmp_3_V_12_reg_12356);

assign xor_ln1545_101_fu_6052_p2 = (xor_ln1545_102_fu_6046_p2 ^ xor_ln1545_100_fu_6042_p2);

assign xor_ln1545_102_fu_6046_p2 = (trunc_ln674_32_fu_5818_p1 ^ tmp_81_fu_5836_p4);

assign xor_ln1545_103_fu_6058_p2 = (tmp_V_32_reg_12266 ^ tmp_3_V_12_reg_12356);

assign xor_ln1545_104_fu_6068_p2 = (xor_ln1545_105_fu_6062_p2 ^ xor_ln1545_103_fu_6058_p2);

assign xor_ln1545_105_fu_6062_p2 = (trunc_ln674_33_fu_5832_p1 ^ tmp_82_fu_5850_p4);

assign xor_ln1545_106_fu_6074_p2 = (tmp_V_33_reg_12296 ^ tmp_V_32_reg_12266);

assign xor_ln1545_107_fu_6084_p2 = (xor_ln1545_108_fu_6078_p2 ^ xor_ln1545_106_fu_6074_p2);

assign xor_ln1545_108_fu_6078_p2 = (trunc_ln674_34_fu_5846_p1 ^ tmp_83_fu_5864_p4);

assign xor_ln1545_109_fu_6090_p2 = (tmp_V_34_reg_12326 ^ tmp_V_33_reg_12296);

assign xor_ln1545_10_fu_4404_p2 = (tmp_V_reg_11754 ^ tmp_V_1_reg_11784);

assign xor_ln1545_110_fu_6100_p2 = (xor_ln1545_111_fu_6094_p2 ^ xor_ln1545_109_fu_6090_p2);

assign xor_ln1545_111_fu_6094_p2 = (trunc_ln674_35_fu_5860_p1 ^ tmp_80_fu_5822_p4);

assign xor_ln1545_112_fu_6106_p2 = (tmp_V_39_reg_12284 ^ tmp_V_38_reg_12350);

assign xor_ln1545_113_fu_6116_p2 = (xor_ln1545_114_fu_6110_p2 ^ xor_ln1545_112_fu_6106_p2);

assign xor_ln1545_114_fu_6110_p2 = (trunc_ln674_36_fu_5874_p1 ^ tmp_85_fu_5892_p4);

assign xor_ln1545_115_fu_6122_p2 = (tmp_V_39_reg_12284 ^ tmp_V_36_reg_12290);

assign xor_ln1545_116_fu_6132_p2 = (xor_ln1545_117_fu_6126_p2 ^ xor_ln1545_115_fu_6122_p2);

assign xor_ln1545_117_fu_6126_p2 = (trunc_ln674_37_fu_5888_p1 ^ tmp_86_fu_5906_p4);

assign xor_ln1545_118_fu_6138_p2 = (tmp_V_37_reg_12320 ^ tmp_V_36_reg_12290);

assign xor_ln1545_119_fu_6148_p2 = (xor_ln1545_120_fu_6142_p2 ^ xor_ln1545_118_fu_6138_p2);

assign xor_ln1545_11_fu_4414_p2 = (xor_ln1545_12_fu_4408_p2 ^ xor_ln1545_10_fu_4404_p2);

assign xor_ln1545_120_fu_6142_p2 = (trunc_ln674_38_fu_5902_p1 ^ tmp_87_fu_5920_p4);

assign xor_ln1545_121_fu_6154_p2 = (tmp_V_38_reg_12350 ^ tmp_V_37_reg_12320);

assign xor_ln1545_122_fu_6164_p2 = (xor_ln1545_123_fu_6158_p2 ^ xor_ln1545_121_fu_6154_p2);

assign xor_ln1545_123_fu_6158_p2 = (trunc_ln674_39_fu_5916_p1 ^ tmp_84_fu_5878_p4);

assign xor_ln1545_124_fu_6170_p2 = (tmp_V_43_reg_12308 ^ tmp_2_1_V_12_reg_12278);

assign xor_ln1545_125_fu_6180_p2 = (xor_ln1545_126_fu_6174_p2 ^ xor_ln1545_124_fu_6170_p2);

assign xor_ln1545_126_fu_6174_p2 = (trunc_ln674_40_fu_5930_p1 ^ tmp_89_fu_5948_p4);

assign xor_ln1545_127_fu_6186_p2 = (tmp_V_43_reg_12308 ^ tmp_V_40_reg_12314);

assign xor_ln1545_128_fu_6196_p2 = (xor_ln1545_129_fu_6190_p2 ^ xor_ln1545_127_fu_6186_p2);

assign xor_ln1545_129_fu_6190_p2 = (trunc_ln674_41_fu_5944_p1 ^ tmp_90_fu_5962_p4);

assign xor_ln1545_12_fu_4408_p2 = (trunc_ln674_2_fu_4176_p1 ^ tmp_21_fu_4194_p4);

assign xor_ln1545_130_fu_6202_p2 = (tmp_V_41_reg_12344 ^ tmp_V_40_reg_12314);

assign xor_ln1545_131_fu_6212_p2 = (xor_ln1545_132_fu_6206_p2 ^ xor_ln1545_130_fu_6202_p2);

assign xor_ln1545_132_fu_6206_p2 = (trunc_ln674_42_fu_5958_p1 ^ tmp_91_fu_5976_p4);

assign xor_ln1545_133_fu_6218_p2 = (tmp_V_41_reg_12344 ^ tmp_2_1_V_12_reg_12278);

assign xor_ln1545_134_fu_6228_p2 = (xor_ln1545_135_fu_6222_p2 ^ xor_ln1545_133_fu_6218_p2);

assign xor_ln1545_135_fu_6222_p2 = (trunc_ln674_43_fu_5972_p1 ^ tmp_88_fu_5934_p4);

assign xor_ln1545_136_fu_6234_p2 = (tmp_V_47_reg_12332 ^ tmp_2_2_V_12_reg_12302);

assign xor_ln1545_137_fu_6244_p2 = (xor_ln1545_138_fu_6238_p2 ^ xor_ln1545_136_fu_6234_p2);

assign xor_ln1545_138_fu_6238_p2 = (trunc_ln674_44_fu_5986_p1 ^ tmp_93_fu_6004_p4);

assign xor_ln1545_139_fu_6250_p2 = (tmp_V_47_reg_12332 ^ tmp_V_44_reg_12338);

assign xor_ln1545_13_fu_4420_p2 = (tmp_V_2_reg_11814 ^ tmp_V_1_reg_11784);

assign xor_ln1545_140_fu_6260_p2 = (xor_ln1545_141_fu_6254_p2 ^ xor_ln1545_139_fu_6250_p2);

assign xor_ln1545_141_fu_6254_p2 = (trunc_ln674_45_fu_6000_p1 ^ tmp_94_fu_6018_p4);

assign xor_ln1545_142_fu_6266_p2 = (tmp_V_44_reg_12338 ^ tmp_1_V_12_reg_12272);

assign xor_ln1545_143_fu_6276_p2 = (xor_ln1545_144_fu_6270_p2 ^ xor_ln1545_142_fu_6266_p2);

assign xor_ln1545_144_fu_6270_p2 = (trunc_ln674_46_fu_6014_p1 ^ tmp_95_fu_6032_p4);

assign xor_ln1545_145_fu_6282_p2 = (tmp_2_2_V_12_reg_12302 ^ tmp_1_V_12_reg_12272);

assign xor_ln1545_146_fu_6292_p2 = (xor_ln1545_147_fu_6286_p2 ^ xor_ln1545_145_fu_6282_p2);

assign xor_ln1545_147_fu_6286_p2 = (trunc_ln674_47_fu_6028_p1 ^ tmp_92_fu_5990_p4);

assign xor_ln1545_148_fu_6877_p2 = (tmp_V_50_reg_12582 ^ tmp_3_V_13_reg_12612);

assign xor_ln1545_149_fu_6887_p2 = (xor_ln1545_150_fu_6881_p2 ^ xor_ln1545_148_fu_6877_p2);

assign xor_ln1545_14_fu_4430_p2 = (xor_ln1545_15_fu_4424_p2 ^ xor_ln1545_13_fu_4420_p2);

assign xor_ln1545_150_fu_6881_p2 = (trunc_ln674_48_fu_6653_p1 ^ tmp_112_fu_6671_p4);

assign xor_ln1545_151_fu_6893_p2 = (tmp_V_48_reg_12522 ^ tmp_3_V_13_reg_12612);

assign xor_ln1545_152_fu_6903_p2 = (xor_ln1545_153_fu_6897_p2 ^ xor_ln1545_151_fu_6893_p2);

assign xor_ln1545_153_fu_6897_p2 = (trunc_ln674_49_fu_6667_p1 ^ tmp_113_fu_6685_p4);

assign xor_ln1545_154_fu_6909_p2 = (tmp_V_49_reg_12552 ^ tmp_V_48_reg_12522);

assign xor_ln1545_155_fu_6919_p2 = (xor_ln1545_156_fu_6913_p2 ^ xor_ln1545_154_fu_6909_p2);

assign xor_ln1545_156_fu_6913_p2 = (trunc_ln674_50_fu_6681_p1 ^ tmp_114_fu_6699_p4);

assign xor_ln1545_157_fu_6925_p2 = (tmp_V_50_reg_12582 ^ tmp_V_49_reg_12552);

assign xor_ln1545_158_fu_6935_p2 = (xor_ln1545_159_fu_6929_p2 ^ xor_ln1545_157_fu_6925_p2);

assign xor_ln1545_159_fu_6929_p2 = (trunc_ln674_51_fu_6695_p1 ^ tmp_111_fu_6657_p4);

assign xor_ln1545_15_fu_4424_p2 = (trunc_ln674_3_fu_4190_p1 ^ tmp_18_fu_4152_p4);

assign xor_ln1545_160_fu_6941_p2 = (tmp_V_55_reg_12540 ^ tmp_V_54_reg_12606);

assign xor_ln1545_161_fu_6951_p2 = (xor_ln1545_162_fu_6945_p2 ^ xor_ln1545_160_fu_6941_p2);

assign xor_ln1545_162_fu_6945_p2 = (trunc_ln674_52_fu_6709_p1 ^ tmp_116_fu_6727_p4);

assign xor_ln1545_163_fu_6957_p2 = (tmp_V_55_reg_12540 ^ tmp_V_52_reg_12546);

assign xor_ln1545_164_fu_6967_p2 = (xor_ln1545_165_fu_6961_p2 ^ xor_ln1545_163_fu_6957_p2);

assign xor_ln1545_165_fu_6961_p2 = (trunc_ln674_53_fu_6723_p1 ^ tmp_117_fu_6741_p4);

assign xor_ln1545_166_fu_6973_p2 = (tmp_V_53_reg_12576 ^ tmp_V_52_reg_12546);

assign xor_ln1545_167_fu_6983_p2 = (xor_ln1545_168_fu_6977_p2 ^ xor_ln1545_166_fu_6973_p2);

assign xor_ln1545_168_fu_6977_p2 = (trunc_ln674_54_fu_6737_p1 ^ tmp_118_fu_6755_p4);

assign xor_ln1545_169_fu_6989_p2 = (tmp_V_54_reg_12606 ^ tmp_V_53_reg_12576);

assign xor_ln1545_16_fu_4436_p2 = (tmp_V_7_reg_11772 ^ tmp_V_6_reg_11838);

assign xor_ln1545_170_fu_6999_p2 = (xor_ln1545_171_fu_6993_p2 ^ xor_ln1545_169_fu_6989_p2);

assign xor_ln1545_171_fu_6993_p2 = (trunc_ln674_55_fu_6751_p1 ^ tmp_115_fu_6713_p4);

assign xor_ln1545_172_fu_7005_p2 = (tmp_V_59_reg_12564 ^ tmp_2_1_V_13_reg_12534);

assign xor_ln1545_173_fu_7015_p2 = (xor_ln1545_174_fu_7009_p2 ^ xor_ln1545_172_fu_7005_p2);

assign xor_ln1545_174_fu_7009_p2 = (trunc_ln674_56_fu_6765_p1 ^ tmp_120_fu_6783_p4);

assign xor_ln1545_175_fu_7021_p2 = (tmp_V_59_reg_12564 ^ tmp_V_56_reg_12570);

assign xor_ln1545_176_fu_7031_p2 = (xor_ln1545_177_fu_7025_p2 ^ xor_ln1545_175_fu_7021_p2);

assign xor_ln1545_177_fu_7025_p2 = (trunc_ln674_57_fu_6779_p1 ^ tmp_121_fu_6797_p4);

assign xor_ln1545_178_fu_7037_p2 = (tmp_V_57_reg_12600 ^ tmp_V_56_reg_12570);

assign xor_ln1545_179_fu_7047_p2 = (xor_ln1545_180_fu_7041_p2 ^ xor_ln1545_178_fu_7037_p2);

assign xor_ln1545_17_fu_4446_p2 = (xor_ln1545_18_fu_4440_p2 ^ xor_ln1545_16_fu_4436_p2);

assign xor_ln1545_180_fu_7041_p2 = (trunc_ln674_58_fu_6793_p1 ^ tmp_122_fu_6811_p4);

assign xor_ln1545_181_fu_7053_p2 = (tmp_V_57_reg_12600 ^ tmp_2_1_V_13_reg_12534);

assign xor_ln1545_182_fu_7063_p2 = (xor_ln1545_183_fu_7057_p2 ^ xor_ln1545_181_fu_7053_p2);

assign xor_ln1545_183_fu_7057_p2 = (trunc_ln674_59_fu_6807_p1 ^ tmp_119_fu_6769_p4);

assign xor_ln1545_184_fu_7069_p2 = (tmp_V_63_reg_12588 ^ tmp_2_2_V_13_reg_12558);

assign xor_ln1545_185_fu_7079_p2 = (xor_ln1545_186_fu_7073_p2 ^ xor_ln1545_184_fu_7069_p2);

assign xor_ln1545_186_fu_7073_p2 = (trunc_ln674_60_fu_6821_p1 ^ tmp_124_fu_6839_p4);

assign xor_ln1545_187_fu_7085_p2 = (tmp_V_63_reg_12588 ^ tmp_V_60_reg_12594);

assign xor_ln1545_188_fu_7095_p2 = (xor_ln1545_189_fu_7089_p2 ^ xor_ln1545_187_fu_7085_p2);

assign xor_ln1545_189_fu_7089_p2 = (trunc_ln674_61_fu_6835_p1 ^ tmp_125_fu_6853_p4);

assign xor_ln1545_18_fu_4440_p2 = (trunc_ln674_4_fu_4204_p1 ^ tmp_23_fu_4222_p4);

assign xor_ln1545_190_fu_7101_p2 = (tmp_V_60_reg_12594 ^ tmp_1_V_13_reg_12528);

assign xor_ln1545_191_fu_7111_p2 = (xor_ln1545_192_fu_7105_p2 ^ xor_ln1545_190_fu_7101_p2);

assign xor_ln1545_192_fu_7105_p2 = (trunc_ln674_62_fu_6849_p1 ^ tmp_126_fu_6867_p4);

assign xor_ln1545_193_fu_7117_p2 = (tmp_2_2_V_13_reg_12558 ^ tmp_1_V_13_reg_12528);

assign xor_ln1545_194_fu_7127_p2 = (xor_ln1545_195_fu_7121_p2 ^ xor_ln1545_193_fu_7117_p2);

assign xor_ln1545_195_fu_7121_p2 = (trunc_ln674_63_fu_6863_p1 ^ tmp_123_fu_6825_p4);

assign xor_ln1545_196_fu_7712_p2 = (tmp_V_66_reg_12838 ^ tmp_3_V_14_reg_12868);

assign xor_ln1545_197_fu_7722_p2 = (xor_ln1545_198_fu_7716_p2 ^ xor_ln1545_196_fu_7712_p2);

assign xor_ln1545_198_fu_7716_p2 = (trunc_ln674_64_fu_7488_p1 ^ tmp_143_fu_7506_p4);

assign xor_ln1545_199_fu_7728_p2 = (tmp_V_64_reg_12778 ^ tmp_3_V_14_reg_12868);

assign xor_ln1545_19_fu_4452_p2 = (tmp_V_7_reg_11772 ^ tmp_V_4_reg_11778);

assign xor_ln1545_200_fu_7738_p2 = (xor_ln1545_201_fu_7732_p2 ^ xor_ln1545_199_fu_7728_p2);

assign xor_ln1545_201_fu_7732_p2 = (trunc_ln674_65_fu_7502_p1 ^ tmp_144_fu_7520_p4);

assign xor_ln1545_202_fu_7744_p2 = (tmp_V_65_reg_12808 ^ tmp_V_64_reg_12778);

assign xor_ln1545_203_fu_7754_p2 = (xor_ln1545_204_fu_7748_p2 ^ xor_ln1545_202_fu_7744_p2);

assign xor_ln1545_204_fu_7748_p2 = (trunc_ln674_66_fu_7516_p1 ^ tmp_145_fu_7534_p4);

assign xor_ln1545_205_fu_7760_p2 = (tmp_V_66_reg_12838 ^ tmp_V_65_reg_12808);

assign xor_ln1545_206_fu_7770_p2 = (xor_ln1545_207_fu_7764_p2 ^ xor_ln1545_205_fu_7760_p2);

assign xor_ln1545_207_fu_7764_p2 = (trunc_ln674_67_fu_7530_p1 ^ tmp_142_fu_7492_p4);

assign xor_ln1545_208_fu_7776_p2 = (tmp_V_71_reg_12796 ^ tmp_V_70_reg_12862);

assign xor_ln1545_209_fu_7786_p2 = (xor_ln1545_210_fu_7780_p2 ^ xor_ln1545_208_fu_7776_p2);

assign xor_ln1545_20_fu_4462_p2 = (xor_ln1545_21_fu_4456_p2 ^ xor_ln1545_19_fu_4452_p2);

assign xor_ln1545_210_fu_7780_p2 = (trunc_ln674_68_fu_7544_p1 ^ tmp_147_fu_7562_p4);

assign xor_ln1545_211_fu_7792_p2 = (tmp_V_71_reg_12796 ^ tmp_V_68_reg_12802);

assign xor_ln1545_212_fu_7802_p2 = (xor_ln1545_213_fu_7796_p2 ^ xor_ln1545_211_fu_7792_p2);

assign xor_ln1545_213_fu_7796_p2 = (trunc_ln674_69_fu_7558_p1 ^ tmp_148_fu_7576_p4);

assign xor_ln1545_214_fu_7808_p2 = (tmp_V_69_reg_12832 ^ tmp_V_68_reg_12802);

assign xor_ln1545_215_fu_7818_p2 = (xor_ln1545_216_fu_7812_p2 ^ xor_ln1545_214_fu_7808_p2);

assign xor_ln1545_216_fu_7812_p2 = (trunc_ln674_70_fu_7572_p1 ^ tmp_149_fu_7590_p4);

assign xor_ln1545_217_fu_7824_p2 = (tmp_V_70_reg_12862 ^ tmp_V_69_reg_12832);

assign xor_ln1545_218_fu_7834_p2 = (xor_ln1545_219_fu_7828_p2 ^ xor_ln1545_217_fu_7824_p2);

assign xor_ln1545_219_fu_7828_p2 = (trunc_ln674_71_fu_7586_p1 ^ tmp_146_fu_7548_p4);

assign xor_ln1545_21_fu_4456_p2 = (trunc_ln674_5_fu_4218_p1 ^ tmp_24_fu_4236_p4);

assign xor_ln1545_220_fu_7840_p2 = (tmp_V_75_reg_12820 ^ tmp_2_1_V_14_reg_12790);

assign xor_ln1545_221_fu_7850_p2 = (xor_ln1545_222_fu_7844_p2 ^ xor_ln1545_220_fu_7840_p2);

assign xor_ln1545_222_fu_7844_p2 = (trunc_ln674_72_fu_7600_p1 ^ tmp_151_fu_7618_p4);

assign xor_ln1545_223_fu_7856_p2 = (tmp_V_75_reg_12820 ^ tmp_V_72_reg_12826);

assign xor_ln1545_224_fu_7866_p2 = (xor_ln1545_225_fu_7860_p2 ^ xor_ln1545_223_fu_7856_p2);

assign xor_ln1545_225_fu_7860_p2 = (trunc_ln674_73_fu_7614_p1 ^ tmp_152_fu_7632_p4);

assign xor_ln1545_226_fu_7872_p2 = (tmp_V_73_reg_12856 ^ tmp_V_72_reg_12826);

assign xor_ln1545_227_fu_7882_p2 = (xor_ln1545_228_fu_7876_p2 ^ xor_ln1545_226_fu_7872_p2);

assign xor_ln1545_228_fu_7876_p2 = (trunc_ln674_74_fu_7628_p1 ^ tmp_153_fu_7646_p4);

assign xor_ln1545_229_fu_7888_p2 = (tmp_V_73_reg_12856 ^ tmp_2_1_V_14_reg_12790);

assign xor_ln1545_22_fu_4468_p2 = (tmp_V_5_reg_11808 ^ tmp_V_4_reg_11778);

assign xor_ln1545_230_fu_7898_p2 = (xor_ln1545_231_fu_7892_p2 ^ xor_ln1545_229_fu_7888_p2);

assign xor_ln1545_231_fu_7892_p2 = (trunc_ln674_75_fu_7642_p1 ^ tmp_150_fu_7604_p4);

assign xor_ln1545_232_fu_7904_p2 = (tmp_V_79_reg_12844 ^ tmp_2_2_V_14_reg_12814);

assign xor_ln1545_233_fu_7914_p2 = (xor_ln1545_234_fu_7908_p2 ^ xor_ln1545_232_fu_7904_p2);

assign xor_ln1545_234_fu_7908_p2 = (trunc_ln674_76_fu_7656_p1 ^ tmp_155_fu_7674_p4);

assign xor_ln1545_235_fu_7920_p2 = (tmp_V_79_reg_12844 ^ tmp_V_76_reg_12850);

assign xor_ln1545_236_fu_7930_p2 = (xor_ln1545_237_fu_7924_p2 ^ xor_ln1545_235_fu_7920_p2);

assign xor_ln1545_237_fu_7924_p2 = (trunc_ln674_77_fu_7670_p1 ^ tmp_156_fu_7688_p4);

assign xor_ln1545_238_fu_7936_p2 = (tmp_V_76_reg_12850 ^ tmp_1_V_14_reg_12784);

assign xor_ln1545_239_fu_7946_p2 = (xor_ln1545_240_fu_7940_p2 ^ xor_ln1545_238_fu_7936_p2);

assign xor_ln1545_23_fu_4478_p2 = (xor_ln1545_24_fu_4472_p2 ^ xor_ln1545_22_fu_4468_p2);

assign xor_ln1545_240_fu_7940_p2 = (trunc_ln674_78_fu_7684_p1 ^ tmp_157_fu_7702_p4);

assign xor_ln1545_241_fu_7952_p2 = (tmp_2_2_V_14_reg_12814 ^ tmp_1_V_14_reg_12784);

assign xor_ln1545_242_fu_7962_p2 = (xor_ln1545_243_fu_7956_p2 ^ xor_ln1545_241_fu_7952_p2);

assign xor_ln1545_243_fu_7956_p2 = (trunc_ln674_79_fu_7698_p1 ^ tmp_154_fu_7660_p4);

assign xor_ln1545_244_fu_8547_p2 = (tmp_V_82_reg_13094 ^ tmp_3_V_15_reg_13124);

assign xor_ln1545_245_fu_8557_p2 = (xor_ln1545_246_fu_8551_p2 ^ xor_ln1545_244_fu_8547_p2);

assign xor_ln1545_246_fu_8551_p2 = (trunc_ln674_80_fu_8323_p1 ^ tmp_174_fu_8341_p4);

assign xor_ln1545_247_fu_8563_p2 = (tmp_V_80_reg_13034 ^ tmp_3_V_15_reg_13124);

assign xor_ln1545_248_fu_8573_p2 = (xor_ln1545_249_fu_8567_p2 ^ xor_ln1545_247_fu_8563_p2);

assign xor_ln1545_249_fu_8567_p2 = (trunc_ln674_81_fu_8337_p1 ^ tmp_175_fu_8355_p4);

assign xor_ln1545_24_fu_4472_p2 = (trunc_ln674_6_fu_4232_p1 ^ tmp_25_fu_4250_p4);

assign xor_ln1545_250_fu_8579_p2 = (tmp_V_81_reg_13064 ^ tmp_V_80_reg_13034);

assign xor_ln1545_251_fu_8589_p2 = (xor_ln1545_252_fu_8583_p2 ^ xor_ln1545_250_fu_8579_p2);

assign xor_ln1545_252_fu_8583_p2 = (trunc_ln674_82_fu_8351_p1 ^ tmp_176_fu_8369_p4);

assign xor_ln1545_253_fu_8595_p2 = (tmp_V_82_reg_13094 ^ tmp_V_81_reg_13064);

assign xor_ln1545_254_fu_8605_p2 = (xor_ln1545_255_fu_8599_p2 ^ xor_ln1545_253_fu_8595_p2);

assign xor_ln1545_255_fu_8599_p2 = (trunc_ln674_83_fu_8365_p1 ^ tmp_173_fu_8327_p4);

assign xor_ln1545_256_fu_8611_p2 = (tmp_V_87_reg_13052 ^ tmp_V_86_reg_13118);

assign xor_ln1545_257_fu_8621_p2 = (xor_ln1545_258_fu_8615_p2 ^ xor_ln1545_256_fu_8611_p2);

assign xor_ln1545_258_fu_8615_p2 = (trunc_ln674_84_fu_8379_p1 ^ tmp_178_fu_8397_p4);

assign xor_ln1545_259_fu_8627_p2 = (tmp_V_87_reg_13052 ^ tmp_V_84_reg_13058);

assign xor_ln1545_25_fu_4484_p2 = (tmp_V_6_reg_11838 ^ tmp_V_5_reg_11808);

assign xor_ln1545_260_fu_8637_p2 = (xor_ln1545_261_fu_8631_p2 ^ xor_ln1545_259_fu_8627_p2);

assign xor_ln1545_261_fu_8631_p2 = (trunc_ln674_85_fu_8393_p1 ^ tmp_179_fu_8411_p4);

assign xor_ln1545_262_fu_8643_p2 = (tmp_V_85_reg_13088 ^ tmp_V_84_reg_13058);

assign xor_ln1545_263_fu_8653_p2 = (xor_ln1545_264_fu_8647_p2 ^ xor_ln1545_262_fu_8643_p2);

assign xor_ln1545_264_fu_8647_p2 = (trunc_ln674_86_fu_8407_p1 ^ tmp_180_fu_8425_p4);

assign xor_ln1545_265_fu_8659_p2 = (tmp_V_86_reg_13118 ^ tmp_V_85_reg_13088);

assign xor_ln1545_266_fu_8669_p2 = (xor_ln1545_267_fu_8663_p2 ^ xor_ln1545_265_fu_8659_p2);

assign xor_ln1545_267_fu_8663_p2 = (trunc_ln674_87_fu_8421_p1 ^ tmp_177_fu_8383_p4);

assign xor_ln1545_268_fu_8675_p2 = (tmp_V_91_reg_13076 ^ tmp_2_1_V_15_reg_13046);

assign xor_ln1545_269_fu_8685_p2 = (xor_ln1545_270_fu_8679_p2 ^ xor_ln1545_268_fu_8675_p2);

assign xor_ln1545_26_fu_4494_p2 = (xor_ln1545_27_fu_4488_p2 ^ xor_ln1545_25_fu_4484_p2);

assign xor_ln1545_270_fu_8679_p2 = (trunc_ln674_88_fu_8435_p1 ^ tmp_182_fu_8453_p4);

assign xor_ln1545_271_fu_8691_p2 = (tmp_V_91_reg_13076 ^ tmp_V_88_reg_13082);

assign xor_ln1545_272_fu_8701_p2 = (xor_ln1545_273_fu_8695_p2 ^ xor_ln1545_271_fu_8691_p2);

assign xor_ln1545_273_fu_8695_p2 = (trunc_ln674_89_fu_8449_p1 ^ tmp_183_fu_8467_p4);

assign xor_ln1545_274_fu_8707_p2 = (tmp_V_89_reg_13112 ^ tmp_V_88_reg_13082);

assign xor_ln1545_275_fu_8717_p2 = (xor_ln1545_276_fu_8711_p2 ^ xor_ln1545_274_fu_8707_p2);

assign xor_ln1545_276_fu_8711_p2 = (trunc_ln674_90_fu_8463_p1 ^ tmp_184_fu_8481_p4);

assign xor_ln1545_277_fu_8723_p2 = (tmp_V_89_reg_13112 ^ tmp_2_1_V_15_reg_13046);

assign xor_ln1545_278_fu_8733_p2 = (xor_ln1545_279_fu_8727_p2 ^ xor_ln1545_277_fu_8723_p2);

assign xor_ln1545_279_fu_8727_p2 = (trunc_ln674_91_fu_8477_p1 ^ tmp_181_fu_8439_p4);

assign xor_ln1545_27_fu_4488_p2 = (trunc_ln674_7_fu_4246_p1 ^ tmp_22_fu_4208_p4);

assign xor_ln1545_280_fu_8739_p2 = (tmp_V_95_reg_13100 ^ tmp_2_2_V_15_reg_13070);

assign xor_ln1545_281_fu_8749_p2 = (xor_ln1545_282_fu_8743_p2 ^ xor_ln1545_280_fu_8739_p2);

assign xor_ln1545_282_fu_8743_p2 = (trunc_ln674_92_fu_8491_p1 ^ tmp_186_fu_8509_p4);

assign xor_ln1545_283_fu_8755_p2 = (tmp_V_95_reg_13100 ^ tmp_V_92_reg_13106);

assign xor_ln1545_284_fu_8765_p2 = (xor_ln1545_285_fu_8759_p2 ^ xor_ln1545_283_fu_8755_p2);

assign xor_ln1545_285_fu_8759_p2 = (trunc_ln674_93_fu_8505_p1 ^ tmp_187_fu_8523_p4);

assign xor_ln1545_286_fu_8771_p2 = (tmp_V_92_reg_13106 ^ tmp_1_V_15_reg_13040);

assign xor_ln1545_287_fu_8781_p2 = (xor_ln1545_288_fu_8775_p2 ^ xor_ln1545_286_fu_8771_p2);

assign xor_ln1545_288_fu_8775_p2 = (trunc_ln674_94_fu_8519_p1 ^ tmp_188_fu_8537_p4);

assign xor_ln1545_289_fu_8787_p2 = (tmp_2_2_V_15_reg_13070 ^ tmp_1_V_15_reg_13040);

assign xor_ln1545_28_fu_4500_p2 = (tmp_V_11_reg_11796 ^ tmp_2_1_V_10_reg_11766);

assign xor_ln1545_290_fu_8797_p2 = (xor_ln1545_291_fu_8791_p2 ^ xor_ln1545_289_fu_8787_p2);

assign xor_ln1545_291_fu_8791_p2 = (trunc_ln674_95_fu_8533_p1 ^ tmp_185_fu_8495_p4);

assign xor_ln1545_292_fu_9382_p2 = (tmp_V_98_reg_13350 ^ tmp_3_V_16_reg_13380);

assign xor_ln1545_293_fu_9392_p2 = (xor_ln1545_294_fu_9386_p2 ^ xor_ln1545_292_fu_9382_p2);

assign xor_ln1545_294_fu_9386_p2 = (trunc_ln674_96_fu_9158_p1 ^ tmp_205_fu_9176_p4);

assign xor_ln1545_295_fu_9398_p2 = (tmp_V_96_reg_13290 ^ tmp_3_V_16_reg_13380);

assign xor_ln1545_296_fu_9408_p2 = (xor_ln1545_297_fu_9402_p2 ^ xor_ln1545_295_fu_9398_p2);

assign xor_ln1545_297_fu_9402_p2 = (trunc_ln674_97_fu_9172_p1 ^ tmp_206_fu_9190_p4);

assign xor_ln1545_298_fu_9414_p2 = (tmp_V_97_reg_13320 ^ tmp_V_96_reg_13290);

assign xor_ln1545_299_fu_9424_p2 = (xor_ln1545_300_fu_9418_p2 ^ xor_ln1545_298_fu_9414_p2);

assign xor_ln1545_29_fu_4510_p2 = (xor_ln1545_30_fu_4504_p2 ^ xor_ln1545_28_fu_4500_p2);

assign xor_ln1545_300_fu_9418_p2 = (trunc_ln674_98_fu_9186_p1 ^ tmp_207_fu_9204_p4);

assign xor_ln1545_301_fu_9430_p2 = (tmp_V_98_reg_13350 ^ tmp_V_97_reg_13320);

assign xor_ln1545_302_fu_9440_p2 = (xor_ln1545_303_fu_9434_p2 ^ xor_ln1545_301_fu_9430_p2);

assign xor_ln1545_303_fu_9434_p2 = (trunc_ln674_99_fu_9200_p1 ^ tmp_204_fu_9162_p4);

assign xor_ln1545_304_fu_9446_p2 = (tmp_V_103_reg_13308 ^ tmp_V_102_reg_13374);

assign xor_ln1545_305_fu_9456_p2 = (xor_ln1545_306_fu_9450_p2 ^ xor_ln1545_304_fu_9446_p2);

assign xor_ln1545_306_fu_9450_p2 = (trunc_ln674_100_fu_9214_p1 ^ tmp_209_fu_9232_p4);

assign xor_ln1545_307_fu_9462_p2 = (tmp_V_103_reg_13308 ^ tmp_V_100_reg_13314);

assign xor_ln1545_308_fu_9472_p2 = (xor_ln1545_309_fu_9466_p2 ^ xor_ln1545_307_fu_9462_p2);

assign xor_ln1545_309_fu_9466_p2 = (trunc_ln674_101_fu_9228_p1 ^ tmp_210_fu_9246_p4);

assign xor_ln1545_30_fu_4504_p2 = (trunc_ln674_8_fu_4260_p1 ^ tmp_27_fu_4278_p4);

assign xor_ln1545_310_fu_9478_p2 = (tmp_V_101_reg_13344 ^ tmp_V_100_reg_13314);

assign xor_ln1545_311_fu_9488_p2 = (xor_ln1545_312_fu_9482_p2 ^ xor_ln1545_310_fu_9478_p2);

assign xor_ln1545_312_fu_9482_p2 = (trunc_ln674_102_fu_9242_p1 ^ tmp_211_fu_9260_p4);

assign xor_ln1545_313_fu_9494_p2 = (tmp_V_102_reg_13374 ^ tmp_V_101_reg_13344);

assign xor_ln1545_314_fu_9504_p2 = (xor_ln1545_315_fu_9498_p2 ^ xor_ln1545_313_fu_9494_p2);

assign xor_ln1545_315_fu_9498_p2 = (trunc_ln674_103_fu_9256_p1 ^ tmp_208_fu_9218_p4);

assign xor_ln1545_316_fu_9510_p2 = (tmp_V_107_reg_13332 ^ tmp_2_1_V_16_reg_13302);

assign xor_ln1545_317_fu_9520_p2 = (xor_ln1545_318_fu_9514_p2 ^ xor_ln1545_316_fu_9510_p2);

assign xor_ln1545_318_fu_9514_p2 = (trunc_ln674_104_fu_9270_p1 ^ tmp_213_fu_9288_p4);

assign xor_ln1545_319_fu_9526_p2 = (tmp_V_107_reg_13332 ^ tmp_V_104_reg_13338);

assign xor_ln1545_31_fu_4516_p2 = (tmp_V_8_reg_11802 ^ tmp_V_11_reg_11796);

assign xor_ln1545_320_fu_9536_p2 = (xor_ln1545_321_fu_9530_p2 ^ xor_ln1545_319_fu_9526_p2);

assign xor_ln1545_321_fu_9530_p2 = (trunc_ln674_105_fu_9284_p1 ^ tmp_214_fu_9302_p4);

assign xor_ln1545_322_fu_9542_p2 = (tmp_V_105_reg_13368 ^ tmp_V_104_reg_13338);

assign xor_ln1545_323_fu_9552_p2 = (xor_ln1545_324_fu_9546_p2 ^ xor_ln1545_322_fu_9542_p2);

assign xor_ln1545_324_fu_9546_p2 = (trunc_ln674_106_fu_9298_p1 ^ tmp_215_fu_9316_p4);

assign xor_ln1545_325_fu_9558_p2 = (tmp_V_105_reg_13368 ^ tmp_2_1_V_16_reg_13302);

assign xor_ln1545_326_fu_9568_p2 = (xor_ln1545_327_fu_9562_p2 ^ xor_ln1545_325_fu_9558_p2);

assign xor_ln1545_327_fu_9562_p2 = (trunc_ln674_107_fu_9312_p1 ^ tmp_212_fu_9274_p4);

assign xor_ln1545_328_fu_9574_p2 = (tmp_V_111_reg_13356 ^ tmp_2_2_V_16_reg_13326);

assign xor_ln1545_329_fu_9584_p2 = (xor_ln1545_330_fu_9578_p2 ^ xor_ln1545_328_fu_9574_p2);

assign xor_ln1545_32_fu_4526_p2 = (xor_ln1545_33_fu_4520_p2 ^ xor_ln1545_31_fu_4516_p2);

assign xor_ln1545_330_fu_9578_p2 = (trunc_ln674_108_fu_9326_p1 ^ tmp_217_fu_9344_p4);

assign xor_ln1545_331_fu_9590_p2 = (tmp_V_111_reg_13356 ^ tmp_V_108_reg_13362);

assign xor_ln1545_332_fu_9600_p2 = (xor_ln1545_333_fu_9594_p2 ^ xor_ln1545_331_fu_9590_p2);

assign xor_ln1545_333_fu_9594_p2 = (trunc_ln674_109_fu_9340_p1 ^ tmp_218_fu_9358_p4);

assign xor_ln1545_334_fu_9606_p2 = (tmp_V_108_reg_13362 ^ tmp_1_V_16_reg_13296);

assign xor_ln1545_335_fu_9616_p2 = (xor_ln1545_336_fu_9610_p2 ^ xor_ln1545_334_fu_9606_p2);

assign xor_ln1545_336_fu_9610_p2 = (trunc_ln674_110_fu_9354_p1 ^ tmp_219_fu_9372_p4);

assign xor_ln1545_337_fu_9622_p2 = (tmp_2_2_V_16_reg_13326 ^ tmp_1_V_16_reg_13296);

assign xor_ln1545_338_fu_9632_p2 = (xor_ln1545_339_fu_9626_p2 ^ xor_ln1545_337_fu_9622_p2);

assign xor_ln1545_339_fu_9626_p2 = (trunc_ln674_111_fu_9368_p1 ^ tmp_216_fu_9330_p4);

assign xor_ln1545_33_fu_4520_p2 = (trunc_ln674_9_fu_4274_p1 ^ tmp_28_fu_4292_p4);

assign xor_ln1545_340_fu_10217_p2 = (tmp_V_114_reg_13606 ^ tmp_3_V_17_reg_13636);

assign xor_ln1545_341_fu_10227_p2 = (xor_ln1545_342_fu_10221_p2 ^ xor_ln1545_340_fu_10217_p2);

assign xor_ln1545_342_fu_10221_p2 = (trunc_ln674_112_fu_9993_p1 ^ tmp_236_fu_10011_p4);

assign xor_ln1545_343_fu_10233_p2 = (tmp_V_112_reg_13546 ^ tmp_3_V_17_reg_13636);

assign xor_ln1545_344_fu_10243_p2 = (xor_ln1545_345_fu_10237_p2 ^ xor_ln1545_343_fu_10233_p2);

assign xor_ln1545_345_fu_10237_p2 = (trunc_ln674_113_fu_10007_p1 ^ tmp_237_fu_10025_p4);

assign xor_ln1545_346_fu_10249_p2 = (tmp_V_113_reg_13576 ^ tmp_V_112_reg_13546);

assign xor_ln1545_347_fu_10259_p2 = (xor_ln1545_348_fu_10253_p2 ^ xor_ln1545_346_fu_10249_p2);

assign xor_ln1545_348_fu_10253_p2 = (trunc_ln674_114_fu_10021_p1 ^ tmp_238_fu_10039_p4);

assign xor_ln1545_349_fu_10265_p2 = (tmp_V_114_reg_13606 ^ tmp_V_113_reg_13576);

assign xor_ln1545_34_fu_4532_p2 = (tmp_V_9_reg_11832 ^ tmp_V_8_reg_11802);

assign xor_ln1545_350_fu_10275_p2 = (xor_ln1545_351_fu_10269_p2 ^ xor_ln1545_349_fu_10265_p2);

assign xor_ln1545_351_fu_10269_p2 = (trunc_ln674_115_fu_10035_p1 ^ tmp_235_fu_9997_p4);

assign xor_ln1545_352_fu_10281_p2 = (tmp_V_119_reg_13564 ^ tmp_V_118_reg_13630);

assign xor_ln1545_353_fu_10291_p2 = (xor_ln1545_354_fu_10285_p2 ^ xor_ln1545_352_fu_10281_p2);

assign xor_ln1545_354_fu_10285_p2 = (trunc_ln674_116_fu_10049_p1 ^ tmp_240_fu_10067_p4);

assign xor_ln1545_355_fu_10297_p2 = (tmp_V_119_reg_13564 ^ tmp_V_116_reg_13570);

assign xor_ln1545_356_fu_10307_p2 = (xor_ln1545_357_fu_10301_p2 ^ xor_ln1545_355_fu_10297_p2);

assign xor_ln1545_357_fu_10301_p2 = (trunc_ln674_117_fu_10063_p1 ^ tmp_241_fu_10081_p4);

assign xor_ln1545_358_fu_10313_p2 = (tmp_V_117_reg_13600 ^ tmp_V_116_reg_13570);

assign xor_ln1545_359_fu_10323_p2 = (xor_ln1545_360_fu_10317_p2 ^ xor_ln1545_358_fu_10313_p2);

assign xor_ln1545_35_fu_4542_p2 = (xor_ln1545_36_fu_4536_p2 ^ xor_ln1545_34_fu_4532_p2);

assign xor_ln1545_360_fu_10317_p2 = (trunc_ln674_118_fu_10077_p1 ^ tmp_242_fu_10095_p4);

assign xor_ln1545_361_fu_10329_p2 = (tmp_V_118_reg_13630 ^ tmp_V_117_reg_13600);

assign xor_ln1545_362_fu_10339_p2 = (xor_ln1545_363_fu_10333_p2 ^ xor_ln1545_361_fu_10329_p2);

assign xor_ln1545_363_fu_10333_p2 = (trunc_ln674_119_fu_10091_p1 ^ tmp_239_fu_10053_p4);

assign xor_ln1545_364_fu_10345_p2 = (tmp_V_123_reg_13588 ^ tmp_2_1_V_17_reg_13558);

assign xor_ln1545_365_fu_10355_p2 = (xor_ln1545_366_fu_10349_p2 ^ xor_ln1545_364_fu_10345_p2);

assign xor_ln1545_366_fu_10349_p2 = (trunc_ln674_120_fu_10105_p1 ^ tmp_244_fu_10123_p4);

assign xor_ln1545_367_fu_10361_p2 = (tmp_V_123_reg_13588 ^ tmp_V_120_reg_13594);

assign xor_ln1545_368_fu_10371_p2 = (xor_ln1545_369_fu_10365_p2 ^ xor_ln1545_367_fu_10361_p2);

assign xor_ln1545_369_fu_10365_p2 = (trunc_ln674_121_fu_10119_p1 ^ tmp_245_fu_10137_p4);

assign xor_ln1545_36_fu_4536_p2 = (trunc_ln674_10_fu_4288_p1 ^ tmp_29_fu_4306_p4);

assign xor_ln1545_370_fu_10377_p2 = (tmp_V_121_reg_13624 ^ tmp_V_120_reg_13594);

assign xor_ln1545_371_fu_10387_p2 = (xor_ln1545_372_fu_10381_p2 ^ xor_ln1545_370_fu_10377_p2);

assign xor_ln1545_372_fu_10381_p2 = (trunc_ln674_122_fu_10133_p1 ^ tmp_246_fu_10151_p4);

assign xor_ln1545_373_fu_10393_p2 = (tmp_V_121_reg_13624 ^ tmp_2_1_V_17_reg_13558);

assign xor_ln1545_374_fu_10403_p2 = (xor_ln1545_375_fu_10397_p2 ^ xor_ln1545_373_fu_10393_p2);

assign xor_ln1545_375_fu_10397_p2 = (trunc_ln674_123_fu_10147_p1 ^ tmp_243_fu_10109_p4);

assign xor_ln1545_376_fu_10409_p2 = (tmp_V_127_reg_13612 ^ tmp_2_2_V_17_reg_13582);

assign xor_ln1545_377_fu_10419_p2 = (xor_ln1545_378_fu_10413_p2 ^ xor_ln1545_376_fu_10409_p2);

assign xor_ln1545_378_fu_10413_p2 = (trunc_ln674_124_fu_10161_p1 ^ tmp_248_fu_10179_p4);

assign xor_ln1545_379_fu_10425_p2 = (tmp_V_127_reg_13612 ^ tmp_V_124_reg_13618);

assign xor_ln1545_37_fu_4548_p2 = (tmp_V_9_reg_11832 ^ tmp_2_1_V_10_reg_11766);

assign xor_ln1545_380_fu_10435_p2 = (xor_ln1545_381_fu_10429_p2 ^ xor_ln1545_379_fu_10425_p2);

assign xor_ln1545_381_fu_10429_p2 = (trunc_ln674_125_fu_10175_p1 ^ tmp_249_fu_10193_p4);

assign xor_ln1545_382_fu_10441_p2 = (tmp_V_124_reg_13618 ^ tmp_1_V_17_reg_13552);

assign xor_ln1545_383_fu_10451_p2 = (xor_ln1545_384_fu_10445_p2 ^ xor_ln1545_382_fu_10441_p2);

assign xor_ln1545_384_fu_10445_p2 = (trunc_ln674_126_fu_10189_p1 ^ tmp_250_fu_10207_p4);

assign xor_ln1545_385_fu_10457_p2 = (tmp_2_2_V_17_reg_13582 ^ tmp_1_V_17_reg_13552);

assign xor_ln1545_386_fu_10467_p2 = (xor_ln1545_387_fu_10461_p2 ^ xor_ln1545_385_fu_10457_p2);

assign xor_ln1545_387_fu_10461_p2 = (trunc_ln674_127_fu_10203_p1 ^ tmp_247_fu_10165_p4);

assign xor_ln1545_388_fu_11052_p2 = (tmp_V_130_reg_13862 ^ tmp_3_V_18_reg_13892);

assign xor_ln1545_389_fu_11062_p2 = (xor_ln1545_390_fu_11056_p2 ^ xor_ln1545_388_fu_11052_p2);

assign xor_ln1545_38_fu_4558_p2 = (xor_ln1545_39_fu_4552_p2 ^ xor_ln1545_37_fu_4548_p2);

assign xor_ln1545_390_fu_11056_p2 = (trunc_ln674_128_fu_10828_p1 ^ tmp_267_fu_10846_p4);

assign xor_ln1545_391_fu_11068_p2 = (tmp_V_128_reg_13802 ^ tmp_3_V_18_reg_13892);

assign xor_ln1545_392_fu_11078_p2 = (xor_ln1545_393_fu_11072_p2 ^ xor_ln1545_391_fu_11068_p2);

assign xor_ln1545_393_fu_11072_p2 = (trunc_ln674_129_fu_10842_p1 ^ tmp_268_fu_10860_p4);

assign xor_ln1545_394_fu_11084_p2 = (tmp_V_129_reg_13832 ^ tmp_V_128_reg_13802);

assign xor_ln1545_395_fu_11094_p2 = (xor_ln1545_396_fu_11088_p2 ^ xor_ln1545_394_fu_11084_p2);

assign xor_ln1545_396_fu_11088_p2 = (trunc_ln674_130_fu_10856_p1 ^ tmp_269_fu_10874_p4);

assign xor_ln1545_397_fu_11100_p2 = (tmp_V_130_reg_13862 ^ tmp_V_129_reg_13832);

assign xor_ln1545_398_fu_11110_p2 = (xor_ln1545_399_fu_11104_p2 ^ xor_ln1545_397_fu_11100_p2);

assign xor_ln1545_399_fu_11104_p2 = (trunc_ln674_131_fu_10870_p1 ^ tmp_266_fu_10832_p4);

assign xor_ln1545_39_fu_4552_p2 = (trunc_ln674_11_fu_4302_p1 ^ tmp_26_fu_4264_p4);

assign xor_ln1545_400_fu_11116_p2 = (tmp_V_135_reg_13820 ^ tmp_V_134_reg_13886);

assign xor_ln1545_401_fu_11126_p2 = (xor_ln1545_402_fu_11120_p2 ^ xor_ln1545_400_fu_11116_p2);

assign xor_ln1545_402_fu_11120_p2 = (trunc_ln674_132_fu_10884_p1 ^ tmp_271_fu_10902_p4);

assign xor_ln1545_403_fu_11132_p2 = (tmp_V_135_reg_13820 ^ tmp_V_132_reg_13826);

assign xor_ln1545_404_fu_11142_p2 = (xor_ln1545_405_fu_11136_p2 ^ xor_ln1545_403_fu_11132_p2);

assign xor_ln1545_405_fu_11136_p2 = (trunc_ln674_133_fu_10898_p1 ^ tmp_272_fu_10916_p4);

assign xor_ln1545_406_fu_11148_p2 = (tmp_V_133_reg_13856 ^ tmp_V_132_reg_13826);

assign xor_ln1545_407_fu_11158_p2 = (xor_ln1545_408_fu_11152_p2 ^ xor_ln1545_406_fu_11148_p2);

assign xor_ln1545_408_fu_11152_p2 = (trunc_ln674_134_fu_10912_p1 ^ tmp_273_fu_10930_p4);

assign xor_ln1545_409_fu_11164_p2 = (tmp_V_134_reg_13886 ^ tmp_V_133_reg_13856);

assign xor_ln1545_40_fu_4564_p2 = (tmp_V_15_reg_11820 ^ tmp_2_2_V_10_reg_11790);

assign xor_ln1545_410_fu_11174_p2 = (xor_ln1545_411_fu_11168_p2 ^ xor_ln1545_409_fu_11164_p2);

assign xor_ln1545_411_fu_11168_p2 = (trunc_ln674_135_fu_10926_p1 ^ tmp_270_fu_10888_p4);

assign xor_ln1545_412_fu_11180_p2 = (tmp_V_139_reg_13844 ^ tmp_2_1_V_18_reg_13814);

assign xor_ln1545_413_fu_11190_p2 = (xor_ln1545_414_fu_11184_p2 ^ xor_ln1545_412_fu_11180_p2);

assign xor_ln1545_414_fu_11184_p2 = (trunc_ln674_136_fu_10940_p1 ^ tmp_275_fu_10958_p4);

assign xor_ln1545_415_fu_11196_p2 = (tmp_V_139_reg_13844 ^ tmp_V_136_reg_13850);

assign xor_ln1545_416_fu_11206_p2 = (xor_ln1545_417_fu_11200_p2 ^ xor_ln1545_415_fu_11196_p2);

assign xor_ln1545_417_fu_11200_p2 = (trunc_ln674_137_fu_10954_p1 ^ tmp_276_fu_10972_p4);

assign xor_ln1545_418_fu_11212_p2 = (tmp_V_137_reg_13880 ^ tmp_V_136_reg_13850);

assign xor_ln1545_419_fu_11222_p2 = (xor_ln1545_420_fu_11216_p2 ^ xor_ln1545_418_fu_11212_p2);

assign xor_ln1545_41_fu_4574_p2 = (xor_ln1545_42_fu_4568_p2 ^ xor_ln1545_40_fu_4564_p2);

assign xor_ln1545_420_fu_11216_p2 = (trunc_ln674_138_fu_10968_p1 ^ tmp_277_fu_10986_p4);

assign xor_ln1545_421_fu_11228_p2 = (tmp_V_137_reg_13880 ^ tmp_2_1_V_18_reg_13814);

assign xor_ln1545_422_fu_11238_p2 = (xor_ln1545_423_fu_11232_p2 ^ xor_ln1545_421_fu_11228_p2);

assign xor_ln1545_423_fu_11232_p2 = (trunc_ln674_139_fu_10982_p1 ^ tmp_274_fu_10944_p4);

assign xor_ln1545_424_fu_11244_p2 = (tmp_V_143_reg_13868 ^ tmp_2_2_V_18_reg_13838);

assign xor_ln1545_425_fu_11254_p2 = (xor_ln1545_426_fu_11248_p2 ^ xor_ln1545_424_fu_11244_p2);

assign xor_ln1545_426_fu_11248_p2 = (trunc_ln674_140_fu_10996_p1 ^ tmp_279_fu_11014_p4);

assign xor_ln1545_427_fu_11260_p2 = (tmp_V_143_reg_13868 ^ tmp_V_140_reg_13874);

assign xor_ln1545_428_fu_11270_p2 = (xor_ln1545_429_fu_11264_p2 ^ xor_ln1545_427_fu_11260_p2);

assign xor_ln1545_429_fu_11264_p2 = (trunc_ln674_141_fu_11010_p1 ^ tmp_280_fu_11028_p4);

assign xor_ln1545_42_fu_4568_p2 = (trunc_ln674_12_fu_4316_p1 ^ tmp_31_fu_4334_p4);

assign xor_ln1545_430_fu_11276_p2 = (tmp_V_140_reg_13874 ^ tmp_1_V_18_reg_13808);

assign xor_ln1545_431_fu_11286_p2 = (xor_ln1545_432_fu_11280_p2 ^ xor_ln1545_430_fu_11276_p2);

assign xor_ln1545_432_fu_11280_p2 = (trunc_ln674_142_fu_11024_p1 ^ tmp_281_fu_11042_p4);

assign xor_ln1545_433_fu_11292_p2 = (tmp_2_2_V_18_reg_13838 ^ tmp_1_V_18_reg_13808);

assign xor_ln1545_434_fu_11302_p2 = (xor_ln1545_435_fu_11296_p2 ^ xor_ln1545_433_fu_11292_p2);

assign xor_ln1545_435_fu_11296_p2 = (trunc_ln674_143_fu_11038_p1 ^ tmp_278_fu_11000_p4);

assign xor_ln1545_43_fu_4580_p2 = (tmp_V_15_reg_11820 ^ tmp_V_12_reg_11826);

assign xor_ln1545_44_fu_4590_p2 = (xor_ln1545_45_fu_4584_p2 ^ xor_ln1545_43_fu_4580_p2);

assign xor_ln1545_45_fu_4584_p2 = (trunc_ln674_13_fu_4330_p1 ^ tmp_32_fu_4348_p4);

assign xor_ln1545_46_fu_4596_p2 = (tmp_V_12_reg_11826 ^ tmp_1_V_10_reg_11760);

assign xor_ln1545_47_fu_4606_p2 = (xor_ln1545_48_fu_4600_p2 ^ xor_ln1545_46_fu_4596_p2);

assign xor_ln1545_48_fu_4600_p2 = (trunc_ln674_14_fu_4344_p1 ^ tmp_33_fu_4362_p4);

assign xor_ln1545_49_fu_4612_p2 = (tmp_2_2_V_10_reg_11790 ^ tmp_1_V_10_reg_11760);

assign xor_ln1545_50_fu_4622_p2 = (xor_ln1545_51_fu_4616_p2 ^ xor_ln1545_49_fu_4612_p2);

assign xor_ln1545_51_fu_4616_p2 = (trunc_ln674_15_fu_4358_p1 ^ tmp_30_fu_4320_p4);

assign xor_ln1545_52_fu_5207_p2 = (tmp_V_18_reg_12070 ^ tmp_3_V_11_reg_12100);

assign xor_ln1545_53_fu_5217_p2 = (xor_ln1545_54_fu_5211_p2 ^ xor_ln1545_52_fu_5207_p2);

assign xor_ln1545_54_fu_5211_p2 = (trunc_ln674_16_fu_4983_p1 ^ tmp_50_fu_5001_p4);

assign xor_ln1545_55_fu_5223_p2 = (tmp_V_16_reg_12010 ^ tmp_3_V_11_reg_12100);

assign xor_ln1545_56_fu_5233_p2 = (xor_ln1545_57_fu_5227_p2 ^ xor_ln1545_55_fu_5223_p2);

assign xor_ln1545_57_fu_5227_p2 = (trunc_ln674_17_fu_4997_p1 ^ tmp_51_fu_5015_p4);

assign xor_ln1545_58_fu_5239_p2 = (tmp_V_17_reg_12040 ^ tmp_V_16_reg_12010);

assign xor_ln1545_59_fu_5249_p2 = (xor_ln1545_60_fu_5243_p2 ^ xor_ln1545_58_fu_5239_p2);

assign xor_ln1545_5_fu_4382_p2 = (xor_ln1545_fu_4372_p2 ^ xor_ln1545_6_fu_4376_p2);

assign xor_ln1545_60_fu_5243_p2 = (trunc_ln674_18_fu_5011_p1 ^ tmp_52_fu_5029_p4);

assign xor_ln1545_61_fu_5255_p2 = (tmp_V_18_reg_12070 ^ tmp_V_17_reg_12040);

assign xor_ln1545_62_fu_5265_p2 = (xor_ln1545_63_fu_5259_p2 ^ xor_ln1545_61_fu_5255_p2);

assign xor_ln1545_63_fu_5259_p2 = (trunc_ln674_19_fu_5025_p1 ^ tmp_49_fu_4987_p4);

assign xor_ln1545_64_fu_5271_p2 = (tmp_V_23_reg_12028 ^ tmp_V_22_reg_12094);

assign xor_ln1545_65_fu_5281_p2 = (xor_ln1545_66_fu_5275_p2 ^ xor_ln1545_64_fu_5271_p2);

assign xor_ln1545_66_fu_5275_p2 = (trunc_ln674_20_fu_5039_p1 ^ tmp_54_fu_5057_p4);

assign xor_ln1545_67_fu_5287_p2 = (tmp_V_23_reg_12028 ^ tmp_V_20_reg_12034);

assign xor_ln1545_68_fu_5297_p2 = (xor_ln1545_69_fu_5291_p2 ^ xor_ln1545_67_fu_5287_p2);

assign xor_ln1545_69_fu_5291_p2 = (trunc_ln674_21_fu_5053_p1 ^ tmp_55_fu_5071_p4);

assign xor_ln1545_6_fu_4376_p2 = (trunc_ln674_fu_4148_p1 ^ tmp_19_fu_4166_p4);

assign xor_ln1545_70_fu_5303_p2 = (tmp_V_21_reg_12064 ^ tmp_V_20_reg_12034);

assign xor_ln1545_71_fu_5313_p2 = (xor_ln1545_72_fu_5307_p2 ^ xor_ln1545_70_fu_5303_p2);

assign xor_ln1545_72_fu_5307_p2 = (trunc_ln674_22_fu_5067_p1 ^ tmp_56_fu_5085_p4);

assign xor_ln1545_73_fu_5319_p2 = (tmp_V_22_reg_12094 ^ tmp_V_21_reg_12064);

assign xor_ln1545_74_fu_5329_p2 = (xor_ln1545_75_fu_5323_p2 ^ xor_ln1545_73_fu_5319_p2);

assign xor_ln1545_75_fu_5323_p2 = (trunc_ln674_23_fu_5081_p1 ^ tmp_53_fu_5043_p4);

assign xor_ln1545_76_fu_5335_p2 = (tmp_V_27_reg_12052 ^ tmp_2_1_V_11_reg_12022);

assign xor_ln1545_77_fu_5345_p2 = (xor_ln1545_78_fu_5339_p2 ^ xor_ln1545_76_fu_5335_p2);

assign xor_ln1545_78_fu_5339_p2 = (trunc_ln674_24_fu_5095_p1 ^ tmp_58_fu_5113_p4);

assign xor_ln1545_79_fu_5351_p2 = (tmp_V_27_reg_12052 ^ tmp_V_24_reg_12058);

assign xor_ln1545_7_fu_4388_p2 = (tmp_V_reg_11754 ^ tmp_3_V_10_reg_11844);

assign xor_ln1545_80_fu_5361_p2 = (xor_ln1545_81_fu_5355_p2 ^ xor_ln1545_79_fu_5351_p2);

assign xor_ln1545_81_fu_5355_p2 = (trunc_ln674_25_fu_5109_p1 ^ tmp_59_fu_5127_p4);

assign xor_ln1545_82_fu_5367_p2 = (tmp_V_25_reg_12088 ^ tmp_V_24_reg_12058);

assign xor_ln1545_83_fu_5377_p2 = (xor_ln1545_84_fu_5371_p2 ^ xor_ln1545_82_fu_5367_p2);

assign xor_ln1545_84_fu_5371_p2 = (trunc_ln674_26_fu_5123_p1 ^ tmp_60_fu_5141_p4);

assign xor_ln1545_85_fu_5383_p2 = (tmp_V_25_reg_12088 ^ tmp_2_1_V_11_reg_12022);

assign xor_ln1545_86_fu_5393_p2 = (xor_ln1545_87_fu_5387_p2 ^ xor_ln1545_85_fu_5383_p2);

assign xor_ln1545_87_fu_5387_p2 = (trunc_ln674_27_fu_5137_p1 ^ tmp_57_fu_5099_p4);

assign xor_ln1545_88_fu_5399_p2 = (tmp_V_31_reg_12076 ^ tmp_2_2_V_11_reg_12046);

assign xor_ln1545_89_fu_5409_p2 = (xor_ln1545_90_fu_5403_p2 ^ xor_ln1545_88_fu_5399_p2);

assign xor_ln1545_8_fu_4398_p2 = (xor_ln1545_9_fu_4392_p2 ^ xor_ln1545_7_fu_4388_p2);

assign xor_ln1545_90_fu_5403_p2 = (trunc_ln674_28_fu_5151_p1 ^ tmp_62_fu_5169_p4);

assign xor_ln1545_91_fu_5415_p2 = (tmp_V_31_reg_12076 ^ tmp_V_28_reg_12082);

assign xor_ln1545_92_fu_5425_p2 = (xor_ln1545_93_fu_5419_p2 ^ xor_ln1545_91_fu_5415_p2);

assign xor_ln1545_93_fu_5419_p2 = (trunc_ln674_29_fu_5165_p1 ^ tmp_63_fu_5183_p4);

assign xor_ln1545_94_fu_5431_p2 = (tmp_V_28_reg_12082 ^ tmp_1_V_11_reg_12016);

assign xor_ln1545_95_fu_5441_p2 = (xor_ln1545_96_fu_5435_p2 ^ xor_ln1545_94_fu_5431_p2);

assign xor_ln1545_96_fu_5435_p2 = (trunc_ln674_30_fu_5179_p1 ^ tmp_64_fu_5197_p4);

assign xor_ln1545_97_fu_5447_p2 = (tmp_2_2_V_11_reg_12046 ^ tmp_1_V_11_reg_12016);

assign xor_ln1545_98_fu_5457_p2 = (xor_ln1545_99_fu_5451_p2 ^ xor_ln1545_97_fu_5447_p2);

assign xor_ln1545_99_fu_5451_p2 = (trunc_ln674_31_fu_5193_p1 ^ tmp_61_fu_5155_p4);

assign xor_ln1545_9_fu_4392_p2 = (trunc_ln674_1_fu_4162_p1 ^ tmp_20_fu_4180_p4);

assign xor_ln1545_fu_4372_p2 = (tmp_V_2_reg_11814 ^ tmp_3_V_10_reg_11844);

assign zext_ln587_100_fu_9098_p1 = cipher_0_ssbox_q59;

assign zext_ln587_101_fu_9103_p1 = cipher_0_ssbox_q54;

assign zext_ln587_102_fu_9108_p1 = cipher_0_ssbox_q49;

assign zext_ln587_103_fu_9113_p1 = cipher_0_ssbox_q60;

assign zext_ln587_104_fu_9118_p1 = cipher_0_ssbox_q55;

assign zext_ln587_105_fu_9123_p1 = cipher_0_ssbox_q50;

assign zext_ln587_106_fu_9128_p1 = cipher_0_ssbox_q61;

assign zext_ln587_107_fu_9133_p1 = cipher_0_ssbox_q56;

assign zext_ln587_108_fu_9138_p1 = cipher_0_ssbox_q51;

assign zext_ln587_109_fu_9143_p1 = cipher_0_ssbox_q62;

assign zext_ln587_10_fu_4118_p1 = cipher_0_ssbox_q157;

assign zext_ln587_110_fu_9148_p1 = cipher_0_ssbox_q57;

assign zext_ln587_111_fu_9153_p1 = cipher_0_ssbox_q52;

assign zext_ln587_112_fu_9913_p1 = cipher_0_ssbox_q47;

assign zext_ln587_113_fu_9918_p1 = cipher_0_ssbox_q42;

assign zext_ln587_114_fu_9923_p1 = cipher_0_ssbox_q37;

assign zext_ln587_115_fu_9928_p1 = cipher_0_ssbox_q32;

assign zext_ln587_116_fu_9933_p1 = cipher_0_ssbox_q43;

assign zext_ln587_117_fu_9938_p1 = cipher_0_ssbox_q38;

assign zext_ln587_118_fu_9943_p1 = cipher_0_ssbox_q33;

assign zext_ln587_119_fu_9948_p1 = cipher_0_ssbox_q44;

assign zext_ln587_11_fu_4123_p1 = cipher_0_ssbox_q152;

assign zext_ln587_120_fu_9953_p1 = cipher_0_ssbox_q39;

assign zext_ln587_121_fu_9958_p1 = cipher_0_ssbox_q34;

assign zext_ln587_122_fu_9963_p1 = cipher_0_ssbox_q45;

assign zext_ln587_123_fu_9968_p1 = cipher_0_ssbox_q40;

assign zext_ln587_124_fu_9973_p1 = cipher_0_ssbox_q35;

assign zext_ln587_125_fu_9978_p1 = cipher_0_ssbox_q46;

assign zext_ln587_126_fu_9983_p1 = cipher_0_ssbox_q41;

assign zext_ln587_127_fu_9988_p1 = cipher_0_ssbox_q36;

assign zext_ln587_128_fu_10748_p1 = cipher_0_ssbox_q31;

assign zext_ln587_129_fu_10753_p1 = cipher_0_ssbox_q26;

assign zext_ln587_12_fu_4128_p1 = cipher_0_ssbox_q147;

assign zext_ln587_130_fu_10758_p1 = cipher_0_ssbox_q21;

assign zext_ln587_131_fu_10763_p1 = cipher_0_ssbox_q16;

assign zext_ln587_132_fu_10768_p1 = cipher_0_ssbox_q27;

assign zext_ln587_133_fu_10773_p1 = cipher_0_ssbox_q22;

assign zext_ln587_134_fu_10778_p1 = cipher_0_ssbox_q17;

assign zext_ln587_135_fu_10783_p1 = cipher_0_ssbox_q28;

assign zext_ln587_136_fu_10788_p1 = cipher_0_ssbox_q23;

assign zext_ln587_137_fu_10793_p1 = cipher_0_ssbox_q18;

assign zext_ln587_138_fu_10798_p1 = cipher_0_ssbox_q29;

assign zext_ln587_139_fu_10803_p1 = cipher_0_ssbox_q24;

assign zext_ln587_13_fu_4133_p1 = cipher_0_ssbox_q158;

assign zext_ln587_140_fu_10808_p1 = cipher_0_ssbox_q19;

assign zext_ln587_141_fu_10813_p1 = cipher_0_ssbox_q30;

assign zext_ln587_142_fu_10818_p1 = cipher_0_ssbox_q25;

assign zext_ln587_143_fu_10823_p1 = cipher_0_ssbox_q20;

assign zext_ln587_14_fu_4138_p1 = cipher_0_ssbox_q153;

assign zext_ln587_15_fu_4143_p1 = cipher_0_ssbox_q148;

assign zext_ln587_16_fu_4903_p1 = cipher_0_ssbox_q143;

assign zext_ln587_17_fu_4908_p1 = cipher_0_ssbox_q138;

assign zext_ln587_18_fu_4913_p1 = cipher_0_ssbox_q133;

assign zext_ln587_19_fu_4918_p1 = cipher_0_ssbox_q128;

assign zext_ln587_1_fu_4073_p1 = cipher_0_ssbox_q154;

assign zext_ln587_20_fu_4923_p1 = cipher_0_ssbox_q139;

assign zext_ln587_21_fu_4928_p1 = cipher_0_ssbox_q134;

assign zext_ln587_22_fu_4933_p1 = cipher_0_ssbox_q129;

assign zext_ln587_23_fu_4938_p1 = cipher_0_ssbox_q140;

assign zext_ln587_24_fu_4943_p1 = cipher_0_ssbox_q135;

assign zext_ln587_25_fu_4948_p1 = cipher_0_ssbox_q130;

assign zext_ln587_26_fu_4953_p1 = cipher_0_ssbox_q141;

assign zext_ln587_27_fu_4958_p1 = cipher_0_ssbox_q136;

assign zext_ln587_28_fu_4963_p1 = cipher_0_ssbox_q131;

assign zext_ln587_29_fu_4968_p1 = cipher_0_ssbox_q142;

assign zext_ln587_2_fu_4078_p1 = cipher_0_ssbox_q149;

assign zext_ln587_30_fu_4973_p1 = cipher_0_ssbox_q137;

assign zext_ln587_31_fu_4978_p1 = cipher_0_ssbox_q132;

assign zext_ln587_32_fu_5738_p1 = cipher_0_ssbox_q127;

assign zext_ln587_33_fu_5743_p1 = cipher_0_ssbox_q122;

assign zext_ln587_34_fu_5748_p1 = cipher_0_ssbox_q117;

assign zext_ln587_35_fu_5753_p1 = cipher_0_ssbox_q112;

assign zext_ln587_36_fu_5758_p1 = cipher_0_ssbox_q123;

assign zext_ln587_37_fu_5763_p1 = cipher_0_ssbox_q118;

assign zext_ln587_38_fu_5768_p1 = cipher_0_ssbox_q113;

assign zext_ln587_39_fu_5773_p1 = cipher_0_ssbox_q124;

assign zext_ln587_3_fu_4083_p1 = cipher_0_ssbox_q144;

assign zext_ln587_40_fu_5778_p1 = cipher_0_ssbox_q119;

assign zext_ln587_41_fu_5783_p1 = cipher_0_ssbox_q114;

assign zext_ln587_42_fu_5788_p1 = cipher_0_ssbox_q125;

assign zext_ln587_43_fu_5793_p1 = cipher_0_ssbox_q120;

assign zext_ln587_44_fu_5798_p1 = cipher_0_ssbox_q115;

assign zext_ln587_45_fu_5803_p1 = cipher_0_ssbox_q126;

assign zext_ln587_46_fu_5808_p1 = cipher_0_ssbox_q121;

assign zext_ln587_47_fu_5813_p1 = cipher_0_ssbox_q116;

assign zext_ln587_48_fu_6573_p1 = cipher_0_ssbox_q111;

assign zext_ln587_49_fu_6578_p1 = cipher_0_ssbox_q106;

assign zext_ln587_4_fu_4088_p1 = cipher_0_ssbox_q155;

assign zext_ln587_50_fu_6583_p1 = cipher_0_ssbox_q101;

assign zext_ln587_51_fu_6588_p1 = cipher_0_ssbox_q96;

assign zext_ln587_52_fu_6593_p1 = cipher_0_ssbox_q107;

assign zext_ln587_53_fu_6598_p1 = cipher_0_ssbox_q102;

assign zext_ln587_54_fu_6603_p1 = cipher_0_ssbox_q97;

assign zext_ln587_55_fu_6608_p1 = cipher_0_ssbox_q108;

assign zext_ln587_56_fu_6613_p1 = cipher_0_ssbox_q103;

assign zext_ln587_57_fu_6618_p1 = cipher_0_ssbox_q98;

assign zext_ln587_58_fu_6623_p1 = cipher_0_ssbox_q109;

assign zext_ln587_59_fu_6628_p1 = cipher_0_ssbox_q104;

assign zext_ln587_5_fu_4093_p1 = cipher_0_ssbox_q150;

assign zext_ln587_60_fu_6633_p1 = cipher_0_ssbox_q99;

assign zext_ln587_61_fu_6638_p1 = cipher_0_ssbox_q110;

assign zext_ln587_62_fu_6643_p1 = cipher_0_ssbox_q105;

assign zext_ln587_63_fu_6648_p1 = cipher_0_ssbox_q100;

assign zext_ln587_64_fu_7408_p1 = cipher_0_ssbox_q95;

assign zext_ln587_65_fu_7413_p1 = cipher_0_ssbox_q90;

assign zext_ln587_66_fu_7418_p1 = cipher_0_ssbox_q85;

assign zext_ln587_67_fu_7423_p1 = cipher_0_ssbox_q80;

assign zext_ln587_68_fu_7428_p1 = cipher_0_ssbox_q91;

assign zext_ln587_69_fu_7433_p1 = cipher_0_ssbox_q86;

assign zext_ln587_6_fu_4098_p1 = cipher_0_ssbox_q145;

assign zext_ln587_70_fu_7438_p1 = cipher_0_ssbox_q81;

assign zext_ln587_71_fu_7443_p1 = cipher_0_ssbox_q92;

assign zext_ln587_72_fu_7448_p1 = cipher_0_ssbox_q87;

assign zext_ln587_73_fu_7453_p1 = cipher_0_ssbox_q82;

assign zext_ln587_74_fu_7458_p1 = cipher_0_ssbox_q93;

assign zext_ln587_75_fu_7463_p1 = cipher_0_ssbox_q88;

assign zext_ln587_76_fu_7468_p1 = cipher_0_ssbox_q83;

assign zext_ln587_77_fu_7473_p1 = cipher_0_ssbox_q94;

assign zext_ln587_78_fu_7478_p1 = cipher_0_ssbox_q89;

assign zext_ln587_79_fu_7483_p1 = cipher_0_ssbox_q84;

assign zext_ln587_7_fu_4103_p1 = cipher_0_ssbox_q156;

assign zext_ln587_80_fu_8243_p1 = cipher_0_ssbox_q79;

assign zext_ln587_81_fu_8248_p1 = cipher_0_ssbox_q74;

assign zext_ln587_82_fu_8253_p1 = cipher_0_ssbox_q69;

assign zext_ln587_83_fu_8258_p1 = cipher_0_ssbox_q64;

assign zext_ln587_84_fu_8263_p1 = cipher_0_ssbox_q75;

assign zext_ln587_85_fu_8268_p1 = cipher_0_ssbox_q70;

assign zext_ln587_86_fu_8273_p1 = cipher_0_ssbox_q65;

assign zext_ln587_87_fu_8278_p1 = cipher_0_ssbox_q76;

assign zext_ln587_88_fu_8283_p1 = cipher_0_ssbox_q71;

assign zext_ln587_89_fu_8288_p1 = cipher_0_ssbox_q66;

assign zext_ln587_8_fu_4108_p1 = cipher_0_ssbox_q151;

assign zext_ln587_90_fu_8293_p1 = cipher_0_ssbox_q77;

assign zext_ln587_91_fu_8298_p1 = cipher_0_ssbox_q72;

assign zext_ln587_92_fu_8303_p1 = cipher_0_ssbox_q67;

assign zext_ln587_93_fu_8308_p1 = cipher_0_ssbox_q78;

assign zext_ln587_94_fu_8313_p1 = cipher_0_ssbox_q73;

assign zext_ln587_95_fu_8318_p1 = cipher_0_ssbox_q68;

assign zext_ln587_96_fu_9078_p1 = cipher_0_ssbox_q63;

assign zext_ln587_97_fu_9083_p1 = cipher_0_ssbox_q58;

assign zext_ln587_98_fu_9088_p1 = cipher_0_ssbox_q53;

assign zext_ln587_99_fu_9093_p1 = cipher_0_ssbox_q48;

assign zext_ln587_9_fu_4113_p1 = cipher_0_ssbox_q146;

assign zext_ln587_fu_4068_p1 = cipher_0_ssbox_q159;

assign zext_ln708_100_fu_8863_p1 = tmp_189_fu_8853_p4;

assign zext_ln708_101_fu_8878_p1 = tmp_190_fu_8868_p4;

assign zext_ln708_102_fu_8893_p1 = tmp_191_fu_8883_p4;

assign zext_ln708_103_fu_8908_p1 = tmp_192_fu_8898_p4;

assign zext_ln708_104_fu_8923_p1 = tmp_193_fu_8913_p4;

assign zext_ln708_105_fu_8938_p1 = tmp_194_fu_8928_p4;

assign zext_ln708_106_fu_8953_p1 = tmp_195_fu_8943_p4;

assign zext_ln708_107_fu_8968_p1 = tmp_196_fu_8958_p4;

assign zext_ln708_108_fu_8983_p1 = tmp_197_fu_8973_p4;

assign zext_ln708_109_fu_8998_p1 = tmp_198_fu_8988_p4;

assign zext_ln708_10_fu_3943_p1 = tmp_9_fu_3933_p4;

assign zext_ln708_110_fu_9013_p1 = tmp_199_fu_9003_p4;

assign zext_ln708_111_fu_9028_p1 = tmp_200_fu_9018_p4;

assign zext_ln708_112_fu_9043_p1 = tmp_201_fu_9033_p4;

assign zext_ln708_113_fu_9058_p1 = tmp_202_fu_9048_p4;

assign zext_ln708_114_fu_9073_p1 = tmp_203_fu_9063_p4;

assign zext_ln708_115_fu_9683_p1 = trunc_ln708_7_fu_9679_p1;

assign zext_ln708_116_fu_9698_p1 = tmp_220_fu_9688_p4;

assign zext_ln708_117_fu_9713_p1 = tmp_221_fu_9703_p4;

assign zext_ln708_118_fu_9728_p1 = tmp_222_fu_9718_p4;

assign zext_ln708_119_fu_9743_p1 = tmp_223_fu_9733_p4;

assign zext_ln708_11_fu_3958_p1 = tmp_10_fu_3948_p4;

assign zext_ln708_120_fu_9758_p1 = tmp_224_fu_9748_p4;

assign zext_ln708_121_fu_9773_p1 = tmp_225_fu_9763_p4;

assign zext_ln708_122_fu_9788_p1 = tmp_226_fu_9778_p4;

assign zext_ln708_123_fu_9803_p1 = tmp_227_fu_9793_p4;

assign zext_ln708_124_fu_9818_p1 = tmp_228_fu_9808_p4;

assign zext_ln708_125_fu_9833_p1 = tmp_229_fu_9823_p4;

assign zext_ln708_126_fu_9848_p1 = tmp_230_fu_9838_p4;

assign zext_ln708_127_fu_9863_p1 = tmp_231_fu_9853_p4;

assign zext_ln708_128_fu_9878_p1 = tmp_232_fu_9868_p4;

assign zext_ln708_129_fu_9893_p1 = tmp_233_fu_9883_p4;

assign zext_ln708_12_fu_3973_p1 = tmp_11_fu_3963_p4;

assign zext_ln708_130_fu_9908_p1 = tmp_234_fu_9898_p4;

assign zext_ln708_131_fu_10518_p1 = trunc_ln708_8_fu_10514_p1;

assign zext_ln708_132_fu_10533_p1 = tmp_251_fu_10523_p4;

assign zext_ln708_133_fu_10548_p1 = tmp_252_fu_10538_p4;

assign zext_ln708_134_fu_10563_p1 = tmp_253_fu_10553_p4;

assign zext_ln708_135_fu_10578_p1 = tmp_254_fu_10568_p4;

assign zext_ln708_136_fu_10593_p1 = tmp_255_fu_10583_p4;

assign zext_ln708_137_fu_10608_p1 = tmp_256_fu_10598_p4;

assign zext_ln708_138_fu_10623_p1 = tmp_257_fu_10613_p4;

assign zext_ln708_139_fu_10638_p1 = tmp_258_fu_10628_p4;

assign zext_ln708_13_fu_3988_p1 = tmp_12_fu_3978_p4;

assign zext_ln708_140_fu_10653_p1 = tmp_259_fu_10643_p4;

assign zext_ln708_141_fu_10668_p1 = tmp_260_fu_10658_p4;

assign zext_ln708_142_fu_10683_p1 = tmp_261_fu_10673_p4;

assign zext_ln708_143_fu_10698_p1 = tmp_262_fu_10688_p4;

assign zext_ln708_144_fu_10713_p1 = tmp_263_fu_10703_p4;

assign zext_ln708_145_fu_10728_p1 = tmp_264_fu_10718_p4;

assign zext_ln708_146_fu_10743_p1 = tmp_265_fu_10733_p4;

assign zext_ln708_147_fu_11353_p1 = trunc_ln708_9_fu_11349_p1;

assign zext_ln708_148_fu_11368_p1 = tmp_282_fu_11358_p4;

assign zext_ln708_149_fu_11383_p1 = tmp_283_fu_11373_p4;

assign zext_ln708_14_fu_4003_p1 = tmp_13_fu_3993_p4;

assign zext_ln708_150_fu_11398_p1 = tmp_284_fu_11388_p4;

assign zext_ln708_151_fu_11413_p1 = tmp_285_fu_11403_p4;

assign zext_ln708_152_fu_11428_p1 = tmp_286_fu_11418_p4;

assign zext_ln708_153_fu_11443_p1 = tmp_287_fu_11433_p4;

assign zext_ln708_154_fu_11458_p1 = tmp_288_fu_11448_p4;

assign zext_ln708_155_fu_11473_p1 = tmp_289_fu_11463_p4;

assign zext_ln708_156_fu_11488_p1 = tmp_290_fu_11478_p4;

assign zext_ln708_157_fu_11503_p1 = tmp_291_fu_11493_p4;

assign zext_ln708_158_fu_11518_p1 = tmp_292_fu_11508_p4;

assign zext_ln708_159_fu_11533_p1 = tmp_293_fu_11523_p4;

assign zext_ln708_15_fu_4018_p1 = tmp_14_fu_4008_p4;

assign zext_ln708_160_fu_11548_p1 = tmp_294_fu_11538_p4;

assign zext_ln708_161_fu_11563_p1 = tmp_295_fu_11553_p4;

assign zext_ln708_162_fu_11578_p1 = tmp_296_fu_11568_p4;

assign zext_ln708_16_fu_4033_p1 = tmp_15_fu_4023_p4;

assign zext_ln708_17_fu_4048_p1 = tmp_16_fu_4038_p4;

assign zext_ln708_18_fu_4063_p1 = tmp_17_fu_4053_p4;

assign zext_ln708_19_fu_4673_p1 = trunc_ln708_1_fu_4669_p1;

assign zext_ln708_20_fu_4688_p1 = tmp_34_fu_4678_p4;

assign zext_ln708_21_fu_4703_p1 = tmp_35_fu_4693_p4;

assign zext_ln708_22_fu_4718_p1 = tmp_36_fu_4708_p4;

assign zext_ln708_23_fu_4733_p1 = tmp_37_fu_4723_p4;

assign zext_ln708_24_fu_4748_p1 = tmp_38_fu_4738_p4;

assign zext_ln708_25_fu_4763_p1 = tmp_39_fu_4753_p4;

assign zext_ln708_26_fu_4778_p1 = tmp_40_fu_4768_p4;

assign zext_ln708_27_fu_4793_p1 = tmp_41_fu_4783_p4;

assign zext_ln708_28_fu_4808_p1 = tmp_42_fu_4798_p4;

assign zext_ln708_29_fu_4823_p1 = tmp_43_fu_4813_p4;

assign zext_ln708_30_fu_4838_p1 = tmp_44_fu_4828_p4;

assign zext_ln708_31_fu_4853_p1 = tmp_45_fu_4843_p4;

assign zext_ln708_32_fu_4868_p1 = tmp_46_fu_4858_p4;

assign zext_ln708_33_fu_4883_p1 = tmp_47_fu_4873_p4;

assign zext_ln708_34_fu_4898_p1 = tmp_48_fu_4888_p4;

assign zext_ln708_35_fu_5508_p1 = trunc_ln708_2_fu_5504_p1;

assign zext_ln708_36_fu_5523_p1 = tmp_65_fu_5513_p4;

assign zext_ln708_37_fu_5538_p1 = tmp_66_fu_5528_p4;

assign zext_ln708_38_fu_5553_p1 = tmp_67_fu_5543_p4;

assign zext_ln708_39_fu_5568_p1 = tmp_68_fu_5558_p4;

assign zext_ln708_40_fu_5583_p1 = tmp_69_fu_5573_p4;

assign zext_ln708_41_fu_5598_p1 = tmp_70_fu_5588_p4;

assign zext_ln708_42_fu_5613_p1 = tmp_71_fu_5603_p4;

assign zext_ln708_43_fu_5628_p1 = tmp_72_fu_5618_p4;

assign zext_ln708_44_fu_5643_p1 = tmp_73_fu_5633_p4;

assign zext_ln708_45_fu_5658_p1 = tmp_74_fu_5648_p4;

assign zext_ln708_46_fu_5673_p1 = tmp_75_fu_5663_p4;

assign zext_ln708_47_fu_5688_p1 = tmp_76_fu_5678_p4;

assign zext_ln708_48_fu_5703_p1 = tmp_77_fu_5693_p4;

assign zext_ln708_49_fu_5718_p1 = tmp_78_fu_5708_p4;

assign zext_ln708_4_fu_3853_p1 = tmp_s_fu_3843_p4;

assign zext_ln708_50_fu_5733_p1 = tmp_79_fu_5723_p4;

assign zext_ln708_51_fu_6343_p1 = trunc_ln708_3_fu_6339_p1;

assign zext_ln708_52_fu_6358_p1 = tmp_96_fu_6348_p4;

assign zext_ln708_53_fu_6373_p1 = tmp_97_fu_6363_p4;

assign zext_ln708_54_fu_6388_p1 = tmp_98_fu_6378_p4;

assign zext_ln708_55_fu_6403_p1 = tmp_99_fu_6393_p4;

assign zext_ln708_56_fu_6418_p1 = tmp_100_fu_6408_p4;

assign zext_ln708_57_fu_6433_p1 = tmp_101_fu_6423_p4;

assign zext_ln708_58_fu_6448_p1 = tmp_102_fu_6438_p4;

assign zext_ln708_59_fu_6463_p1 = tmp_103_fu_6453_p4;

assign zext_ln708_5_fu_3868_p1 = tmp_4_fu_3858_p4;

assign zext_ln708_60_fu_6478_p1 = tmp_104_fu_6468_p4;

assign zext_ln708_61_fu_6493_p1 = tmp_105_fu_6483_p4;

assign zext_ln708_62_fu_6508_p1 = tmp_106_fu_6498_p4;

assign zext_ln708_63_fu_6523_p1 = tmp_107_fu_6513_p4;

assign zext_ln708_64_fu_6538_p1 = tmp_108_fu_6528_p4;

assign zext_ln708_65_fu_6553_p1 = tmp_109_fu_6543_p4;

assign zext_ln708_66_fu_6568_p1 = tmp_110_fu_6558_p4;

assign zext_ln708_67_fu_7178_p1 = trunc_ln708_4_fu_7174_p1;

assign zext_ln708_68_fu_7193_p1 = tmp_127_fu_7183_p4;

assign zext_ln708_69_fu_7208_p1 = tmp_128_fu_7198_p4;

assign zext_ln708_6_fu_3883_p1 = tmp_5_fu_3873_p4;

assign zext_ln708_70_fu_7223_p1 = tmp_129_fu_7213_p4;

assign zext_ln708_71_fu_7238_p1 = tmp_130_fu_7228_p4;

assign zext_ln708_72_fu_7253_p1 = tmp_131_fu_7243_p4;

assign zext_ln708_73_fu_7268_p1 = tmp_132_fu_7258_p4;

assign zext_ln708_74_fu_7283_p1 = tmp_133_fu_7273_p4;

assign zext_ln708_75_fu_7298_p1 = tmp_134_fu_7288_p4;

assign zext_ln708_76_fu_7313_p1 = tmp_135_fu_7303_p4;

assign zext_ln708_77_fu_7328_p1 = tmp_136_fu_7318_p4;

assign zext_ln708_78_fu_7343_p1 = tmp_137_fu_7333_p4;

assign zext_ln708_79_fu_7358_p1 = tmp_138_fu_7348_p4;

assign zext_ln708_7_fu_3898_p1 = tmp_6_fu_3888_p4;

assign zext_ln708_80_fu_7373_p1 = tmp_139_fu_7363_p4;

assign zext_ln708_81_fu_7388_p1 = tmp_140_fu_7378_p4;

assign zext_ln708_82_fu_7403_p1 = tmp_141_fu_7393_p4;

assign zext_ln708_83_fu_8013_p1 = trunc_ln708_5_fu_8009_p1;

assign zext_ln708_84_fu_8028_p1 = tmp_158_fu_8018_p4;

assign zext_ln708_85_fu_8043_p1 = tmp_159_fu_8033_p4;

assign zext_ln708_86_fu_8058_p1 = tmp_160_fu_8048_p4;

assign zext_ln708_87_fu_8073_p1 = tmp_161_fu_8063_p4;

assign zext_ln708_88_fu_8088_p1 = tmp_162_fu_8078_p4;

assign zext_ln708_89_fu_8103_p1 = tmp_163_fu_8093_p4;

assign zext_ln708_8_fu_3913_p1 = tmp_7_fu_3903_p4;

assign zext_ln708_90_fu_8118_p1 = tmp_164_fu_8108_p4;

assign zext_ln708_91_fu_8133_p1 = tmp_165_fu_8123_p4;

assign zext_ln708_92_fu_8148_p1 = tmp_166_fu_8138_p4;

assign zext_ln708_93_fu_8163_p1 = tmp_167_fu_8153_p4;

assign zext_ln708_94_fu_8178_p1 = tmp_168_fu_8168_p4;

assign zext_ln708_95_fu_8193_p1 = tmp_169_fu_8183_p4;

assign zext_ln708_96_fu_8208_p1 = tmp_170_fu_8198_p4;

assign zext_ln708_97_fu_8223_p1 = tmp_171_fu_8213_p4;

assign zext_ln708_98_fu_8238_p1 = tmp_172_fu_8228_p4;

assign zext_ln708_99_fu_8848_p1 = trunc_ln708_6_fu_8844_p1;

assign zext_ln708_9_fu_3928_p1 = tmp_8_fu_3918_p4;

assign zext_ln708_fu_3838_p1 = trunc_ln708_fu_3834_p1;

endmodule //testEnc_process_r
