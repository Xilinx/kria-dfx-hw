   
    parameter PROC_NUM = 33;
    parameter ST_IDLE = 2'b0;
    parameter ST_DL_DETECTED = 2'b1;
    parameter ST_DL_REPORT = 2'b10;
   

    reg find_df_deadlock = 0;
    reg [1:0] CS_fsm;
    reg [1:0] NS_fsm;
    reg [PROC_NUM - 1:0] dl_detect_reg;
    reg [PROC_NUM - 1:0] dl_done_reg;
    reg [PROC_NUM - 1:0] origin_reg;
    reg [PROC_NUM - 1:0] dl_in_vec_reg;
    integer i;
    integer fp;

    // FSM State machine
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            CS_fsm <= ST_IDLE;
        end
        else begin
            CS_fsm <= NS_fsm;
        end
    end
    always @ (CS_fsm or dl_in_vec or dl_detect_reg or dl_done_reg or dl_in_vec or origin_reg) begin
        NS_fsm = CS_fsm;
        case (CS_fsm)
            ST_IDLE : begin
                if (|dl_in_vec) begin
                    NS_fsm = ST_DL_DETECTED;
                end
            end
            ST_DL_DETECTED: begin
                // has unreported deadlock cycle
                if (dl_detect_reg != dl_done_reg) begin
                    NS_fsm = ST_DL_REPORT;
                end
            end
            ST_DL_REPORT: begin
                if (|(dl_in_vec & origin_reg)) begin
                    NS_fsm = ST_DL_DETECTED;
                end
            end
        endcase
    end

    // dl_detect_reg record the procs that first detect deadlock
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            dl_detect_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_IDLE) begin
                dl_detect_reg <= dl_in_vec;
            end
        end
    end

    // dl_detect_out keeps in high after deadlock detected
    assign dl_detect_out = |dl_detect_reg;

    // dl_done_reg record the cycles has been reported
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            dl_done_reg <= 'b0;
        end
        else begin
            if ((CS_fsm == ST_DL_REPORT) && (|(dl_in_vec & dl_detect_reg) == 'b1)) begin
                dl_done_reg <= dl_done_reg | dl_in_vec;
            end
        end
    end

    // clear token once a cycle is done
    assign token_clear = (CS_fsm == ST_DL_REPORT) ? ((|(dl_in_vec & origin_reg)) ? 'b1 : 'b0) : 'b0;

    // origin_reg record the current cycle start id
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            origin_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                origin_reg <= origin;
            end
        end
    end
   
    // origin will be valid for only one cycle
    always @ (CS_fsm or dl_detect_reg or dl_done_reg) begin
        if (CS_fsm == ST_DL_DETECTED) begin
            for (i = 0; i < PROC_NUM; i = i + 1) begin
                if (dl_detect_reg[i] & ~dl_done_reg[i] & ~(|origin)) begin
                    origin = 'b1 << i;
                end
            end
        end
        else begin
            origin = 'b0;
        end
    end
    
    // dl_in_vec_reg record the current cycle dl_in_vec
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            dl_in_vec_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                dl_in_vec_reg <= origin;
            end
            else if (CS_fsm == ST_DL_REPORT) begin
                dl_in_vec_reg <= dl_in_vec;
            end
        end
    end
    
    // get the first valid proc index in dl vector
    function integer proc_index(input [PROC_NUM - 1:0] dl_vec);
        begin
            proc_index = 0;
            for (i = 0; i < PROC_NUM; i = i + 1) begin
                if (dl_vec[i]) begin
                    proc_index = i;
                end
            end
        end
    endfunction

    // get the proc path based on dl vector
    function [1048:0] proc_path(input [PROC_NUM - 1:0] dl_vec);
        integer index;
        begin
            index = proc_index(dl_vec);
            case (index)
                0 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0";
                end
                1 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0";
                end
                2 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0";
                end
                3 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0";
                end
                4 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0";
                end
                5 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_pxl_width_1_U0";
                end
                6 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0";
                end
                7 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.addrbound_2_U0";
                end
                8 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split48_proc_U0";
                end
                9 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2AxiStream_1_U0";
                end
                10 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.AxiStream2MatStream_1_U0";
                end
                11 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit2022_proc_U0";
                end
                12 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0";
                end
                13 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0";
                end
                14 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0";
                end
                15 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_pxl_width_U0";
                end
                16 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split35_proc_U0";
                end
                17 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.addrbound_1_U0";
                end
                18 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split37_proc_U0";
                end
                19 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2AxiStream_U0";
                end
                20 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.AxiStream2MatStream_U0";
                end
                21 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.nv122bgr_0_6_9_2160_3840_1_1_U0";
                end
                22 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.resize_1_9_2160_3840_720_720_1_9_U0";
                end
                23 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.preProcess_9_9_720_720_1_8_8_8_4_8_8_U0";
                end
                24 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0";
                end
                25 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0";
                end
                26 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split2_proc_U0";
                end
                27 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.addrbound_U0";
                end
                28 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split24_proc_U0";
                end
                29 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0";
                end
                30 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0";
                end
                31 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.MatStream2AxiStream_U0";
                end
                32 : begin
                    proc_path = "pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.AxiStream2Axi_U0";
                end
                default : begin
                    proc_path = "unknown";
                end
            endcase
        end
    endfunction

    // print the headlines of deadlock detection
    task print_dl_head;
        begin
            $display("\n//////////////////////////////////////////////////////////////////////////////");
            $display("// ERROR!!! DEADLOCK DETECTED at %0t ns! SIMULATION WILL BE STOPPED! //", $time);
            $display("//////////////////////////////////////////////////////////////////////////////");
            fp = $fopen("deadlock_db.dat", "w");
        end
    endtask

    // print the start of a cycle
    task print_cycle_start(input reg [1048:0] proc_path, input integer cycle_id);
        begin
            $display("/////////////////////////");
            $display("// Dependence cycle %0d:", cycle_id);
            $display("// (1): Process: %0s", proc_path);
            $fdisplay(fp, "Dependence_Cycle_ID %0d", cycle_id);
            $fdisplay(fp, "Dependence_Process_ID 1");
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print the end of deadlock detection
    task print_dl_end(input integer num, input integer record_time);
        begin
            $display("////////////////////////////////////////////////////////////////////////");
            $display("// Totally %0d cycles detected!", num);
            $display("////////////////////////////////////////////////////////////////////////");
            $display("// ERROR!!! DEADLOCK DETECTED at %0t ns! SIMULATION WILL BE STOPPED! //", record_time);
            $display("//////////////////////////////////////////////////////////////////////////////");
            $fdisplay(fp, "Dependence_Cycle_Number %0d", num);
            $fclose(fp);
        end
    endtask

    // print one proc component in the cycle
    task print_cycle_proc_comp(input reg [1048:0] proc_path, input integer cycle_comp_id);
        begin
            $display("// (%0d): Process: %0s", cycle_comp_id, proc_path);
            $fdisplay(fp, "Dependence_Process_ID %0d", cycle_comp_id);
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print one channel component in the cycle
    task print_cycle_chan_comp(input [PROC_NUM - 1:0] dl_vec1, input [PROC_NUM - 1:0] dl_vec2);
        reg [1072:0] chan_path;
        integer index1;
        integer index2;
        begin
            index1 = proc_index(dl_vec1);
            index2 = proc_index(dl_vec2);
            case (index1)
                0 : begin
                    case(index2)
                    2: begin
                        if (~pp_pipeline_accel_entry33_U0.img_inp_y_out_blk_n) begin
                            if (~img_inp_y_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.img_inp_y_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.img_inp_y_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~img_inp_y_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.img_inp_y_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.img_inp_y_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~pp_pipeline_accel_entry33_U0.in_img_linestride_out_blk_n) begin
                            if (~in_img_linestride_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.in_img_linestride_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.in_img_linestride_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~in_img_linestride_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.in_img_linestride_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.in_img_linestride_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_pp_pipeline_accel_entry33_U0_ap_ready & pp_pipeline_accel_entry33_U0.ap_idle & ~ap_sync_Array2xfMat_64_0_2160_3840_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0'");
                        end
                    end
                    12: begin
                        if (~pp_pipeline_accel_entry33_U0.img_inp_uv_out_blk_n) begin
                            if (~img_inp_uv_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.img_inp_uv_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.img_inp_uv_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~img_inp_uv_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.img_inp_uv_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.img_inp_uv_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_pp_pipeline_accel_entry33_U0_ap_ready & pp_pipeline_accel_entry33_U0.ap_idle & ~ap_sync_Array2xfMat_64_6_1080_1920_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0'");
                        end
                    end
                    24: begin
                        if (~pp_pipeline_accel_entry33_U0.img_out_out_blk_n) begin
                            if (~img_out_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.img_out_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.img_out_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~img_out_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.img_out_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.img_out_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~pp_pipeline_accel_entry33_U0.out_img_linestride_out_blk_n) begin
                            if (~out_img_linestride_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.out_img_linestride_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.out_img_linestride_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~out_img_linestride_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.out_img_linestride_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.out_img_linestride_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_xfMat2Array_64_9_720_720_1_1_U0_U.if_full_n & pp_pipeline_accel_entry33_U0.ap_start & ~pp_pipeline_accel_entry33_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_xfMat2Array_64_9_720_720_1_1_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'pp_pipeline_accel_pp_pipeline_accel.start_for_xfMat2Array_64_9_720_720_1_1_U0_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0',");
                        end
                    end
                    23: begin
                        if (~pp_pipeline_accel_entry33_U0.params_out_blk_n) begin
                            if (~params_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.params_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.preProcess_9_9_720_720_1_8_8_8_4_8_8_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.params_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~params_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.params_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.preProcess_9_9_720_720_1_8_8_8_4_8_8_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.params_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_pp_pipeline_accel_entry33_U0_ap_ready & pp_pipeline_accel_entry33_U0.ap_idle & ~ap_sync_preProcess_9_9_720_720_1_8_8_8_4_8_8_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'pp_pipeline_accel_pp_pipeline_accel.preProcess_9_9_720_720_1_8_8_8_4_8_8_U0'");
                        end
                    end
                    1: begin
                        if (~pp_pipeline_accel_entry33_U0.in_img_width_out_blk_n) begin
                            if (~in_img_width_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.in_img_width_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.in_img_width_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~in_img_width_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.in_img_width_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.in_img_width_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~pp_pipeline_accel_entry33_U0.in_img_height_out_blk_n) begin
                            if (~in_img_height_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.in_img_height_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.in_img_height_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~in_img_height_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.in_img_height_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.in_img_height_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~pp_pipeline_accel_entry33_U0.out_img_width_out_blk_n) begin
                            if (~out_img_width_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.out_img_width_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.out_img_width_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~out_img_width_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.out_img_width_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.out_img_width_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~pp_pipeline_accel_entry33_U0.out_img_height_out_blk_n) begin
                            if (~out_img_height_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.out_img_height_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.out_img_height_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~out_img_height_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.out_img_height_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.out_img_height_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0_U.if_full_n & pp_pipeline_accel_entry33_U0.ap_start & ~pp_pipeline_accel_entry33_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'pp_pipeline_accel_pp_pipeline_accel.start_for_Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0',");
                        end
                    end
                    11: begin
                        if (~pp_pipeline_accel_entry33_U0.in_img_linestride_out1_blk_n) begin
                            if (~in_img_linestride_c36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.in_img_linestride_c36_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit2022_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.in_img_linestride_c36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~in_img_linestride_c36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.in_img_linestride_c36_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit2022_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.in_img_linestride_c36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit2022_proc_U0_U.if_full_n & pp_pipeline_accel_entry33_U0.ap_start & ~pp_pipeline_accel_entry33_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit2022_proc_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'pp_pipeline_accel_pp_pipeline_accel.start_for_Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit2022_proc_U0_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit2022_proc_U0',");
                        end
                    end
                    endcase
                end
                1 : begin
                    case(index2)
                    0: begin
                        if (~Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.in_img_height_blk_n) begin
                            if (~in_img_height_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.in_img_height_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.in_img_height_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~in_img_height_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.in_img_height_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.in_img_height_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.in_img_width_blk_n) begin
                            if (~in_img_width_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.in_img_width_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.in_img_width_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~in_img_width_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.in_img_width_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.in_img_width_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.out_img_height_blk_n) begin
                            if (~out_img_height_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.out_img_height_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.out_img_height_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~out_img_height_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.out_img_height_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.out_img_height_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.out_img_width_blk_n) begin
                            if (~out_img_width_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.out_img_width_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.out_img_width_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~out_img_width_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.out_img_width_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.out_img_width_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0_U.if_empty_n & Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.ap_idle & ~start_for_Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'pp_pipeline_accel_pp_pipeline_accel.start_for_Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0',");
                        end
                    end
                    2: begin
                        if (~Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.imgInput_y_rows_out_blk_n) begin
                            if (~imgInput_y_rows_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.imgInput_y_rows_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.imgInput_y_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgInput_y_rows_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.imgInput_y_rows_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.imgInput_y_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.imgInput_y_cols_out_blk_n) begin
                            if (~imgInput_y_cols_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.imgInput_y_cols_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.imgInput_y_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgInput_y_cols_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.imgInput_y_cols_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.imgInput_y_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    22: begin
                        if (~Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.rgb_mat_rows_out_blk_n) begin
                            if (~rgb_mat_rows_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.rgb_mat_rows_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.resize_1_9_2160_3840_720_720_1_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.rgb_mat_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rgb_mat_rows_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.rgb_mat_rows_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.resize_1_9_2160_3840_720_720_1_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.rgb_mat_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.rgb_mat_cols_out_blk_n) begin
                            if (~rgb_mat_cols_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.rgb_mat_cols_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.resize_1_9_2160_3840_720_720_1_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.rgb_mat_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rgb_mat_cols_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.rgb_mat_cols_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.resize_1_9_2160_3840_720_720_1_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.rgb_mat_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.resize_out_mat_rows_out_blk_n) begin
                            if (~resize_out_mat_rows_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_rows_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.resize_1_9_2160_3840_720_720_1_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~resize_out_mat_rows_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_rows_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.resize_1_9_2160_3840_720_720_1_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.resize_out_mat_cols_out_blk_n) begin
                            if (~resize_out_mat_cols_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_cols_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.resize_1_9_2160_3840_720_720_1_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~resize_out_mat_cols_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_cols_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.resize_1_9_2160_3840_720_720_1_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_resize_1_9_2160_3840_720_720_1_9_U0_U.if_full_n & Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.ap_start & ~Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.real_start & (trans_in_cnt_8 == trans_out_cnt_8) & ~start_for_resize_1_9_2160_3840_720_720_1_9_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'pp_pipeline_accel_pp_pipeline_accel.start_for_resize_1_9_2160_3840_720_720_1_9_U0_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.resize_1_9_2160_3840_720_720_1_9_U0',");
                        end
                    end
                    24: begin
                        if (~Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.out_mat_rows_out_blk_n) begin
                            if (~out_mat_rows_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.out_mat_rows_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.out_mat_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~out_mat_rows_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.out_mat_rows_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.out_mat_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.out_mat_cols_out_blk_n) begin
                            if (~out_mat_cols_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.out_mat_cols_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.out_mat_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~out_mat_cols_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.out_mat_cols_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.out_mat_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                2 : begin
                    case(index2)
                    21: begin
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.AxiStream2MatStream_1_U0.imgInput_y_466_blk_n) begin
                            if (~imgInput_y_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.imgInput_y_data_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.nv122bgr_0_6_9_2160_3840_1_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.imgInput_y_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgInput_y_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.imgInput_y_data_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.nv122bgr_0_6_9_2160_3840_1_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.imgInput_y_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_0_2160_3840_1_U0.dstMat_1_out_blk_n) begin
                            if (~imgInput_y_rows_c37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.imgInput_y_rows_c37_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.nv122bgr_0_6_9_2160_3840_1_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.imgInput_y_rows_c37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgInput_y_rows_c37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.imgInput_y_rows_c37_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.nv122bgr_0_6_9_2160_3840_1_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.imgInput_y_rows_c37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_0_2160_3840_1_U0.dstMat_2_out_blk_n) begin
                            if (~imgInput_y_cols_c38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.imgInput_y_cols_c38_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.nv122bgr_0_6_9_2160_3840_1_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.imgInput_y_cols_c38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgInput_y_cols_c38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.imgInput_y_cols_c38_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.nv122bgr_0_6_9_2160_3840_1_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.imgInput_y_cols_c38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_nv122bgr_0_6_9_2160_3840_1_1_U0_U.if_full_n & Array2xfMat_64_0_2160_3840_1_U0.ap_start & ~Array2xfMat_64_0_2160_3840_1_U0.real_start & (trans_in_cnt_7 == trans_out_cnt_7) & ~start_for_nv122bgr_0_6_9_2160_3840_1_1_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'pp_pipeline_accel_pp_pipeline_accel.start_for_nv122bgr_0_6_9_2160_3840_1_1_U0_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.nv122bgr_0_6_9_2160_3840_1_1_U0',");
                        end
                    end
                    0: begin
                        if (~Array2xfMat_64_0_2160_3840_1_U0.srcPtr_blk_n) begin
                            if (~img_inp_y_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.img_inp_y_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.img_inp_y_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~img_inp_y_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.img_inp_y_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.img_inp_y_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_0_2160_3840_1_U0.stride_blk_n) begin
                            if (~in_img_linestride_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.in_img_linestride_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.in_img_linestride_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~in_img_linestride_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.in_img_linestride_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.in_img_linestride_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_Array2xfMat_64_0_2160_3840_1_U0_ap_ready & Array2xfMat_64_0_2160_3840_1_U0.ap_idle & ~ap_sync_pp_pipeline_accel_entry33_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0'");
                        end
                    end
                    1: begin
                        if (~Array2xfMat_64_0_2160_3840_1_U0.dstMat_1_blk_n) begin
                            if (~imgInput_y_rows_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.imgInput_y_rows_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.imgInput_y_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgInput_y_rows_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.imgInput_y_rows_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.imgInput_y_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_0_2160_3840_1_U0.dstMat_2_blk_n) begin
                            if (~imgInput_y_cols_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.imgInput_y_cols_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.imgInput_y_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgInput_y_cols_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.imgInput_y_cols_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.imgInput_y_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    12: begin
                        if (ap_sync_Array2xfMat_64_0_2160_3840_1_U0_ap_ready & Array2xfMat_64_0_2160_3840_1_U0.ap_idle & ~ap_sync_Array2xfMat_64_6_1080_1920_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0'");
                        end
                    end
                    23: begin
                        if (ap_sync_Array2xfMat_64_0_2160_3840_1_U0_ap_ready & Array2xfMat_64_0_2160_3840_1_U0.ap_idle & ~ap_sync_preProcess_9_9_720_720_1_8_8_8_4_8_8_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'pp_pipeline_accel_pp_pipeline_accel.preProcess_9_9_720_720_1_8_8_8_4_8_8_U0'");
                        end
                    end
                    endcase
                end
                3 : begin
                    case(index2)
                    4: begin
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0.din_out_blk_n) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.din_c1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.din_c1_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.din_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.din_c1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.din_c1_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.din_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0.rows_out_blk_n) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c2_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c2_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0.cols_out_blk_n) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c3_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c3_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0.stride_out_blk_n) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c4_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c4_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_Axi2Mat_entry12_U0_U.if_full_n & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0.ap_start & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0.real_start & (trans_in_cnt_1 == trans_out_cnt_1) & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_Axi2Mat_entry12_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_Axi2Mat_entry12_U0_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0',");
                        end
                    end
                    5: begin
                        if (Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ap_sync_Axi2Mat_1_entry3_U0_ap_ready & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0.ap_idle & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ap_sync_last_blk_pxl_width_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_pxl_width_1_U0'");
                        end
                    end
                    9: begin
                        if (Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ap_sync_Axi2Mat_1_entry3_U0_ap_ready & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0.ap_idle & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ap_sync_Axi2AxiStream_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2AxiStream_1_U0'");
                        end
                    end
                    endcase
                end
                4 : begin
                    case(index2)
                    3: begin
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0.din_blk_n) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.din_c1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.din_c1_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.din_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.din_c1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.din_c1_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.din_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0.rows_blk_n) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c2_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c2_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0.cols_blk_n) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c3_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c3_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0.stride_blk_n) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c4_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c4_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_Axi2Mat_entry12_U0_U.if_empty_n & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0.ap_idle & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_Axi2Mat_entry12_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_Axi2Mat_entry12_U0_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0',");
                        end
                    end
                    9: begin
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0.din_out_blk_n) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.din_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.din_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2AxiStream_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.din_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.din_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.din_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2AxiStream_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.din_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    6: begin
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0.rows_out_blk_n) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0.cols_out_blk_n) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0.stride_out_blk_n) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_Axi2Mat_Block_split46_proc_U0_U.if_full_n & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0.ap_start & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0.real_start & (trans_in_cnt_2 == trans_out_cnt_2) & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_Axi2Mat_Block_split46_proc_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_Axi2Mat_Block_split46_proc_U0_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0',");
                        end
                    end
                    endcase
                end
                5 : begin
                    case(index2)
                    10: begin
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_pxl_width_1_U0.ret_out_blk_n) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_width_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_width_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.AxiStream2MatStream_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_width_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_width_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_width_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.AxiStream2MatStream_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_width_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_AxiStream2MatStream_1_U0_U.if_full_n & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_pxl_width_1_U0.ap_start & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_pxl_width_1_U0.real_start & (trans_in_cnt_3 == trans_out_cnt_3) & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_AxiStream2MatStream_1_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_AxiStream2MatStream_1_U0_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.AxiStream2MatStream_1_U0',");
                        end
                    end
                    3: begin
                        if (Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ap_sync_last_blk_pxl_width_1_U0_ap_ready & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_pxl_width_1_U0.ap_idle & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ap_sync_Axi2Mat_1_entry3_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0'");
                        end
                    end
                    9: begin
                        if (Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ap_sync_last_blk_pxl_width_1_U0_ap_ready & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_pxl_width_1_U0.ap_idle & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ap_sync_Axi2AxiStream_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2AxiStream_1_U0'");
                        end
                    end
                    endcase
                end
                6 : begin
                    case(index2)
                    4: begin
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0.stride_blk_n) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0.cols_blk_n) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0.rows_blk_n) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_Axi2Mat_Block_split46_proc_U0_U.if_empty_n & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0.ap_idle & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_Axi2Mat_Block_split46_proc_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_Axi2Mat_Block_split46_proc_U0_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0',");
                        end
                    end
                    10: begin
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0.stride_out_blk_n) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c17_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.AxiStream2MatStream_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c17_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.AxiStream2MatStream_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0.cols_out_blk_n) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c18_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.AxiStream2MatStream_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c18_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.AxiStream2MatStream_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0.rows_out_blk_n) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c19_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.AxiStream2MatStream_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c19_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.AxiStream2MatStream_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                7 : begin
                    case(index2)
                    6: begin
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_cast_loc_channel_U.if_empty_n & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.addrbound_2_U0.ap_idle & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_cast_loc_channel_U.if_write) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_cast_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_cast_loc_channel_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_cast_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_cast_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_cast_loc_channel_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_cast_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_tmp_loc_channel_U.if_empty_n & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.addrbound_2_U0.ap_idle & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_tmp_loc_channel_U.if_write) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_tmp_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_tmp_loc_channel_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_tmp_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_tmp_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_tmp_loc_channel_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_tmp_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                8 : begin
                    case(index2)
                    7: begin
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.p_channel_U.if_empty_n & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split48_proc_U0.ap_idle & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.p_channel_U.if_write) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.p_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.p_channel_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.addrbound_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.p_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.p_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.p_channel_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.addrbound_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.p_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                9 : begin
                    case(index2)
                    10: begin
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2AxiStream_1_U0.ldata1_blk_n) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ldata_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ldata_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.AxiStream2MatStream_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ldata_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ldata_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ldata_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.AxiStream2MatStream_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ldata_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    4: begin
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2AxiStream_1_U0.din_blk_n) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.din_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.din_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.din_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.din_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.din_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.din_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    8: begin
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.axibound_V_U.if_empty_n & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2AxiStream_1_U0.ap_idle & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.axibound_V_U.if_write) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.axibound_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.axibound_V_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split48_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.axibound_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.axibound_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.axibound_V_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split48_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.axibound_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    3: begin
                        if (Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ap_sync_Axi2AxiStream_1_U0_ap_ready & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2AxiStream_1_U0.ap_idle & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ap_sync_Axi2Mat_1_entry3_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0'");
                        end
                    end
                    5: begin
                        if (Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ap_sync_Axi2AxiStream_1_U0_ap_ready & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2AxiStream_1_U0.ap_idle & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ap_sync_last_blk_pxl_width_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_pxl_width_1_U0'");
                        end
                    end
                    endcase
                end
                10 : begin
                    case(index2)
                    9: begin
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.AxiStream2MatStream_1_U0.ldata1_blk_n) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ldata_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ldata_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2AxiStream_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ldata_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ldata_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ldata_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2AxiStream_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ldata_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    6: begin
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.AxiStream2MatStream_1_U0.rows_blk_n) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c19_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c19_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c19_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c19_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_c19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.AxiStream2MatStream_1_U0.cols_bound_per_npc_blk_n) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c18_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c18_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_c18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.AxiStream2MatStream_1_U0.stride_blk_n) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c17_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c17_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.stride_c17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    5: begin
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.AxiStream2MatStream_1_U0.last_blk_width_blk_n) begin
                            if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_width_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_width_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_pxl_width_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_width_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_width_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_width_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_pxl_width_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_width_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_AxiStream2MatStream_1_U0_U.if_empty_n & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.AxiStream2MatStream_1_U0.ap_idle & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_AxiStream2MatStream_1_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_AxiStream2MatStream_1_U0_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_pxl_width_1_U0',");
                        end
                    end
                    endcase
                end
                11 : begin
                    case(index2)
                    0: begin
                        if (~Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit2022_proc_U0.in_img_linestride_blk_n) begin
                            if (~in_img_linestride_c36_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.in_img_linestride_c36_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.in_img_linestride_c36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~in_img_linestride_c36_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.in_img_linestride_c36_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.in_img_linestride_c36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit2022_proc_U0_U.if_empty_n & Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit2022_proc_U0.ap_idle & ~start_for_Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit2022_proc_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'pp_pipeline_accel_pp_pipeline_accel.start_for_Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit2022_proc_U0_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0',");
                        end
                    end
                    endcase
                end
                12 : begin
                    case(index2)
                    21: begin
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.AxiStream2MatStream_U0.imgInput_uv_467_blk_n) begin
                            if (~imgInput_uv_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.imgInput_uv_data_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.nv122bgr_0_6_9_2160_3840_1_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.imgInput_uv_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgInput_uv_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.imgInput_uv_data_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.nv122bgr_0_6_9_2160_3840_1_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.imgInput_uv_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin
                        if (~Array2xfMat_64_6_1080_1920_1_U0.img_inp_uv_blk_n) begin
                            if (~img_inp_uv_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.img_inp_uv_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.img_inp_uv_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~img_inp_uv_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.img_inp_uv_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.img_inp_uv_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_Array2xfMat_64_6_1080_1920_1_U0_ap_ready & Array2xfMat_64_6_1080_1920_1_U0.ap_idle & ~ap_sync_pp_pipeline_accel_entry33_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0'");
                        end
                    end
                    1: begin
                        if (~imgInput_uv_rows_channel_U.if_empty_n & Array2xfMat_64_6_1080_1920_1_U0.ap_idle & ~imgInput_uv_rows_channel_U.if_write) begin
                            if (~imgInput_uv_rows_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.imgInput_uv_rows_channel_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.imgInput_uv_rows_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgInput_uv_rows_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.imgInput_uv_rows_channel_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.imgInput_uv_rows_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~imgInput_uv_cols_channel_U.if_empty_n & Array2xfMat_64_6_1080_1920_1_U0.ap_idle & ~imgInput_uv_cols_channel_U.if_write) begin
                            if (~imgInput_uv_cols_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.imgInput_uv_cols_channel_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.imgInput_uv_cols_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgInput_uv_cols_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.imgInput_uv_cols_channel_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.imgInput_uv_cols_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    11: begin
                        if (~select_ln59_loc_channel_U.if_empty_n & Array2xfMat_64_6_1080_1920_1_U0.ap_idle & ~select_ln59_loc_channel_U.if_write) begin
                            if (~select_ln59_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.select_ln59_loc_channel_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit2022_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.select_ln59_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~select_ln59_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.select_ln59_loc_channel_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit2022_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.select_ln59_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    2: begin
                        if (ap_sync_Array2xfMat_64_6_1080_1920_1_U0_ap_ready & Array2xfMat_64_6_1080_1920_1_U0.ap_idle & ~ap_sync_Array2xfMat_64_0_2160_3840_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0'");
                        end
                    end
                    23: begin
                        if (ap_sync_Array2xfMat_64_6_1080_1920_1_U0_ap_ready & Array2xfMat_64_6_1080_1920_1_U0.ap_idle & ~ap_sync_preProcess_9_9_720_720_1_8_8_8_4_8_8_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'pp_pipeline_accel_pp_pipeline_accel.preProcess_9_9_720_720_1_8_8_8_4_8_8_U0'");
                        end
                    end
                    endcase
                end
                13 : begin
                    case(index2)
                    14: begin
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0.din_out_blk_n) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.din_c1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.din_c1_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.din_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.din_c1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.din_c1_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.din_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0.rows_out_blk_n) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c2_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c2_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0.cols_out_blk_n) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c3_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c3_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0.stride_out_blk_n) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c4_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c4_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_Axi2Mat_entry18_U0_U.if_full_n & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0.ap_start & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0.real_start & (trans_in_cnt_4 == trans_out_cnt_4) & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_Axi2Mat_entry18_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_Axi2Mat_entry18_U0_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0',");
                        end
                    end
                    15: begin
                        if (Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ap_sync_Axi2Mat_entry6_U0_ap_ready & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0.ap_idle & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ap_sync_last_blk_pxl_width_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_pxl_width_U0'");
                        end
                    end
                    19: begin
                        if (Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ap_sync_Axi2Mat_entry6_U0_ap_ready & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0.ap_idle & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ap_sync_Axi2AxiStream_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2AxiStream_U0'");
                        end
                    end
                    endcase
                end
                14 : begin
                    case(index2)
                    13: begin
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0.din_blk_n) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.din_c1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.din_c1_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.din_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.din_c1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.din_c1_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.din_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0.rows_blk_n) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c2_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c2_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0.cols_blk_n) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c3_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c3_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0.stride_blk_n) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c4_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c4_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_Axi2Mat_entry18_U0_U.if_empty_n & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0.ap_idle & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_Axi2Mat_entry18_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_Axi2Mat_entry18_U0_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0',");
                        end
                    end
                    19: begin
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0.din_out_blk_n) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.din_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.din_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2AxiStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.din_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.din_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.din_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2AxiStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.din_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    17: begin
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0.rows_out_blk_n) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.addrbound_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.addrbound_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    16: begin
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0.cols_out_blk_n) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split35_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split35_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0.stride_out_blk_n) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split35_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split35_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_Axi2Mat_Block_split35_proc_U0_U.if_full_n & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0.ap_start & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0.real_start & (trans_in_cnt_5 == trans_out_cnt_5) & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_Axi2Mat_Block_split35_proc_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_Axi2Mat_Block_split35_proc_U0_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split35_proc_U0',");
                        end
                    end
                    endcase
                end
                15 : begin
                    case(index2)
                    20: begin
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_pxl_width_U0.ret_out_blk_n) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_width_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_width_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.AxiStream2MatStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_width_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_width_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_width_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.AxiStream2MatStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_width_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_AxiStream2MatStream_U0_U.if_full_n & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_pxl_width_U0.ap_start & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_pxl_width_U0.real_start & (trans_in_cnt_6 == trans_out_cnt_6) & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_AxiStream2MatStream_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_AxiStream2MatStream_U0_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.AxiStream2MatStream_U0',");
                        end
                    end
                    13: begin
                        if (Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ap_sync_last_blk_pxl_width_U0_ap_ready & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_pxl_width_U0.ap_idle & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ap_sync_Axi2Mat_entry6_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0'");
                        end
                    end
                    19: begin
                        if (Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ap_sync_last_blk_pxl_width_U0_ap_ready & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_pxl_width_U0.ap_idle & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ap_sync_Axi2AxiStream_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2AxiStream_U0'");
                        end
                    end
                    endcase
                end
                16 : begin
                    case(index2)
                    14: begin
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split35_proc_U0.stride_blk_n) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split35_proc_U0.cols_blk_n) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_Axi2Mat_Block_split35_proc_U0_U.if_empty_n & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split35_proc_U0.ap_idle & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_Axi2Mat_Block_split35_proc_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_Axi2Mat_Block_split35_proc_U0_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0',");
                        end
                    end
                    20: begin
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split35_proc_U0.stride_out_blk_n) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c16_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.AxiStream2MatStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c16_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.AxiStream2MatStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split35_proc_U0.cols_out_blk_n) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c17_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.AxiStream2MatStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c17_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.AxiStream2MatStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                17 : begin
                    case(index2)
                    14: begin
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.addrbound_1_U0.rows_blk_n) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    16: begin
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_tmp_loc_channel_U.if_empty_n & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.addrbound_1_U0.ap_idle & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_tmp_loc_channel_U.if_write) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_tmp_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_tmp_loc_channel_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split35_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_tmp_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_tmp_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_tmp_loc_channel_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split35_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_tmp_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    20: begin
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.addrbound_1_U0.rows_out_blk_n) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c18_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.AxiStream2MatStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c18_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.AxiStream2MatStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                18 : begin
                    case(index2)
                    17: begin
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.p_channel_U.if_empty_n & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split37_proc_U0.ap_idle & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.p_channel_U.if_write) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.p_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.p_channel_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.addrbound_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.p_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.p_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.p_channel_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.addrbound_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.p_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                19 : begin
                    case(index2)
                    20: begin
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2AxiStream_U0.ldata1_blk_n) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ldata_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ldata_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.AxiStream2MatStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ldata_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ldata_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ldata_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.AxiStream2MatStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ldata_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    14: begin
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2AxiStream_U0.din_blk_n) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.din_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.din_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.din_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.din_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.din_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.din_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    18: begin
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.axibound_V_U.if_empty_n & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2AxiStream_U0.ap_idle & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.axibound_V_U.if_write) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.axibound_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.axibound_V_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split37_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.axibound_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.axibound_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.axibound_V_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split37_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.axibound_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    13: begin
                        if (Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ap_sync_Axi2AxiStream_U0_ap_ready & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2AxiStream_U0.ap_idle & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ap_sync_Axi2Mat_entry6_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0'");
                        end
                    end
                    15: begin
                        if (Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ap_sync_Axi2AxiStream_U0_ap_ready & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2AxiStream_U0.ap_idle & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ap_sync_last_blk_pxl_width_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_pxl_width_U0'");
                        end
                    end
                    endcase
                end
                20 : begin
                    case(index2)
                    19: begin
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.AxiStream2MatStream_U0.ldata1_blk_n) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ldata_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ldata_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2AxiStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ldata_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ldata_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ldata_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2AxiStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ldata_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    17: begin
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.AxiStream2MatStream_U0.rows_blk_n) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c18_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c18_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.addrbound_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c18_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c18_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.addrbound_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.rows_c18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    16: begin
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.AxiStream2MatStream_U0.cols_bound_per_npc_blk_n) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c17_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c17_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split35_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c17_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c17_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split35_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_c17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.AxiStream2MatStream_U0.stride_blk_n) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c16_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c16_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split35_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c16_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c16_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split35_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.stride_c16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    15: begin
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.AxiStream2MatStream_U0.last_blk_width_blk_n) begin
                            if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_width_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_width_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_pxl_width_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_width_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_width_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_width_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_pxl_width_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_width_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_AxiStream2MatStream_U0_U.if_empty_n & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.AxiStream2MatStream_U0.ap_idle & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_AxiStream2MatStream_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_AxiStream2MatStream_U0_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_pxl_width_U0',");
                        end
                    end
                    endcase
                end
                21 : begin
                    case(index2)
                    2: begin
                        if (~nv122bgr_0_6_9_2160_3840_1_1_U0.grp_KernNv122bgr_0_6_9_2160_3840_1_1_1_5_9_s_fu_44.imgInput_y_466_blk_n) begin
                            if (~imgInput_y_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.imgInput_y_data_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.imgInput_y_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgInput_y_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.imgInput_y_data_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.imgInput_y_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~nv122bgr_0_6_9_2160_3840_1_1_U0.src_y_rows_blk_n) begin
                            if (~imgInput_y_rows_c37_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.imgInput_y_rows_c37_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.imgInput_y_rows_c37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgInput_y_rows_c37_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.imgInput_y_rows_c37_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.imgInput_y_rows_c37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~nv122bgr_0_6_9_2160_3840_1_1_U0.src_y_cols_blk_n) begin
                            if (~imgInput_y_cols_c38_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.imgInput_y_cols_c38_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.imgInput_y_cols_c38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgInput_y_cols_c38_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.imgInput_y_cols_c38_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.imgInput_y_cols_c38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_nv122bgr_0_6_9_2160_3840_1_1_U0_U.if_empty_n & nv122bgr_0_6_9_2160_3840_1_1_U0.ap_idle & ~start_for_nv122bgr_0_6_9_2160_3840_1_1_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'pp_pipeline_accel_pp_pipeline_accel.start_for_nv122bgr_0_6_9_2160_3840_1_1_U0_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0',");
                        end
                    end
                    12: begin
                        if (~nv122bgr_0_6_9_2160_3840_1_1_U0.grp_KernNv122bgr_0_6_9_2160_3840_1_1_1_5_9_s_fu_44.imgInput_uv_467_blk_n) begin
                            if (~imgInput_uv_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.imgInput_uv_data_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.imgInput_uv_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~imgInput_uv_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.imgInput_uv_data_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.imgInput_uv_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    22: begin
                        if (~nv122bgr_0_6_9_2160_3840_1_1_U0.grp_KernNv122bgr_0_6_9_2160_3840_1_1_1_5_9_s_fu_44.rgb_mat_468_blk_n) begin
                            if (~rgb_mat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.rgb_mat_data_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.resize_1_9_2160_3840_720_720_1_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.rgb_mat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rgb_mat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.rgb_mat_data_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.resize_1_9_2160_3840_720_720_1_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.rgb_mat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                22 : begin
                    case(index2)
                    21: begin
                        if (~resize_1_9_2160_3840_720_720_1_9_U0.grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_80.rgb_mat_468_blk_n) begin
                            if (~rgb_mat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.rgb_mat_data_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.nv122bgr_0_6_9_2160_3840_1_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.rgb_mat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rgb_mat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.rgb_mat_data_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.nv122bgr_0_6_9_2160_3840_1_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.rgb_mat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    23: begin
                        if (~resize_1_9_2160_3840_720_720_1_9_U0.grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_80.resize_out_mat_469_blk_n) begin
                            if (~resize_out_mat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_data_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.preProcess_9_9_720_720_1_8_8_8_4_8_8_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~resize_out_mat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_data_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.preProcess_9_9_720_720_1_8_8_8_4_8_8_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~resize_1_9_2160_3840_720_720_1_9_U0.p_dst_rows_out_blk_n) begin
                            if (~resize_out_mat_rows_c39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_rows_c39_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.preProcess_9_9_720_720_1_8_8_8_4_8_8_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_rows_c39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~resize_out_mat_rows_c39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_rows_c39_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.preProcess_9_9_720_720_1_8_8_8_4_8_8_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_rows_c39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~resize_1_9_2160_3840_720_720_1_9_U0.p_dst_cols_out_blk_n) begin
                            if (~resize_out_mat_cols_c40_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_cols_c40_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.preProcess_9_9_720_720_1_8_8_8_4_8_8_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_cols_c40_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~resize_out_mat_cols_c40_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_cols_c40_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.preProcess_9_9_720_720_1_8_8_8_4_8_8_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_cols_c40_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin
                        if (~resize_1_9_2160_3840_720_720_1_9_U0.p_src_rows_blk_n) begin
                            if (~rgb_mat_rows_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.rgb_mat_rows_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.rgb_mat_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rgb_mat_rows_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.rgb_mat_rows_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.rgb_mat_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~resize_1_9_2160_3840_720_720_1_9_U0.p_src_cols_blk_n) begin
                            if (~rgb_mat_cols_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.rgb_mat_cols_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.rgb_mat_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rgb_mat_cols_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.rgb_mat_cols_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.rgb_mat_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~resize_1_9_2160_3840_720_720_1_9_U0.p_dst_rows_blk_n) begin
                            if (~resize_out_mat_rows_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_rows_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~resize_out_mat_rows_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_rows_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~resize_1_9_2160_3840_720_720_1_9_U0.p_dst_cols_blk_n) begin
                            if (~resize_out_mat_cols_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_cols_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~resize_out_mat_cols_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_cols_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_resize_1_9_2160_3840_720_720_1_9_U0_U.if_empty_n & resize_1_9_2160_3840_720_720_1_9_U0.ap_idle & ~start_for_resize_1_9_2160_3840_720_720_1_9_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'pp_pipeline_accel_pp_pipeline_accel.start_for_resize_1_9_2160_3840_720_720_1_9_U0_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0',");
                        end
                    end
                    endcase
                end
                23 : begin
                    case(index2)
                    22: begin
                        if (~preProcess_9_9_720_720_1_8_8_8_4_8_8_U0.resize_out_mat_469_blk_n) begin
                            if (~resize_out_mat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_data_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.resize_1_9_2160_3840_720_720_1_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~resize_out_mat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_data_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.resize_1_9_2160_3840_720_720_1_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~preProcess_9_9_720_720_1_8_8_8_4_8_8_U0.in_mat_rows_blk_n) begin
                            if (~resize_out_mat_rows_c39_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_rows_c39_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.resize_1_9_2160_3840_720_720_1_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_rows_c39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~resize_out_mat_rows_c39_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_rows_c39_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.resize_1_9_2160_3840_720_720_1_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_rows_c39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~preProcess_9_9_720_720_1_8_8_8_4_8_8_U0.in_mat_cols_blk_n) begin
                            if (~resize_out_mat_cols_c40_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_cols_c40_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.resize_1_9_2160_3840_720_720_1_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_cols_c40_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~resize_out_mat_cols_c40_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_cols_c40_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.resize_1_9_2160_3840_720_720_1_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.resize_out_mat_cols_c40_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    24: begin
                        if (~preProcess_9_9_720_720_1_8_8_8_4_8_8_U0.out_mat_470_blk_n) begin
                            if (~out_mat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.out_mat_data_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.out_mat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~out_mat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.out_mat_data_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.out_mat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin
                        if (~preProcess_9_9_720_720_1_8_8_8_4_8_8_U0.params_blk_n) begin
                            if (~params_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.params_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.params_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~params_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.params_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.params_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_preProcess_9_9_720_720_1_8_8_8_4_8_8_U0_ap_ready & preProcess_9_9_720_720_1_8_8_8_4_8_8_U0.ap_idle & ~ap_sync_pp_pipeline_accel_entry33_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0'");
                        end
                    end
                    2: begin
                        if (ap_sync_preProcess_9_9_720_720_1_8_8_8_4_8_8_U0_ap_ready & preProcess_9_9_720_720_1_8_8_8_4_8_8_U0.ap_idle & ~ap_sync_Array2xfMat_64_0_2160_3840_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_0_2160_3840_1_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_preProcess_9_9_720_720_1_8_8_8_4_8_8_U0_ap_ready & preProcess_9_9_720_720_1_8_8_8_4_8_8_U0.ap_idle & ~ap_sync_Array2xfMat_64_6_1080_1920_1_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'pp_pipeline_accel_pp_pipeline_accel.Array2xfMat_64_6_1080_1920_1_U0'");
                        end
                    end
                    endcase
                end
                24 : begin
                    case(index2)
                    23: begin
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.MatStream2AxiStream_U0.out_mat_470_blk_n) begin
                            if (~out_mat_data_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.out_mat_data_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.preProcess_9_9_720_720_1_8_8_8_4_8_8_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.out_mat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~out_mat_data_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.out_mat_data_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.preProcess_9_9_720_720_1_8_8_8_4_8_8_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.out_mat_data_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin
                        if (~xfMat2Array_64_9_720_720_1_1_U0.srcMat_rows_blk_n) begin
                            if (~out_mat_rows_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.out_mat_rows_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.out_mat_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~out_mat_rows_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.out_mat_rows_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.out_mat_rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~xfMat2Array_64_9_720_720_1_1_U0.srcMat_cols_blk_n) begin
                            if (~out_mat_cols_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.out_mat_cols_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.out_mat_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~out_mat_cols_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.out_mat_cols_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.out_mat_cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin
                        if (~xfMat2Array_64_9_720_720_1_1_U0.dstPtr_blk_n) begin
                            if (~img_out_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.img_out_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.img_out_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~img_out_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.img_out_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.img_out_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~xfMat2Array_64_9_720_720_1_1_U0.stride_blk_n) begin
                            if (~out_img_linestride_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.out_img_linestride_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.out_img_linestride_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~out_img_linestride_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.out_img_linestride_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.out_img_linestride_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_xfMat2Array_64_9_720_720_1_1_U0_U.if_empty_n & xfMat2Array_64_9_720_720_1_1_U0.ap_idle & ~start_for_xfMat2Array_64_9_720_720_1_1_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'pp_pipeline_accel_pp_pipeline_accel.start_for_xfMat2Array_64_9_720_720_1_1_U0_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.pp_pipeline_accel_entry33_U0',");
                        end
                    end
                    endcase
                end
                25 : begin
                    case(index2)
                    32: begin
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0.dout_out_blk_n) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.dout_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.dout_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.AxiStream2Axi_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.dout_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.dout_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.dout_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.AxiStream2Axi_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.dout_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    26: begin
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0.rows_out_blk_n) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0.cols_out_blk_n) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0.stride_out_blk_n) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.start_for_Mat2Axi_Block_split2_proc_U0_U.if_full_n & xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0.ap_start & ~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0.real_start & (trans_in_cnt_9 == trans_out_cnt_9) & ~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.start_for_Mat2Axi_Block_split2_proc_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.start_for_Mat2Axi_Block_split2_proc_U0_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split2_proc_U0',");
                        end
                    end
                    30: begin
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0.rows_out1_blk_n) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c12_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c12_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0.cols_out2_blk_n) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c13_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c13_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0.stride_out3_blk_n) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c14_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c14_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    29: begin
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.start_for_Mat2AxiStream_U0_U.if_full_n & xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0.ap_start & ~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0.real_start & (trans_in_cnt_9 == trans_out_cnt_9) & ~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.start_for_Mat2AxiStream_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.start_for_Mat2AxiStream_U0_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0',");
                        end
                    end
                    endcase
                end
                26 : begin
                    case(index2)
                    25: begin
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split2_proc_U0.stride_blk_n) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split2_proc_U0.cols_blk_n) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split2_proc_U0.rows_blk_n) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.start_for_Mat2Axi_Block_split2_proc_U0_U.if_empty_n & xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split2_proc_U0.ap_idle & ~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.start_for_Mat2Axi_Block_split2_proc_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.start_for_Mat2Axi_Block_split2_proc_U0_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0',");
                        end
                    end
                    endcase
                end
                27 : begin
                    case(index2)
                    26: begin
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_cast_loc_channel_U.if_empty_n & xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.addrbound_U0.ap_idle & ~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_cast_loc_channel_U.if_write) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_cast_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_cast_loc_channel_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_cast_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_cast_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_cast_loc_channel_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_cast_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_tmp_loc_channel_U.if_empty_n & xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.addrbound_U0.ap_idle & ~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_tmp_loc_channel_U.if_write) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_tmp_loc_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_tmp_loc_channel_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_tmp_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_tmp_loc_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_tmp_loc_channel_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_tmp_loc_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                28 : begin
                    case(index2)
                    27: begin
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.p_channel_U.if_empty_n & xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split24_proc_U0.ap_idle & ~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.p_channel_U.if_write) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.p_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.p_channel_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.addrbound_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.p_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.p_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.p_channel_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.addrbound_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.p_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                29 : begin
                    case(index2)
                    32: begin
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.MatStream2AxiStream_U0.ldata1_blk_n) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.ldata_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.ldata_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.AxiStream2Axi_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.ldata_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.ldata_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.ldata_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.AxiStream2Axi_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.ldata_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    25: begin
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0.rows_blk_n) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c12_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c12_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0.cols_blk_n) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c13_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c13_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0.stride_blk_n) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c14_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c14_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.start_for_Mat2AxiStream_U0_U.if_empty_n & xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.ap_idle & ~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.start_for_Mat2AxiStream_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.start_for_Mat2AxiStream_U0_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0',");
                        end
                    end
                    endcase
                end
                30 : begin
                    case(index2)
                    25: begin
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0.rows_blk_n) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c12_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c12_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c12_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c12_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_c12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0.cols_blk_n) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c13_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c13_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c13_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c13_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_c13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0.stride_blk_n) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c14_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c14_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c14_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c14_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.stride_c14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    31: begin
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0.rows_out_blk_n) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.rows_c_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.rows_c_i_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.MatStream2AxiStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.rows_c_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.rows_c_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.rows_c_i_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.MatStream2AxiStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.rows_c_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0.cols_out_blk_n) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.cols_c_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.cols_c_i_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.MatStream2AxiStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.cols_c_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.cols_c_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.cols_c_i_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.MatStream2AxiStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.cols_c_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0.stride_out_blk_n) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.stride_c_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.stride_c_i_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.MatStream2AxiStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.stride_c_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.stride_c_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.stride_c_i_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.MatStream2AxiStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.stride_c_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                31 : begin
                    case(index2)
                    32: begin
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.MatStream2AxiStream_U0.ldata1_blk_n) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.ldata_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.ldata_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.AxiStream2Axi_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.ldata_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.ldata_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.ldata_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.AxiStream2Axi_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.ldata_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    30: begin
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.MatStream2AxiStream_U0.rows_blk_n) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.rows_c_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.rows_c_i_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.rows_c_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.rows_c_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.rows_c_i_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.rows_c_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.MatStream2AxiStream_U0.cols_bound_per_npc_blk_n) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.cols_c_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.cols_c_i_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.cols_c_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.cols_c_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.cols_c_i_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.cols_c_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.p_channel_U.if_empty_n & xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.MatStream2AxiStream_U0.ap_idle & ~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.p_channel_U.if_write) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.p_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.p_channel_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.p_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.p_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.p_channel_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.p_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.MatStream2AxiStream_U0.stride_blk_n) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.stride_c_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.stride_c_i_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.stride_c_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.stride_c_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.stride_c_i_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.stride_c_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                32 : begin
                    case(index2)
                    31: begin
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.AxiStream2Axi_U0.ldata1_blk_n) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.ldata_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.ldata_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.MatStream2AxiStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.ldata_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.ldata_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.ldata_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.MatStream2AxiStream_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.ldata_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    25: begin
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.AxiStream2Axi_U0.dout_blk_n) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.dout_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.dout_c_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.dout_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.dout_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.dout_c_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.dout_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    28: begin
                        if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.axibound_V_U.if_empty_n & xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.AxiStream2Axi_U0.ap_idle & ~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.axibound_V_U.if_write) begin
                            if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.axibound_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.axibound_V_U' written by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split24_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.axibound_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.axibound_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.axibound_V_U' read by process 'pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split24_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path pp_pipeline_accel_pp_pipeline_accel.xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.axibound_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
            endcase
        end
    endtask

    // report
    initial begin : report_deadlock
        integer cycle_id;
        integer cycle_comp_id;
        integer record_time;
        wait (reset == 1);
        cycle_id = 1;
        record_time = 0;
        while (1) begin
            @ (negedge clock);
            case (CS_fsm)
                ST_DL_DETECTED: begin
                    cycle_comp_id = 2;
                    if (dl_detect_reg != dl_done_reg) begin
                        if (dl_done_reg == 'b0) begin
                            print_dl_head;
                            record_time = $time;
                        end
                        print_cycle_start(proc_path(origin), cycle_id);
                        cycle_id = cycle_id + 1;
                    end
                    else begin
                        print_dl_end((cycle_id - 1),record_time);
                        find_df_deadlock = 1;
                        @(negedge clock);
                        $finish;
                    end
                end
                ST_DL_REPORT: begin
                    if ((|(dl_in_vec)) & ~(|(dl_in_vec & origin_reg))) begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                        print_cycle_proc_comp(proc_path(dl_in_vec), cycle_comp_id);
                        cycle_comp_id = cycle_comp_id + 1;
                    end
                    else begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                    end
                end
            endcase
        end
    end
 
