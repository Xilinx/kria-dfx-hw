// Copyright (C) 2022, Advanced Micro Devices, Inc. All rights reserved.
// SPDX-License-Identifier: MIT
// ==============================================================
// Version: 2022.1.0
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module testDec_process_r (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        p_read,
        p_read1,
        p_read2,
        p_read3,
        p_read4,
        p_read5,
        p_read6,
        p_read7,
        p_read8,
        p_read9,
        p_read10,
        p_read11,
        p_read12,
        ciphertext,
        ap_return
);

parameter    ap_ST_fsm_pp0_stage0 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [127:0] p_read;
input  [127:0] p_read1;
input  [127:0] p_read2;
input  [127:0] p_read3;
input  [127:0] p_read4;
input  [127:0] p_read5;
input  [127:0] p_read6;
input  [127:0] p_read7;
input  [127:0] p_read8;
input  [127:0] p_read9;
input  [127:0] p_read10;
input  [127:0] p_read11;
input  [127:0] p_read12;
input  [127:0] ciphertext;
output  [127:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;

(* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg    ap_enable_reg_pp0_iter5;
reg    ap_enable_reg_pp0_iter6;
reg    ap_enable_reg_pp0_iter7;
reg    ap_enable_reg_pp0_iter8;
reg    ap_enable_reg_pp0_iter9;
reg    ap_enable_reg_pp0_iter10;
reg    ap_enable_reg_pp0_iter11;
reg    ap_enable_reg_pp0_iter12;
reg    ap_enable_reg_pp0_iter13;
reg    ap_enable_reg_pp0_iter14;
reg    ap_enable_reg_pp0_iter15;
reg    ap_enable_reg_pp0_iter16;
reg    ap_enable_reg_pp0_iter17;
reg    ap_enable_reg_pp0_iter18;
reg    ap_enable_reg_pp0_iter19;
reg    ap_enable_reg_pp0_iter20;
reg    ap_enable_reg_pp0_iter21;
reg    ap_enable_reg_pp0_iter22;
reg    ap_enable_reg_pp0_iter23;
reg    ap_idle_pp0;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_state4_pp0_stage0_iter3;
wire    ap_block_state5_pp0_stage0_iter4;
wire    ap_block_state6_pp0_stage0_iter5;
wire    ap_block_state7_pp0_stage0_iter6;
wire    ap_block_state8_pp0_stage0_iter7;
wire    ap_block_state9_pp0_stage0_iter8;
wire    ap_block_state10_pp0_stage0_iter9;
wire    ap_block_state11_pp0_stage0_iter10;
wire    ap_block_state12_pp0_stage0_iter11;
wire    ap_block_state13_pp0_stage0_iter12;
wire    ap_block_state14_pp0_stage0_iter13;
wire    ap_block_state15_pp0_stage0_iter14;
wire    ap_block_state16_pp0_stage0_iter15;
wire    ap_block_state17_pp0_stage0_iter16;
wire    ap_block_state18_pp0_stage0_iter17;
wire    ap_block_state19_pp0_stage0_iter18;
wire    ap_block_state20_pp0_stage0_iter19;
wire    ap_block_state21_pp0_stage0_iter20;
wire    ap_block_state22_pp0_stage0_iter21;
wire    ap_block_state23_pp0_stage0_iter22;
wire    ap_block_state24_pp0_stage0_iter23;
wire    ap_block_pp0_stage0_subdone;
wire   [7:0] decipher_0_iibox_address0;
reg    decipher_0_iibox_ce0;
wire   [7:0] decipher_0_iibox_q0;
wire   [7:0] decipher_0_iibox_address1;
reg    decipher_0_iibox_ce1;
wire   [7:0] decipher_0_iibox_q1;
wire   [7:0] decipher_0_iibox_address2;
reg    decipher_0_iibox_ce2;
wire   [7:0] decipher_0_iibox_q2;
wire   [7:0] decipher_0_iibox_address3;
reg    decipher_0_iibox_ce3;
wire   [7:0] decipher_0_iibox_q3;
wire   [7:0] decipher_0_iibox_address4;
reg    decipher_0_iibox_ce4;
wire   [7:0] decipher_0_iibox_q4;
wire   [7:0] decipher_0_iibox_address5;
reg    decipher_0_iibox_ce5;
wire   [7:0] decipher_0_iibox_q5;
wire   [7:0] decipher_0_iibox_address6;
reg    decipher_0_iibox_ce6;
wire   [7:0] decipher_0_iibox_q6;
wire   [7:0] decipher_0_iibox_address7;
reg    decipher_0_iibox_ce7;
wire   [7:0] decipher_0_iibox_q7;
wire   [7:0] decipher_0_iibox_address8;
reg    decipher_0_iibox_ce8;
wire   [7:0] decipher_0_iibox_q8;
wire   [7:0] decipher_0_iibox_address9;
reg    decipher_0_iibox_ce9;
wire   [7:0] decipher_0_iibox_q9;
wire   [7:0] decipher_0_iibox_address10;
reg    decipher_0_iibox_ce10;
wire   [7:0] decipher_0_iibox_q10;
wire   [7:0] decipher_0_iibox_address11;
reg    decipher_0_iibox_ce11;
wire   [7:0] decipher_0_iibox_q11;
wire   [7:0] decipher_0_iibox_address12;
reg    decipher_0_iibox_ce12;
wire   [7:0] decipher_0_iibox_q12;
wire   [7:0] decipher_0_iibox_address13;
reg    decipher_0_iibox_ce13;
wire   [7:0] decipher_0_iibox_q13;
wire   [7:0] decipher_0_iibox_address14;
reg    decipher_0_iibox_ce14;
wire   [7:0] decipher_0_iibox_q14;
wire   [7:0] decipher_0_iibox_address15;
reg    decipher_0_iibox_ce15;
wire   [7:0] decipher_0_iibox_q15;
wire   [7:0] decipher_0_iibox_address16;
reg    decipher_0_iibox_ce16;
wire   [7:0] decipher_0_iibox_q16;
wire   [7:0] decipher_0_iibox_address17;
reg    decipher_0_iibox_ce17;
wire   [7:0] decipher_0_iibox_q17;
wire   [7:0] decipher_0_iibox_address18;
reg    decipher_0_iibox_ce18;
wire   [7:0] decipher_0_iibox_q18;
wire   [7:0] decipher_0_iibox_address19;
reg    decipher_0_iibox_ce19;
wire   [7:0] decipher_0_iibox_q19;
wire   [7:0] decipher_0_iibox_address20;
reg    decipher_0_iibox_ce20;
wire   [7:0] decipher_0_iibox_q20;
wire   [7:0] decipher_0_iibox_address21;
reg    decipher_0_iibox_ce21;
wire   [7:0] decipher_0_iibox_q21;
wire   [7:0] decipher_0_iibox_address22;
reg    decipher_0_iibox_ce22;
wire   [7:0] decipher_0_iibox_q22;
wire   [7:0] decipher_0_iibox_address23;
reg    decipher_0_iibox_ce23;
wire   [7:0] decipher_0_iibox_q23;
wire   [7:0] decipher_0_iibox_address24;
reg    decipher_0_iibox_ce24;
wire   [7:0] decipher_0_iibox_q24;
wire   [7:0] decipher_0_iibox_address25;
reg    decipher_0_iibox_ce25;
wire   [7:0] decipher_0_iibox_q25;
wire   [7:0] decipher_0_iibox_address26;
reg    decipher_0_iibox_ce26;
wire   [7:0] decipher_0_iibox_q26;
wire   [7:0] decipher_0_iibox_address27;
reg    decipher_0_iibox_ce27;
wire   [7:0] decipher_0_iibox_q27;
wire   [7:0] decipher_0_iibox_address28;
reg    decipher_0_iibox_ce28;
wire   [7:0] decipher_0_iibox_q28;
wire   [7:0] decipher_0_iibox_address29;
reg    decipher_0_iibox_ce29;
wire   [7:0] decipher_0_iibox_q29;
wire   [7:0] decipher_0_iibox_address30;
reg    decipher_0_iibox_ce30;
wire   [7:0] decipher_0_iibox_q30;
wire   [7:0] decipher_0_iibox_address31;
reg    decipher_0_iibox_ce31;
wire   [7:0] decipher_0_iibox_q31;
wire   [7:0] decipher_0_iibox_address32;
reg    decipher_0_iibox_ce32;
wire   [7:0] decipher_0_iibox_q32;
wire   [7:0] decipher_0_iibox_address33;
reg    decipher_0_iibox_ce33;
wire   [7:0] decipher_0_iibox_q33;
wire   [7:0] decipher_0_iibox_address34;
reg    decipher_0_iibox_ce34;
wire   [7:0] decipher_0_iibox_q34;
wire   [7:0] decipher_0_iibox_address35;
reg    decipher_0_iibox_ce35;
wire   [7:0] decipher_0_iibox_q35;
wire   [7:0] decipher_0_iibox_address36;
reg    decipher_0_iibox_ce36;
wire   [7:0] decipher_0_iibox_q36;
wire   [7:0] decipher_0_iibox_address37;
reg    decipher_0_iibox_ce37;
wire   [7:0] decipher_0_iibox_q37;
wire   [7:0] decipher_0_iibox_address38;
reg    decipher_0_iibox_ce38;
wire   [7:0] decipher_0_iibox_q38;
wire   [7:0] decipher_0_iibox_address39;
reg    decipher_0_iibox_ce39;
wire   [7:0] decipher_0_iibox_q39;
wire   [7:0] decipher_0_iibox_address40;
reg    decipher_0_iibox_ce40;
wire   [7:0] decipher_0_iibox_q40;
wire   [7:0] decipher_0_iibox_address41;
reg    decipher_0_iibox_ce41;
wire   [7:0] decipher_0_iibox_q41;
wire   [7:0] decipher_0_iibox_address42;
reg    decipher_0_iibox_ce42;
wire   [7:0] decipher_0_iibox_q42;
wire   [7:0] decipher_0_iibox_address43;
reg    decipher_0_iibox_ce43;
wire   [7:0] decipher_0_iibox_q43;
wire   [7:0] decipher_0_iibox_address44;
reg    decipher_0_iibox_ce44;
wire   [7:0] decipher_0_iibox_q44;
wire   [7:0] decipher_0_iibox_address45;
reg    decipher_0_iibox_ce45;
wire   [7:0] decipher_0_iibox_q45;
wire   [7:0] decipher_0_iibox_address46;
reg    decipher_0_iibox_ce46;
wire   [7:0] decipher_0_iibox_q46;
wire   [7:0] decipher_0_iibox_address47;
reg    decipher_0_iibox_ce47;
wire   [7:0] decipher_0_iibox_q47;
wire   [7:0] decipher_0_iibox_address48;
reg    decipher_0_iibox_ce48;
wire   [7:0] decipher_0_iibox_q48;
wire   [7:0] decipher_0_iibox_address49;
reg    decipher_0_iibox_ce49;
wire   [7:0] decipher_0_iibox_q49;
wire   [7:0] decipher_0_iibox_address50;
reg    decipher_0_iibox_ce50;
wire   [7:0] decipher_0_iibox_q50;
wire   [7:0] decipher_0_iibox_address51;
reg    decipher_0_iibox_ce51;
wire   [7:0] decipher_0_iibox_q51;
wire   [7:0] decipher_0_iibox_address52;
reg    decipher_0_iibox_ce52;
wire   [7:0] decipher_0_iibox_q52;
wire   [7:0] decipher_0_iibox_address53;
reg    decipher_0_iibox_ce53;
wire   [7:0] decipher_0_iibox_q53;
wire   [7:0] decipher_0_iibox_address54;
reg    decipher_0_iibox_ce54;
wire   [7:0] decipher_0_iibox_q54;
wire   [7:0] decipher_0_iibox_address55;
reg    decipher_0_iibox_ce55;
wire   [7:0] decipher_0_iibox_q55;
wire   [7:0] decipher_0_iibox_address56;
reg    decipher_0_iibox_ce56;
wire   [7:0] decipher_0_iibox_q56;
wire   [7:0] decipher_0_iibox_address57;
reg    decipher_0_iibox_ce57;
wire   [7:0] decipher_0_iibox_q57;
wire   [7:0] decipher_0_iibox_address58;
reg    decipher_0_iibox_ce58;
wire   [7:0] decipher_0_iibox_q58;
wire   [7:0] decipher_0_iibox_address59;
reg    decipher_0_iibox_ce59;
wire   [7:0] decipher_0_iibox_q59;
wire   [7:0] decipher_0_iibox_address60;
reg    decipher_0_iibox_ce60;
wire   [7:0] decipher_0_iibox_q60;
wire   [7:0] decipher_0_iibox_address61;
reg    decipher_0_iibox_ce61;
wire   [7:0] decipher_0_iibox_q61;
wire   [7:0] decipher_0_iibox_address62;
reg    decipher_0_iibox_ce62;
wire   [7:0] decipher_0_iibox_q62;
wire   [7:0] decipher_0_iibox_address63;
reg    decipher_0_iibox_ce63;
wire   [7:0] decipher_0_iibox_q63;
wire   [7:0] decipher_0_iibox_address64;
reg    decipher_0_iibox_ce64;
wire   [7:0] decipher_0_iibox_q64;
wire   [7:0] decipher_0_iibox_address65;
reg    decipher_0_iibox_ce65;
wire   [7:0] decipher_0_iibox_q65;
wire   [7:0] decipher_0_iibox_address66;
reg    decipher_0_iibox_ce66;
wire   [7:0] decipher_0_iibox_q66;
wire   [7:0] decipher_0_iibox_address67;
reg    decipher_0_iibox_ce67;
wire   [7:0] decipher_0_iibox_q67;
wire   [7:0] decipher_0_iibox_address68;
reg    decipher_0_iibox_ce68;
wire   [7:0] decipher_0_iibox_q68;
wire   [7:0] decipher_0_iibox_address69;
reg    decipher_0_iibox_ce69;
wire   [7:0] decipher_0_iibox_q69;
wire   [7:0] decipher_0_iibox_address70;
reg    decipher_0_iibox_ce70;
wire   [7:0] decipher_0_iibox_q70;
wire   [7:0] decipher_0_iibox_address71;
reg    decipher_0_iibox_ce71;
wire   [7:0] decipher_0_iibox_q71;
wire   [7:0] decipher_0_iibox_address72;
reg    decipher_0_iibox_ce72;
wire   [7:0] decipher_0_iibox_q72;
wire   [7:0] decipher_0_iibox_address73;
reg    decipher_0_iibox_ce73;
wire   [7:0] decipher_0_iibox_q73;
wire   [7:0] decipher_0_iibox_address74;
reg    decipher_0_iibox_ce74;
wire   [7:0] decipher_0_iibox_q74;
wire   [7:0] decipher_0_iibox_address75;
reg    decipher_0_iibox_ce75;
wire   [7:0] decipher_0_iibox_q75;
wire   [7:0] decipher_0_iibox_address76;
reg    decipher_0_iibox_ce76;
wire   [7:0] decipher_0_iibox_q76;
wire   [7:0] decipher_0_iibox_address77;
reg    decipher_0_iibox_ce77;
wire   [7:0] decipher_0_iibox_q77;
wire   [7:0] decipher_0_iibox_address78;
reg    decipher_0_iibox_ce78;
wire   [7:0] decipher_0_iibox_q78;
wire   [7:0] decipher_0_iibox_address79;
reg    decipher_0_iibox_ce79;
wire   [7:0] decipher_0_iibox_q79;
wire   [7:0] decipher_0_iibox_address80;
reg    decipher_0_iibox_ce80;
wire   [7:0] decipher_0_iibox_q80;
wire   [7:0] decipher_0_iibox_address81;
reg    decipher_0_iibox_ce81;
wire   [7:0] decipher_0_iibox_q81;
wire   [7:0] decipher_0_iibox_address82;
reg    decipher_0_iibox_ce82;
wire   [7:0] decipher_0_iibox_q82;
wire   [7:0] decipher_0_iibox_address83;
reg    decipher_0_iibox_ce83;
wire   [7:0] decipher_0_iibox_q83;
wire   [7:0] decipher_0_iibox_address84;
reg    decipher_0_iibox_ce84;
wire   [7:0] decipher_0_iibox_q84;
wire   [7:0] decipher_0_iibox_address85;
reg    decipher_0_iibox_ce85;
wire   [7:0] decipher_0_iibox_q85;
wire   [7:0] decipher_0_iibox_address86;
reg    decipher_0_iibox_ce86;
wire   [7:0] decipher_0_iibox_q86;
wire   [7:0] decipher_0_iibox_address87;
reg    decipher_0_iibox_ce87;
wire   [7:0] decipher_0_iibox_q87;
wire   [7:0] decipher_0_iibox_address88;
reg    decipher_0_iibox_ce88;
wire   [7:0] decipher_0_iibox_q88;
wire   [7:0] decipher_0_iibox_address89;
reg    decipher_0_iibox_ce89;
wire   [7:0] decipher_0_iibox_q89;
wire   [7:0] decipher_0_iibox_address90;
reg    decipher_0_iibox_ce90;
wire   [7:0] decipher_0_iibox_q90;
wire   [7:0] decipher_0_iibox_address91;
reg    decipher_0_iibox_ce91;
wire   [7:0] decipher_0_iibox_q91;
wire   [7:0] decipher_0_iibox_address92;
reg    decipher_0_iibox_ce92;
wire   [7:0] decipher_0_iibox_q92;
wire   [7:0] decipher_0_iibox_address93;
reg    decipher_0_iibox_ce93;
wire   [7:0] decipher_0_iibox_q93;
wire   [7:0] decipher_0_iibox_address94;
reg    decipher_0_iibox_ce94;
wire   [7:0] decipher_0_iibox_q94;
wire   [7:0] decipher_0_iibox_address95;
reg    decipher_0_iibox_ce95;
wire   [7:0] decipher_0_iibox_q95;
wire   [7:0] decipher_0_iibox_address96;
reg    decipher_0_iibox_ce96;
wire   [7:0] decipher_0_iibox_q96;
wire   [7:0] decipher_0_iibox_address97;
reg    decipher_0_iibox_ce97;
wire   [7:0] decipher_0_iibox_q97;
wire   [7:0] decipher_0_iibox_address98;
reg    decipher_0_iibox_ce98;
wire   [7:0] decipher_0_iibox_q98;
wire   [7:0] decipher_0_iibox_address99;
reg    decipher_0_iibox_ce99;
wire   [7:0] decipher_0_iibox_q99;
wire   [7:0] decipher_0_iibox_address100;
reg    decipher_0_iibox_ce100;
wire   [7:0] decipher_0_iibox_q100;
wire   [7:0] decipher_0_iibox_address101;
reg    decipher_0_iibox_ce101;
wire   [7:0] decipher_0_iibox_q101;
wire   [7:0] decipher_0_iibox_address102;
reg    decipher_0_iibox_ce102;
wire   [7:0] decipher_0_iibox_q102;
wire   [7:0] decipher_0_iibox_address103;
reg    decipher_0_iibox_ce103;
wire   [7:0] decipher_0_iibox_q103;
wire   [7:0] decipher_0_iibox_address104;
reg    decipher_0_iibox_ce104;
wire   [7:0] decipher_0_iibox_q104;
wire   [7:0] decipher_0_iibox_address105;
reg    decipher_0_iibox_ce105;
wire   [7:0] decipher_0_iibox_q105;
wire   [7:0] decipher_0_iibox_address106;
reg    decipher_0_iibox_ce106;
wire   [7:0] decipher_0_iibox_q106;
wire   [7:0] decipher_0_iibox_address107;
reg    decipher_0_iibox_ce107;
wire   [7:0] decipher_0_iibox_q107;
wire   [7:0] decipher_0_iibox_address108;
reg    decipher_0_iibox_ce108;
wire   [7:0] decipher_0_iibox_q108;
wire   [7:0] decipher_0_iibox_address109;
reg    decipher_0_iibox_ce109;
wire   [7:0] decipher_0_iibox_q109;
wire   [7:0] decipher_0_iibox_address110;
reg    decipher_0_iibox_ce110;
wire   [7:0] decipher_0_iibox_q110;
wire   [7:0] decipher_0_iibox_address111;
reg    decipher_0_iibox_ce111;
wire   [7:0] decipher_0_iibox_q111;
wire   [7:0] decipher_0_iibox_address112;
reg    decipher_0_iibox_ce112;
wire   [7:0] decipher_0_iibox_q112;
wire   [7:0] decipher_0_iibox_address113;
reg    decipher_0_iibox_ce113;
wire   [7:0] decipher_0_iibox_q113;
wire   [7:0] decipher_0_iibox_address114;
reg    decipher_0_iibox_ce114;
wire   [7:0] decipher_0_iibox_q114;
wire   [7:0] decipher_0_iibox_address115;
reg    decipher_0_iibox_ce115;
wire   [7:0] decipher_0_iibox_q115;
wire   [7:0] decipher_0_iibox_address116;
reg    decipher_0_iibox_ce116;
wire   [7:0] decipher_0_iibox_q116;
wire   [7:0] decipher_0_iibox_address117;
reg    decipher_0_iibox_ce117;
wire   [7:0] decipher_0_iibox_q117;
wire   [7:0] decipher_0_iibox_address118;
reg    decipher_0_iibox_ce118;
wire   [7:0] decipher_0_iibox_q118;
wire   [7:0] decipher_0_iibox_address119;
reg    decipher_0_iibox_ce119;
wire   [7:0] decipher_0_iibox_q119;
wire   [7:0] decipher_0_iibox_address120;
reg    decipher_0_iibox_ce120;
wire   [7:0] decipher_0_iibox_q120;
wire   [7:0] decipher_0_iibox_address121;
reg    decipher_0_iibox_ce121;
wire   [7:0] decipher_0_iibox_q121;
wire   [7:0] decipher_0_iibox_address122;
reg    decipher_0_iibox_ce122;
wire   [7:0] decipher_0_iibox_q122;
wire   [7:0] decipher_0_iibox_address123;
reg    decipher_0_iibox_ce123;
wire   [7:0] decipher_0_iibox_q123;
wire   [7:0] decipher_0_iibox_address124;
reg    decipher_0_iibox_ce124;
wire   [7:0] decipher_0_iibox_q124;
wire   [7:0] decipher_0_iibox_address125;
reg    decipher_0_iibox_ce125;
wire   [7:0] decipher_0_iibox_q125;
wire   [7:0] decipher_0_iibox_address126;
reg    decipher_0_iibox_ce126;
wire   [7:0] decipher_0_iibox_q126;
wire   [7:0] decipher_0_iibox_address127;
reg    decipher_0_iibox_ce127;
wire   [7:0] decipher_0_iibox_q127;
wire   [7:0] decipher_0_iibox_address128;
reg    decipher_0_iibox_ce128;
wire   [7:0] decipher_0_iibox_q128;
wire   [7:0] decipher_0_iibox_address129;
reg    decipher_0_iibox_ce129;
wire   [7:0] decipher_0_iibox_q129;
wire   [7:0] decipher_0_iibox_address130;
reg    decipher_0_iibox_ce130;
wire   [7:0] decipher_0_iibox_q130;
wire   [7:0] decipher_0_iibox_address131;
reg    decipher_0_iibox_ce131;
wire   [7:0] decipher_0_iibox_q131;
wire   [7:0] decipher_0_iibox_address132;
reg    decipher_0_iibox_ce132;
wire   [7:0] decipher_0_iibox_q132;
wire   [7:0] decipher_0_iibox_address133;
reg    decipher_0_iibox_ce133;
wire   [7:0] decipher_0_iibox_q133;
wire   [7:0] decipher_0_iibox_address134;
reg    decipher_0_iibox_ce134;
wire   [7:0] decipher_0_iibox_q134;
wire   [7:0] decipher_0_iibox_address135;
reg    decipher_0_iibox_ce135;
wire   [7:0] decipher_0_iibox_q135;
wire   [7:0] decipher_0_iibox_address136;
reg    decipher_0_iibox_ce136;
wire   [7:0] decipher_0_iibox_q136;
wire   [7:0] decipher_0_iibox_address137;
reg    decipher_0_iibox_ce137;
wire   [7:0] decipher_0_iibox_q137;
wire   [7:0] decipher_0_iibox_address138;
reg    decipher_0_iibox_ce138;
wire   [7:0] decipher_0_iibox_q138;
wire   [7:0] decipher_0_iibox_address139;
reg    decipher_0_iibox_ce139;
wire   [7:0] decipher_0_iibox_q139;
wire   [7:0] decipher_0_iibox_address140;
reg    decipher_0_iibox_ce140;
wire   [7:0] decipher_0_iibox_q140;
wire   [7:0] decipher_0_iibox_address141;
reg    decipher_0_iibox_ce141;
wire   [7:0] decipher_0_iibox_q141;
wire   [7:0] decipher_0_iibox_address142;
reg    decipher_0_iibox_ce142;
wire   [7:0] decipher_0_iibox_q142;
wire   [7:0] decipher_0_iibox_address143;
reg    decipher_0_iibox_ce143;
wire   [7:0] decipher_0_iibox_q143;
wire   [7:0] decipher_0_iibox_address144;
reg    decipher_0_iibox_ce144;
wire   [7:0] decipher_0_iibox_q144;
wire   [7:0] decipher_0_iibox_address145;
reg    decipher_0_iibox_ce145;
wire   [7:0] decipher_0_iibox_q145;
wire   [7:0] decipher_0_iibox_address146;
reg    decipher_0_iibox_ce146;
wire   [7:0] decipher_0_iibox_q146;
wire   [7:0] decipher_0_iibox_address147;
reg    decipher_0_iibox_ce147;
wire   [7:0] decipher_0_iibox_q147;
wire   [7:0] decipher_0_iibox_address148;
reg    decipher_0_iibox_ce148;
wire   [7:0] decipher_0_iibox_q148;
wire   [7:0] decipher_0_iibox_address149;
reg    decipher_0_iibox_ce149;
wire   [7:0] decipher_0_iibox_q149;
wire   [7:0] decipher_0_iibox_address150;
reg    decipher_0_iibox_ce150;
wire   [7:0] decipher_0_iibox_q150;
wire   [7:0] decipher_0_iibox_address151;
reg    decipher_0_iibox_ce151;
wire   [7:0] decipher_0_iibox_q151;
wire   [7:0] decipher_0_iibox_address152;
reg    decipher_0_iibox_ce152;
wire   [7:0] decipher_0_iibox_q152;
wire   [7:0] decipher_0_iibox_address153;
reg    decipher_0_iibox_ce153;
wire   [7:0] decipher_0_iibox_q153;
wire   [7:0] decipher_0_iibox_address154;
reg    decipher_0_iibox_ce154;
wire   [7:0] decipher_0_iibox_q154;
wire   [7:0] decipher_0_iibox_address155;
reg    decipher_0_iibox_ce155;
wire   [7:0] decipher_0_iibox_q155;
wire   [7:0] decipher_0_iibox_address156;
reg    decipher_0_iibox_ce156;
wire   [7:0] decipher_0_iibox_q156;
wire   [7:0] decipher_0_iibox_address157;
reg    decipher_0_iibox_ce157;
wire   [7:0] decipher_0_iibox_q157;
wire   [7:0] decipher_0_iibox_address158;
reg    decipher_0_iibox_ce158;
wire   [7:0] decipher_0_iibox_q158;
wire   [7:0] decipher_0_iibox_address159;
reg    decipher_0_iibox_ce159;
wire   [7:0] decipher_0_iibox_q159;
wire   [7:0] decipher_0_iibox_address160;
reg    decipher_0_iibox_ce160;
wire   [7:0] decipher_0_iibox_q160;
wire   [7:0] decipher_0_iibox_address161;
reg    decipher_0_iibox_ce161;
wire   [7:0] decipher_0_iibox_q161;
wire   [7:0] decipher_0_iibox_address162;
reg    decipher_0_iibox_ce162;
wire   [7:0] decipher_0_iibox_q162;
wire   [7:0] decipher_0_iibox_address163;
reg    decipher_0_iibox_ce163;
wire   [7:0] decipher_0_iibox_q163;
wire   [7:0] decipher_0_iibox_address164;
reg    decipher_0_iibox_ce164;
wire   [7:0] decipher_0_iibox_q164;
wire   [7:0] decipher_0_iibox_address165;
reg    decipher_0_iibox_ce165;
wire   [7:0] decipher_0_iibox_q165;
wire   [7:0] decipher_0_iibox_address166;
reg    decipher_0_iibox_ce166;
wire   [7:0] decipher_0_iibox_q166;
wire   [7:0] decipher_0_iibox_address167;
reg    decipher_0_iibox_ce167;
wire   [7:0] decipher_0_iibox_q167;
wire   [7:0] decipher_0_iibox_address168;
reg    decipher_0_iibox_ce168;
wire   [7:0] decipher_0_iibox_q168;
wire   [7:0] decipher_0_iibox_address169;
reg    decipher_0_iibox_ce169;
wire   [7:0] decipher_0_iibox_q169;
wire   [7:0] decipher_0_iibox_address170;
reg    decipher_0_iibox_ce170;
wire   [7:0] decipher_0_iibox_q170;
wire   [7:0] decipher_0_iibox_address171;
reg    decipher_0_iibox_ce171;
wire   [7:0] decipher_0_iibox_q171;
wire   [7:0] decipher_0_iibox_address172;
reg    decipher_0_iibox_ce172;
wire   [7:0] decipher_0_iibox_q172;
wire   [7:0] decipher_0_iibox_address173;
reg    decipher_0_iibox_ce173;
wire   [7:0] decipher_0_iibox_q173;
wire   [7:0] decipher_0_iibox_address174;
reg    decipher_0_iibox_ce174;
wire   [7:0] decipher_0_iibox_q174;
wire   [7:0] decipher_0_iibox_address175;
reg    decipher_0_iibox_ce175;
wire   [7:0] decipher_0_iibox_q175;
wire   [7:0] decipher_0_iibox_address176;
reg    decipher_0_iibox_ce176;
wire   [7:0] decipher_0_iibox_q176;
wire   [7:0] decipher_0_iibox_address177;
reg    decipher_0_iibox_ce177;
wire   [7:0] decipher_0_iibox_q177;
wire   [7:0] decipher_0_iibox_address178;
reg    decipher_0_iibox_ce178;
wire   [7:0] decipher_0_iibox_q178;
wire   [7:0] decipher_0_iibox_address179;
reg    decipher_0_iibox_ce179;
wire   [7:0] decipher_0_iibox_q179;
wire   [7:0] decipher_0_iibox_address180;
reg    decipher_0_iibox_ce180;
wire   [7:0] decipher_0_iibox_q180;
wire   [7:0] decipher_0_iibox_address181;
reg    decipher_0_iibox_ce181;
wire   [7:0] decipher_0_iibox_q181;
wire   [7:0] decipher_0_iibox_address182;
reg    decipher_0_iibox_ce182;
wire   [7:0] decipher_0_iibox_q182;
wire   [7:0] decipher_0_iibox_address183;
reg    decipher_0_iibox_ce183;
wire   [7:0] decipher_0_iibox_q183;
wire   [7:0] decipher_0_iibox_address184;
reg    decipher_0_iibox_ce184;
wire   [7:0] decipher_0_iibox_q184;
wire   [7:0] decipher_0_iibox_address185;
reg    decipher_0_iibox_ce185;
wire   [7:0] decipher_0_iibox_q185;
wire   [7:0] decipher_0_iibox_address186;
reg    decipher_0_iibox_ce186;
wire   [7:0] decipher_0_iibox_q186;
wire   [7:0] decipher_0_iibox_address187;
reg    decipher_0_iibox_ce187;
wire   [7:0] decipher_0_iibox_q187;
wire   [7:0] decipher_0_iibox_address188;
reg    decipher_0_iibox_ce188;
wire   [7:0] decipher_0_iibox_q188;
wire   [7:0] decipher_0_iibox_address189;
reg    decipher_0_iibox_ce189;
wire   [7:0] decipher_0_iibox_q189;
wire   [7:0] decipher_0_iibox_address190;
reg    decipher_0_iibox_ce190;
wire   [7:0] decipher_0_iibox_q190;
wire   [7:0] decipher_0_iibox_address191;
reg    decipher_0_iibox_ce191;
wire   [7:0] decipher_0_iibox_q191;
wire   [7:0] decipher_0_i32box_address0;
reg    decipher_0_i32box_ce0;
wire   [31:0] decipher_0_i32box_q0;
wire   [7:0] decipher_0_i32box_address1;
reg    decipher_0_i32box_ce1;
wire   [31:0] decipher_0_i32box_q1;
wire   [7:0] decipher_0_i32box_address2;
reg    decipher_0_i32box_ce2;
wire   [31:0] decipher_0_i32box_q2;
wire   [7:0] decipher_0_i32box_address3;
reg    decipher_0_i32box_ce3;
wire   [31:0] decipher_0_i32box_q3;
wire   [7:0] decipher_0_i32box_address4;
reg    decipher_0_i32box_ce4;
wire   [31:0] decipher_0_i32box_q4;
wire   [7:0] decipher_0_i32box_address5;
reg    decipher_0_i32box_ce5;
wire   [31:0] decipher_0_i32box_q5;
wire   [7:0] decipher_0_i32box_address6;
reg    decipher_0_i32box_ce6;
wire   [31:0] decipher_0_i32box_q6;
wire   [7:0] decipher_0_i32box_address7;
reg    decipher_0_i32box_ce7;
wire   [31:0] decipher_0_i32box_q7;
wire   [7:0] decipher_0_i32box_address8;
reg    decipher_0_i32box_ce8;
wire   [31:0] decipher_0_i32box_q8;
wire   [7:0] decipher_0_i32box_address9;
reg    decipher_0_i32box_ce9;
wire   [31:0] decipher_0_i32box_q9;
wire   [7:0] decipher_0_i32box_address10;
reg    decipher_0_i32box_ce10;
wire   [31:0] decipher_0_i32box_q10;
wire   [7:0] decipher_0_i32box_address11;
reg    decipher_0_i32box_ce11;
wire   [31:0] decipher_0_i32box_q11;
wire   [7:0] decipher_0_i32box_address12;
reg    decipher_0_i32box_ce12;
wire   [31:0] decipher_0_i32box_q12;
wire   [7:0] decipher_0_i32box_address13;
reg    decipher_0_i32box_ce13;
wire   [31:0] decipher_0_i32box_q13;
wire   [7:0] decipher_0_i32box_address14;
reg    decipher_0_i32box_ce14;
wire   [31:0] decipher_0_i32box_q14;
wire   [7:0] decipher_0_i32box_address15;
reg    decipher_0_i32box_ce15;
wire   [31:0] decipher_0_i32box_q15;
wire   [7:0] decipher_0_i32box_address16;
reg    decipher_0_i32box_ce16;
wire   [31:0] decipher_0_i32box_q16;
wire   [7:0] decipher_0_i32box_address17;
reg    decipher_0_i32box_ce17;
wire   [31:0] decipher_0_i32box_q17;
wire   [7:0] decipher_0_i32box_address18;
reg    decipher_0_i32box_ce18;
wire   [31:0] decipher_0_i32box_q18;
wire   [7:0] decipher_0_i32box_address19;
reg    decipher_0_i32box_ce19;
wire   [31:0] decipher_0_i32box_q19;
wire   [7:0] decipher_0_i32box_address20;
reg    decipher_0_i32box_ce20;
wire   [31:0] decipher_0_i32box_q20;
wire   [7:0] decipher_0_i32box_address21;
reg    decipher_0_i32box_ce21;
wire   [31:0] decipher_0_i32box_q21;
wire   [7:0] decipher_0_i32box_address22;
reg    decipher_0_i32box_ce22;
wire   [31:0] decipher_0_i32box_q22;
wire   [7:0] decipher_0_i32box_address23;
reg    decipher_0_i32box_ce23;
wire   [31:0] decipher_0_i32box_q23;
wire   [7:0] decipher_0_i32box_address24;
reg    decipher_0_i32box_ce24;
wire   [31:0] decipher_0_i32box_q24;
wire   [7:0] decipher_0_i32box_address25;
reg    decipher_0_i32box_ce25;
wire   [31:0] decipher_0_i32box_q25;
wire   [7:0] decipher_0_i32box_address26;
reg    decipher_0_i32box_ce26;
wire   [31:0] decipher_0_i32box_q26;
wire   [7:0] decipher_0_i32box_address27;
reg    decipher_0_i32box_ce27;
wire   [31:0] decipher_0_i32box_q27;
wire   [7:0] decipher_0_i32box_address28;
reg    decipher_0_i32box_ce28;
wire   [31:0] decipher_0_i32box_q28;
wire   [7:0] decipher_0_i32box_address29;
reg    decipher_0_i32box_ce29;
wire   [31:0] decipher_0_i32box_q29;
wire   [7:0] decipher_0_i32box_address30;
reg    decipher_0_i32box_ce30;
wire   [31:0] decipher_0_i32box_q30;
wire   [7:0] decipher_0_i32box_address31;
reg    decipher_0_i32box_ce31;
wire   [31:0] decipher_0_i32box_q31;
wire   [7:0] decipher_0_i32box_address32;
reg    decipher_0_i32box_ce32;
wire   [31:0] decipher_0_i32box_q32;
wire   [7:0] decipher_0_i32box_address33;
reg    decipher_0_i32box_ce33;
wire   [31:0] decipher_0_i32box_q33;
wire   [7:0] decipher_0_i32box_address34;
reg    decipher_0_i32box_ce34;
wire   [31:0] decipher_0_i32box_q34;
wire   [7:0] decipher_0_i32box_address35;
reg    decipher_0_i32box_ce35;
wire   [31:0] decipher_0_i32box_q35;
wire   [7:0] decipher_0_i32box_address36;
reg    decipher_0_i32box_ce36;
wire   [31:0] decipher_0_i32box_q36;
wire   [7:0] decipher_0_i32box_address37;
reg    decipher_0_i32box_ce37;
wire   [31:0] decipher_0_i32box_q37;
wire   [7:0] decipher_0_i32box_address38;
reg    decipher_0_i32box_ce38;
wire   [31:0] decipher_0_i32box_q38;
wire   [7:0] decipher_0_i32box_address39;
reg    decipher_0_i32box_ce39;
wire   [31:0] decipher_0_i32box_q39;
wire   [7:0] decipher_0_i32box_address40;
reg    decipher_0_i32box_ce40;
wire   [31:0] decipher_0_i32box_q40;
wire   [7:0] decipher_0_i32box_address41;
reg    decipher_0_i32box_ce41;
wire   [31:0] decipher_0_i32box_q41;
wire   [7:0] decipher_0_i32box_address42;
reg    decipher_0_i32box_ce42;
wire   [31:0] decipher_0_i32box_q42;
wire   [7:0] decipher_0_i32box_address43;
reg    decipher_0_i32box_ce43;
wire   [31:0] decipher_0_i32box_q43;
wire   [7:0] decipher_0_i32box_address44;
reg    decipher_0_i32box_ce44;
wire   [31:0] decipher_0_i32box_q44;
wire   [7:0] decipher_0_i32box_address45;
reg    decipher_0_i32box_ce45;
wire   [31:0] decipher_0_i32box_q45;
wire   [7:0] decipher_0_i32box_address46;
reg    decipher_0_i32box_ce46;
wire   [31:0] decipher_0_i32box_q46;
wire   [7:0] decipher_0_i32box_address47;
reg    decipher_0_i32box_ce47;
wire   [31:0] decipher_0_i32box_q47;
wire   [7:0] decipher_0_i32box_address48;
reg    decipher_0_i32box_ce48;
wire   [31:0] decipher_0_i32box_q48;
wire   [7:0] decipher_0_i32box_address49;
reg    decipher_0_i32box_ce49;
wire   [31:0] decipher_0_i32box_q49;
wire   [7:0] decipher_0_i32box_address50;
reg    decipher_0_i32box_ce50;
wire   [31:0] decipher_0_i32box_q50;
wire   [7:0] decipher_0_i32box_address51;
reg    decipher_0_i32box_ce51;
wire   [31:0] decipher_0_i32box_q51;
wire   [7:0] decipher_0_i32box_address52;
reg    decipher_0_i32box_ce52;
wire   [31:0] decipher_0_i32box_q52;
wire   [7:0] decipher_0_i32box_address53;
reg    decipher_0_i32box_ce53;
wire   [31:0] decipher_0_i32box_q53;
wire   [7:0] decipher_0_i32box_address54;
reg    decipher_0_i32box_ce54;
wire   [31:0] decipher_0_i32box_q54;
wire   [7:0] decipher_0_i32box_address55;
reg    decipher_0_i32box_ce55;
wire   [31:0] decipher_0_i32box_q55;
wire   [7:0] decipher_0_i32box_address56;
reg    decipher_0_i32box_ce56;
wire   [31:0] decipher_0_i32box_q56;
wire   [7:0] decipher_0_i32box_address57;
reg    decipher_0_i32box_ce57;
wire   [31:0] decipher_0_i32box_q57;
wire   [7:0] decipher_0_i32box_address58;
reg    decipher_0_i32box_ce58;
wire   [31:0] decipher_0_i32box_q58;
wire   [7:0] decipher_0_i32box_address59;
reg    decipher_0_i32box_ce59;
wire   [31:0] decipher_0_i32box_q59;
wire   [7:0] decipher_0_i32box_address60;
reg    decipher_0_i32box_ce60;
wire   [31:0] decipher_0_i32box_q60;
wire   [7:0] decipher_0_i32box_address61;
reg    decipher_0_i32box_ce61;
wire   [31:0] decipher_0_i32box_q61;
wire   [7:0] decipher_0_i32box_address62;
reg    decipher_0_i32box_ce62;
wire   [31:0] decipher_0_i32box_q62;
wire   [7:0] decipher_0_i32box_address63;
reg    decipher_0_i32box_ce63;
wire   [31:0] decipher_0_i32box_q63;
wire   [7:0] decipher_0_i32box_address64;
reg    decipher_0_i32box_ce64;
wire   [31:0] decipher_0_i32box_q64;
wire   [7:0] decipher_0_i32box_address65;
reg    decipher_0_i32box_ce65;
wire   [31:0] decipher_0_i32box_q65;
wire   [7:0] decipher_0_i32box_address66;
reg    decipher_0_i32box_ce66;
wire   [31:0] decipher_0_i32box_q66;
wire   [7:0] decipher_0_i32box_address67;
reg    decipher_0_i32box_ce67;
wire   [31:0] decipher_0_i32box_q67;
wire   [7:0] decipher_0_i32box_address68;
reg    decipher_0_i32box_ce68;
wire   [31:0] decipher_0_i32box_q68;
wire   [7:0] decipher_0_i32box_address69;
reg    decipher_0_i32box_ce69;
wire   [31:0] decipher_0_i32box_q69;
wire   [7:0] decipher_0_i32box_address70;
reg    decipher_0_i32box_ce70;
wire   [31:0] decipher_0_i32box_q70;
wire   [7:0] decipher_0_i32box_address71;
reg    decipher_0_i32box_ce71;
wire   [31:0] decipher_0_i32box_q71;
wire   [7:0] decipher_0_i32box_address72;
reg    decipher_0_i32box_ce72;
wire   [31:0] decipher_0_i32box_q72;
wire   [7:0] decipher_0_i32box_address73;
reg    decipher_0_i32box_ce73;
wire   [31:0] decipher_0_i32box_q73;
wire   [7:0] decipher_0_i32box_address74;
reg    decipher_0_i32box_ce74;
wire   [31:0] decipher_0_i32box_q74;
wire   [7:0] decipher_0_i32box_address75;
reg    decipher_0_i32box_ce75;
wire   [31:0] decipher_0_i32box_q75;
wire   [7:0] decipher_0_i32box_address76;
reg    decipher_0_i32box_ce76;
wire   [31:0] decipher_0_i32box_q76;
wire   [7:0] decipher_0_i32box_address77;
reg    decipher_0_i32box_ce77;
wire   [31:0] decipher_0_i32box_q77;
wire   [7:0] decipher_0_i32box_address78;
reg    decipher_0_i32box_ce78;
wire   [31:0] decipher_0_i32box_q78;
wire   [7:0] decipher_0_i32box_address79;
reg    decipher_0_i32box_ce79;
wire   [31:0] decipher_0_i32box_q79;
wire   [7:0] decipher_0_i32box_address80;
reg    decipher_0_i32box_ce80;
wire   [31:0] decipher_0_i32box_q80;
wire   [7:0] decipher_0_i32box_address81;
reg    decipher_0_i32box_ce81;
wire   [31:0] decipher_0_i32box_q81;
wire   [7:0] decipher_0_i32box_address82;
reg    decipher_0_i32box_ce82;
wire   [31:0] decipher_0_i32box_q82;
wire   [7:0] decipher_0_i32box_address83;
reg    decipher_0_i32box_ce83;
wire   [31:0] decipher_0_i32box_q83;
wire   [7:0] decipher_0_i32box_address84;
reg    decipher_0_i32box_ce84;
wire   [31:0] decipher_0_i32box_q84;
wire   [7:0] decipher_0_i32box_address85;
reg    decipher_0_i32box_ce85;
wire   [31:0] decipher_0_i32box_q85;
wire   [7:0] decipher_0_i32box_address86;
reg    decipher_0_i32box_ce86;
wire   [31:0] decipher_0_i32box_q86;
wire   [7:0] decipher_0_i32box_address87;
reg    decipher_0_i32box_ce87;
wire   [31:0] decipher_0_i32box_q87;
wire   [7:0] decipher_0_i32box_address88;
reg    decipher_0_i32box_ce88;
wire   [31:0] decipher_0_i32box_q88;
wire   [7:0] decipher_0_i32box_address89;
reg    decipher_0_i32box_ce89;
wire   [31:0] decipher_0_i32box_q89;
wire   [7:0] decipher_0_i32box_address90;
reg    decipher_0_i32box_ce90;
wire   [31:0] decipher_0_i32box_q90;
wire   [7:0] decipher_0_i32box_address91;
reg    decipher_0_i32box_ce91;
wire   [31:0] decipher_0_i32box_q91;
wire   [7:0] decipher_0_i32box_address92;
reg    decipher_0_i32box_ce92;
wire   [31:0] decipher_0_i32box_q92;
wire   [7:0] decipher_0_i32box_address93;
reg    decipher_0_i32box_ce93;
wire   [31:0] decipher_0_i32box_q93;
wire   [7:0] decipher_0_i32box_address94;
reg    decipher_0_i32box_ce94;
wire   [31:0] decipher_0_i32box_q94;
wire   [7:0] decipher_0_i32box_address95;
reg    decipher_0_i32box_ce95;
wire   [31:0] decipher_0_i32box_q95;
wire   [7:0] decipher_0_i32box_address96;
reg    decipher_0_i32box_ce96;
wire   [31:0] decipher_0_i32box_q96;
wire   [7:0] decipher_0_i32box_address97;
reg    decipher_0_i32box_ce97;
wire   [31:0] decipher_0_i32box_q97;
wire   [7:0] decipher_0_i32box_address98;
reg    decipher_0_i32box_ce98;
wire   [31:0] decipher_0_i32box_q98;
wire   [7:0] decipher_0_i32box_address99;
reg    decipher_0_i32box_ce99;
wire   [31:0] decipher_0_i32box_q99;
wire   [7:0] decipher_0_i32box_address100;
reg    decipher_0_i32box_ce100;
wire   [31:0] decipher_0_i32box_q100;
wire   [7:0] decipher_0_i32box_address101;
reg    decipher_0_i32box_ce101;
wire   [31:0] decipher_0_i32box_q101;
wire   [7:0] decipher_0_i32box_address102;
reg    decipher_0_i32box_ce102;
wire   [31:0] decipher_0_i32box_q102;
wire   [7:0] decipher_0_i32box_address103;
reg    decipher_0_i32box_ce103;
wire   [31:0] decipher_0_i32box_q103;
wire   [7:0] decipher_0_i32box_address104;
reg    decipher_0_i32box_ce104;
wire   [31:0] decipher_0_i32box_q104;
wire   [7:0] decipher_0_i32box_address105;
reg    decipher_0_i32box_ce105;
wire   [31:0] decipher_0_i32box_q105;
wire   [7:0] decipher_0_i32box_address106;
reg    decipher_0_i32box_ce106;
wire   [31:0] decipher_0_i32box_q106;
wire   [7:0] decipher_0_i32box_address107;
reg    decipher_0_i32box_ce107;
wire   [31:0] decipher_0_i32box_q107;
wire   [7:0] decipher_0_i32box_address108;
reg    decipher_0_i32box_ce108;
wire   [31:0] decipher_0_i32box_q108;
wire   [7:0] decipher_0_i32box_address109;
reg    decipher_0_i32box_ce109;
wire   [31:0] decipher_0_i32box_q109;
wire   [7:0] decipher_0_i32box_address110;
reg    decipher_0_i32box_ce110;
wire   [31:0] decipher_0_i32box_q110;
wire   [7:0] decipher_0_i32box_address111;
reg    decipher_0_i32box_ce111;
wire   [31:0] decipher_0_i32box_q111;
wire   [7:0] decipher_0_i32box_address112;
reg    decipher_0_i32box_ce112;
wire   [31:0] decipher_0_i32box_q112;
wire   [7:0] decipher_0_i32box_address113;
reg    decipher_0_i32box_ce113;
wire   [31:0] decipher_0_i32box_q113;
wire   [7:0] decipher_0_i32box_address114;
reg    decipher_0_i32box_ce114;
wire   [31:0] decipher_0_i32box_q114;
wire   [7:0] decipher_0_i32box_address115;
reg    decipher_0_i32box_ce115;
wire   [31:0] decipher_0_i32box_q115;
wire   [7:0] decipher_0_i32box_address116;
reg    decipher_0_i32box_ce116;
wire   [31:0] decipher_0_i32box_q116;
wire   [7:0] decipher_0_i32box_address117;
reg    decipher_0_i32box_ce117;
wire   [31:0] decipher_0_i32box_q117;
wire   [7:0] decipher_0_i32box_address118;
reg    decipher_0_i32box_ce118;
wire   [31:0] decipher_0_i32box_q118;
wire   [7:0] decipher_0_i32box_address119;
reg    decipher_0_i32box_ce119;
wire   [31:0] decipher_0_i32box_q119;
wire   [7:0] decipher_0_i32box_address120;
reg    decipher_0_i32box_ce120;
wire   [31:0] decipher_0_i32box_q120;
wire   [7:0] decipher_0_i32box_address121;
reg    decipher_0_i32box_ce121;
wire   [31:0] decipher_0_i32box_q121;
wire   [7:0] decipher_0_i32box_address122;
reg    decipher_0_i32box_ce122;
wire   [31:0] decipher_0_i32box_q122;
wire   [7:0] decipher_0_i32box_address123;
reg    decipher_0_i32box_ce123;
wire   [31:0] decipher_0_i32box_q123;
wire   [7:0] decipher_0_i32box_address124;
reg    decipher_0_i32box_ce124;
wire   [31:0] decipher_0_i32box_q124;
wire   [7:0] decipher_0_i32box_address125;
reg    decipher_0_i32box_ce125;
wire   [31:0] decipher_0_i32box_q125;
wire   [7:0] decipher_0_i32box_address126;
reg    decipher_0_i32box_ce126;
wire   [31:0] decipher_0_i32box_q126;
wire   [7:0] decipher_0_i32box_address127;
reg    decipher_0_i32box_ce127;
wire   [31:0] decipher_0_i32box_q127;
wire   [7:0] decipher_0_i32box_address128;
reg    decipher_0_i32box_ce128;
wire   [31:0] decipher_0_i32box_q128;
wire   [7:0] decipher_0_i32box_address129;
reg    decipher_0_i32box_ce129;
wire   [31:0] decipher_0_i32box_q129;
wire   [7:0] decipher_0_i32box_address130;
reg    decipher_0_i32box_ce130;
wire   [31:0] decipher_0_i32box_q130;
wire   [7:0] decipher_0_i32box_address131;
reg    decipher_0_i32box_ce131;
wire   [31:0] decipher_0_i32box_q131;
wire   [7:0] decipher_0_i32box_address132;
reg    decipher_0_i32box_ce132;
wire   [31:0] decipher_0_i32box_q132;
wire   [7:0] decipher_0_i32box_address133;
reg    decipher_0_i32box_ce133;
wire   [31:0] decipher_0_i32box_q133;
wire   [7:0] decipher_0_i32box_address134;
reg    decipher_0_i32box_ce134;
wire   [31:0] decipher_0_i32box_q134;
wire   [7:0] decipher_0_i32box_address135;
reg    decipher_0_i32box_ce135;
wire   [31:0] decipher_0_i32box_q135;
wire   [7:0] decipher_0_i32box_address136;
reg    decipher_0_i32box_ce136;
wire   [31:0] decipher_0_i32box_q136;
wire   [7:0] decipher_0_i32box_address137;
reg    decipher_0_i32box_ce137;
wire   [31:0] decipher_0_i32box_q137;
wire   [7:0] decipher_0_i32box_address138;
reg    decipher_0_i32box_ce138;
wire   [31:0] decipher_0_i32box_q138;
wire   [7:0] decipher_0_i32box_address139;
reg    decipher_0_i32box_ce139;
wire   [31:0] decipher_0_i32box_q139;
wire   [7:0] decipher_0_i32box_address140;
reg    decipher_0_i32box_ce140;
wire   [31:0] decipher_0_i32box_q140;
wire   [7:0] decipher_0_i32box_address141;
reg    decipher_0_i32box_ce141;
wire   [31:0] decipher_0_i32box_q141;
wire   [7:0] decipher_0_i32box_address142;
reg    decipher_0_i32box_ce142;
wire   [31:0] decipher_0_i32box_q142;
wire   [7:0] decipher_0_i32box_address143;
reg    decipher_0_i32box_ce143;
wire   [31:0] decipher_0_i32box_q143;
wire   [7:0] decipher_0_i32box_address144;
reg    decipher_0_i32box_ce144;
wire   [31:0] decipher_0_i32box_q144;
wire   [7:0] decipher_0_i32box_address145;
reg    decipher_0_i32box_ce145;
wire   [31:0] decipher_0_i32box_q145;
wire   [7:0] decipher_0_i32box_address146;
reg    decipher_0_i32box_ce146;
wire   [31:0] decipher_0_i32box_q146;
wire   [7:0] decipher_0_i32box_address147;
reg    decipher_0_i32box_ce147;
wire   [31:0] decipher_0_i32box_q147;
wire   [7:0] decipher_0_i32box_address148;
reg    decipher_0_i32box_ce148;
wire   [31:0] decipher_0_i32box_q148;
wire   [7:0] decipher_0_i32box_address149;
reg    decipher_0_i32box_ce149;
wire   [31:0] decipher_0_i32box_q149;
wire   [7:0] decipher_0_i32box_address150;
reg    decipher_0_i32box_ce150;
wire   [31:0] decipher_0_i32box_q150;
wire   [7:0] decipher_0_i32box_address151;
reg    decipher_0_i32box_ce151;
wire   [31:0] decipher_0_i32box_q151;
wire   [7:0] decipher_0_i32box_address152;
reg    decipher_0_i32box_ce152;
wire   [31:0] decipher_0_i32box_q152;
wire   [7:0] decipher_0_i32box_address153;
reg    decipher_0_i32box_ce153;
wire   [31:0] decipher_0_i32box_q153;
wire   [7:0] decipher_0_i32box_address154;
reg    decipher_0_i32box_ce154;
wire   [31:0] decipher_0_i32box_q154;
wire   [7:0] decipher_0_i32box_address155;
reg    decipher_0_i32box_ce155;
wire   [31:0] decipher_0_i32box_q155;
wire   [7:0] decipher_0_i32box_address156;
reg    decipher_0_i32box_ce156;
wire   [31:0] decipher_0_i32box_q156;
wire   [7:0] decipher_0_i32box_address157;
reg    decipher_0_i32box_ce157;
wire   [31:0] decipher_0_i32box_q157;
wire   [7:0] decipher_0_i32box_address158;
reg    decipher_0_i32box_ce158;
wire   [31:0] decipher_0_i32box_q158;
wire   [7:0] decipher_0_i32box_address159;
reg    decipher_0_i32box_ce159;
wire   [31:0] decipher_0_i32box_q159;
wire   [7:0] decipher_0_i32box_address160;
reg    decipher_0_i32box_ce160;
wire   [31:0] decipher_0_i32box_q160;
wire   [7:0] decipher_0_i32box_address161;
reg    decipher_0_i32box_ce161;
wire   [31:0] decipher_0_i32box_q161;
wire   [7:0] decipher_0_i32box_address162;
reg    decipher_0_i32box_ce162;
wire   [31:0] decipher_0_i32box_q162;
wire   [7:0] decipher_0_i32box_address163;
reg    decipher_0_i32box_ce163;
wire   [31:0] decipher_0_i32box_q163;
wire   [7:0] decipher_0_i32box_address164;
reg    decipher_0_i32box_ce164;
wire   [31:0] decipher_0_i32box_q164;
wire   [7:0] decipher_0_i32box_address165;
reg    decipher_0_i32box_ce165;
wire   [31:0] decipher_0_i32box_q165;
wire   [7:0] decipher_0_i32box_address166;
reg    decipher_0_i32box_ce166;
wire   [31:0] decipher_0_i32box_q166;
wire   [7:0] decipher_0_i32box_address167;
reg    decipher_0_i32box_ce167;
wire   [31:0] decipher_0_i32box_q167;
wire   [7:0] decipher_0_i32box_address168;
reg    decipher_0_i32box_ce168;
wire   [31:0] decipher_0_i32box_q168;
wire   [7:0] decipher_0_i32box_address169;
reg    decipher_0_i32box_ce169;
wire   [31:0] decipher_0_i32box_q169;
wire   [7:0] decipher_0_i32box_address170;
reg    decipher_0_i32box_ce170;
wire   [31:0] decipher_0_i32box_q170;
wire   [7:0] decipher_0_i32box_address171;
reg    decipher_0_i32box_ce171;
wire   [31:0] decipher_0_i32box_q171;
wire   [7:0] decipher_0_i32box_address172;
reg    decipher_0_i32box_ce172;
wire   [31:0] decipher_0_i32box_q172;
wire   [7:0] decipher_0_i32box_address173;
reg    decipher_0_i32box_ce173;
wire   [31:0] decipher_0_i32box_q173;
wire   [7:0] decipher_0_i32box_address174;
reg    decipher_0_i32box_ce174;
wire   [31:0] decipher_0_i32box_q174;
wire   [7:0] decipher_0_i32box_address175;
reg    decipher_0_i32box_ce175;
wire   [31:0] decipher_0_i32box_q175;
reg   [127:0] p_read_2_reg_17950;
wire    ap_block_pp0_stage0_11001;
reg   [127:0] p_read_3_reg_17955;
reg   [127:0] p_read_3_reg_17955_pp0_iter1_reg;
reg   [127:0] p_read_3_reg_17955_pp0_iter2_reg;
reg   [127:0] p_read_4_reg_17960;
reg   [127:0] p_read_4_reg_17960_pp0_iter1_reg;
reg   [127:0] p_read_4_reg_17960_pp0_iter2_reg;
reg   [127:0] p_read_4_reg_17960_pp0_iter3_reg;
reg   [127:0] p_read_4_reg_17960_pp0_iter4_reg;
reg   [127:0] p_read_5_reg_17965;
reg   [127:0] p_read_5_reg_17965_pp0_iter1_reg;
reg   [127:0] p_read_5_reg_17965_pp0_iter2_reg;
reg   [127:0] p_read_5_reg_17965_pp0_iter3_reg;
reg   [127:0] p_read_5_reg_17965_pp0_iter4_reg;
reg   [127:0] p_read_5_reg_17965_pp0_iter5_reg;
reg   [127:0] p_read_5_reg_17965_pp0_iter6_reg;
reg   [127:0] p_read_6_reg_17970;
reg   [127:0] p_read_6_reg_17970_pp0_iter1_reg;
reg   [127:0] p_read_6_reg_17970_pp0_iter2_reg;
reg   [127:0] p_read_6_reg_17970_pp0_iter3_reg;
reg   [127:0] p_read_6_reg_17970_pp0_iter4_reg;
reg   [127:0] p_read_6_reg_17970_pp0_iter5_reg;
reg   [127:0] p_read_6_reg_17970_pp0_iter6_reg;
reg   [127:0] p_read_6_reg_17970_pp0_iter7_reg;
reg   [127:0] p_read_6_reg_17970_pp0_iter8_reg;
reg   [127:0] p_read_7_reg_17975;
reg   [127:0] p_read_7_reg_17975_pp0_iter1_reg;
reg   [127:0] p_read_7_reg_17975_pp0_iter2_reg;
reg   [127:0] p_read_7_reg_17975_pp0_iter3_reg;
reg   [127:0] p_read_7_reg_17975_pp0_iter4_reg;
reg   [127:0] p_read_7_reg_17975_pp0_iter5_reg;
reg   [127:0] p_read_7_reg_17975_pp0_iter6_reg;
reg   [127:0] p_read_7_reg_17975_pp0_iter7_reg;
reg   [127:0] p_read_7_reg_17975_pp0_iter8_reg;
reg   [127:0] p_read_7_reg_17975_pp0_iter9_reg;
reg   [127:0] p_read_7_reg_17975_pp0_iter10_reg;
reg   [127:0] p_read_8_reg_17980;
reg   [127:0] p_read_8_reg_17980_pp0_iter1_reg;
reg   [127:0] p_read_8_reg_17980_pp0_iter2_reg;
reg   [127:0] p_read_8_reg_17980_pp0_iter3_reg;
reg   [127:0] p_read_8_reg_17980_pp0_iter4_reg;
reg   [127:0] p_read_8_reg_17980_pp0_iter5_reg;
reg   [127:0] p_read_8_reg_17980_pp0_iter6_reg;
reg   [127:0] p_read_8_reg_17980_pp0_iter7_reg;
reg   [127:0] p_read_8_reg_17980_pp0_iter8_reg;
reg   [127:0] p_read_8_reg_17980_pp0_iter9_reg;
reg   [127:0] p_read_8_reg_17980_pp0_iter10_reg;
reg   [127:0] p_read_8_reg_17980_pp0_iter11_reg;
reg   [127:0] p_read_8_reg_17980_pp0_iter12_reg;
reg   [127:0] p_read_9_reg_17985;
reg   [127:0] p_read_9_reg_17985_pp0_iter1_reg;
reg   [127:0] p_read_9_reg_17985_pp0_iter2_reg;
reg   [127:0] p_read_9_reg_17985_pp0_iter3_reg;
reg   [127:0] p_read_9_reg_17985_pp0_iter4_reg;
reg   [127:0] p_read_9_reg_17985_pp0_iter5_reg;
reg   [127:0] p_read_9_reg_17985_pp0_iter6_reg;
reg   [127:0] p_read_9_reg_17985_pp0_iter7_reg;
reg   [127:0] p_read_9_reg_17985_pp0_iter8_reg;
reg   [127:0] p_read_9_reg_17985_pp0_iter9_reg;
reg   [127:0] p_read_9_reg_17985_pp0_iter10_reg;
reg   [127:0] p_read_9_reg_17985_pp0_iter11_reg;
reg   [127:0] p_read_9_reg_17985_pp0_iter12_reg;
reg   [127:0] p_read_9_reg_17985_pp0_iter13_reg;
reg   [127:0] p_read_9_reg_17985_pp0_iter14_reg;
reg   [127:0] p_read_10_reg_17990;
reg   [127:0] p_read_10_reg_17990_pp0_iter1_reg;
reg   [127:0] p_read_10_reg_17990_pp0_iter2_reg;
reg   [127:0] p_read_10_reg_17990_pp0_iter3_reg;
reg   [127:0] p_read_10_reg_17990_pp0_iter4_reg;
reg   [127:0] p_read_10_reg_17990_pp0_iter5_reg;
reg   [127:0] p_read_10_reg_17990_pp0_iter6_reg;
reg   [127:0] p_read_10_reg_17990_pp0_iter7_reg;
reg   [127:0] p_read_10_reg_17990_pp0_iter8_reg;
reg   [127:0] p_read_10_reg_17990_pp0_iter9_reg;
reg   [127:0] p_read_10_reg_17990_pp0_iter10_reg;
reg   [127:0] p_read_10_reg_17990_pp0_iter11_reg;
reg   [127:0] p_read_10_reg_17990_pp0_iter12_reg;
reg   [127:0] p_read_10_reg_17990_pp0_iter13_reg;
reg   [127:0] p_read_10_reg_17990_pp0_iter14_reg;
reg   [127:0] p_read_10_reg_17990_pp0_iter15_reg;
reg   [127:0] p_read_10_reg_17990_pp0_iter16_reg;
reg   [127:0] p_read_11_reg_17995;
reg   [127:0] p_read_11_reg_17995_pp0_iter1_reg;
reg   [127:0] p_read_11_reg_17995_pp0_iter2_reg;
reg   [127:0] p_read_11_reg_17995_pp0_iter3_reg;
reg   [127:0] p_read_11_reg_17995_pp0_iter4_reg;
reg   [127:0] p_read_11_reg_17995_pp0_iter5_reg;
reg   [127:0] p_read_11_reg_17995_pp0_iter6_reg;
reg   [127:0] p_read_11_reg_17995_pp0_iter7_reg;
reg   [127:0] p_read_11_reg_17995_pp0_iter8_reg;
reg   [127:0] p_read_11_reg_17995_pp0_iter9_reg;
reg   [127:0] p_read_11_reg_17995_pp0_iter10_reg;
reg   [127:0] p_read_11_reg_17995_pp0_iter11_reg;
reg   [127:0] p_read_11_reg_17995_pp0_iter12_reg;
reg   [127:0] p_read_11_reg_17995_pp0_iter13_reg;
reg   [127:0] p_read_11_reg_17995_pp0_iter14_reg;
reg   [127:0] p_read_11_reg_17995_pp0_iter15_reg;
reg   [127:0] p_read_11_reg_17995_pp0_iter16_reg;
reg   [127:0] p_read_11_reg_17995_pp0_iter17_reg;
reg   [127:0] p_read_11_reg_17995_pp0_iter18_reg;
reg   [127:0] p_read_12_reg_18000;
reg   [127:0] p_read_12_reg_18000_pp0_iter1_reg;
reg   [127:0] p_read_12_reg_18000_pp0_iter2_reg;
reg   [127:0] p_read_12_reg_18000_pp0_iter3_reg;
reg   [127:0] p_read_12_reg_18000_pp0_iter4_reg;
reg   [127:0] p_read_12_reg_18000_pp0_iter5_reg;
reg   [127:0] p_read_12_reg_18000_pp0_iter6_reg;
reg   [127:0] p_read_12_reg_18000_pp0_iter7_reg;
reg   [127:0] p_read_12_reg_18000_pp0_iter8_reg;
reg   [127:0] p_read_12_reg_18000_pp0_iter9_reg;
reg   [127:0] p_read_12_reg_18000_pp0_iter10_reg;
reg   [127:0] p_read_12_reg_18000_pp0_iter11_reg;
reg   [127:0] p_read_12_reg_18000_pp0_iter12_reg;
reg   [127:0] p_read_12_reg_18000_pp0_iter13_reg;
reg   [127:0] p_read_12_reg_18000_pp0_iter14_reg;
reg   [127:0] p_read_12_reg_18000_pp0_iter15_reg;
reg   [127:0] p_read_12_reg_18000_pp0_iter16_reg;
reg   [127:0] p_read_12_reg_18000_pp0_iter17_reg;
reg   [127:0] p_read_12_reg_18000_pp0_iter18_reg;
reg   [127:0] p_read_12_reg_18000_pp0_iter19_reg;
reg   [127:0] p_read_12_reg_18000_pp0_iter20_reg;
reg   [127:0] p_read13_reg_18005;
reg   [127:0] p_read13_reg_18005_pp0_iter1_reg;
reg   [127:0] p_read13_reg_18005_pp0_iter2_reg;
reg   [127:0] p_read13_reg_18005_pp0_iter3_reg;
reg   [127:0] p_read13_reg_18005_pp0_iter4_reg;
reg   [127:0] p_read13_reg_18005_pp0_iter5_reg;
reg   [127:0] p_read13_reg_18005_pp0_iter6_reg;
reg   [127:0] p_read13_reg_18005_pp0_iter7_reg;
reg   [127:0] p_read13_reg_18005_pp0_iter8_reg;
reg   [127:0] p_read13_reg_18005_pp0_iter9_reg;
reg   [127:0] p_read13_reg_18005_pp0_iter10_reg;
reg   [127:0] p_read13_reg_18005_pp0_iter11_reg;
reg   [127:0] p_read13_reg_18005_pp0_iter12_reg;
reg   [127:0] p_read13_reg_18005_pp0_iter13_reg;
reg   [127:0] p_read13_reg_18005_pp0_iter14_reg;
reg   [127:0] p_read13_reg_18005_pp0_iter15_reg;
reg   [127:0] p_read13_reg_18005_pp0_iter16_reg;
reg   [127:0] p_read13_reg_18005_pp0_iter17_reg;
reg   [127:0] p_read13_reg_18005_pp0_iter18_reg;
reg   [127:0] p_read13_reg_18005_pp0_iter19_reg;
reg   [127:0] p_read13_reg_18005_pp0_iter20_reg;
reg   [127:0] p_read13_reg_18005_pp0_iter21_reg;
reg   [127:0] p_read13_reg_18005_pp0_iter22_reg;
wire   [63:0] zext_ln708_fu_4622_p1;
wire    ap_block_pp0_stage0;
wire   [63:0] zext_ln708_4_fu_4637_p1;
wire   [63:0] zext_ln708_5_fu_4652_p1;
wire   [63:0] zext_ln708_6_fu_4667_p1;
wire   [63:0] zext_ln708_7_fu_4682_p1;
wire   [63:0] zext_ln708_8_fu_4697_p1;
wire   [63:0] zext_ln708_9_fu_4712_p1;
wire   [63:0] zext_ln708_10_fu_4727_p1;
wire   [63:0] zext_ln708_11_fu_4742_p1;
wire   [63:0] zext_ln708_12_fu_4757_p1;
wire   [63:0] zext_ln708_13_fu_4772_p1;
wire   [63:0] zext_ln708_14_fu_4787_p1;
wire   [63:0] zext_ln708_15_fu_4802_p1;
wire   [63:0] zext_ln708_16_fu_4817_p1;
wire   [63:0] zext_ln708_17_fu_4832_p1;
wire   [63:0] zext_ln708_18_fu_4847_p1;
wire   [63:0] zext_ln708_19_fu_4897_p1;
wire   [63:0] zext_ln708_20_fu_4912_p1;
wire   [63:0] zext_ln708_21_fu_4927_p1;
wire   [63:0] zext_ln708_22_fu_4942_p1;
wire   [63:0] zext_ln708_23_fu_4957_p1;
wire   [63:0] zext_ln708_24_fu_4972_p1;
wire   [63:0] zext_ln708_25_fu_4987_p1;
wire   [63:0] zext_ln708_26_fu_5002_p1;
wire   [63:0] zext_ln708_27_fu_5017_p1;
wire   [63:0] zext_ln708_28_fu_5032_p1;
wire   [63:0] zext_ln708_29_fu_5047_p1;
wire   [63:0] zext_ln708_30_fu_5062_p1;
wire   [63:0] zext_ln708_31_fu_5077_p1;
wire   [63:0] zext_ln708_32_fu_5092_p1;
wire   [63:0] zext_ln708_33_fu_5107_p1;
wire   [63:0] zext_ln708_34_fu_5122_p1;
wire   [63:0] zext_ln708_35_fu_5959_p1;
wire   [63:0] zext_ln708_36_fu_5964_p1;
wire   [63:0] zext_ln708_37_fu_5969_p1;
wire   [63:0] zext_ln708_38_fu_5974_p1;
wire   [63:0] zext_ln708_39_fu_5979_p1;
wire   [63:0] zext_ln708_40_fu_5984_p1;
wire   [63:0] zext_ln708_41_fu_5989_p1;
wire   [63:0] zext_ln708_42_fu_5994_p1;
wire   [63:0] zext_ln708_43_fu_5999_p1;
wire   [63:0] zext_ln708_44_fu_6004_p1;
wire   [63:0] zext_ln708_45_fu_6009_p1;
wire   [63:0] zext_ln708_46_fu_6014_p1;
wire   [63:0] zext_ln708_47_fu_6019_p1;
wire   [63:0] zext_ln708_48_fu_6024_p1;
wire   [63:0] zext_ln708_49_fu_6029_p1;
wire   [63:0] zext_ln708_50_fu_6034_p1;
wire   [63:0] zext_ln708_51_fu_6084_p1;
wire   [63:0] zext_ln708_52_fu_6099_p1;
wire   [63:0] zext_ln708_53_fu_6114_p1;
wire   [63:0] zext_ln708_54_fu_6129_p1;
wire   [63:0] zext_ln708_55_fu_6144_p1;
wire   [63:0] zext_ln708_56_fu_6159_p1;
wire   [63:0] zext_ln708_57_fu_6174_p1;
wire   [63:0] zext_ln708_58_fu_6189_p1;
wire   [63:0] zext_ln708_59_fu_6204_p1;
wire   [63:0] zext_ln708_60_fu_6219_p1;
wire   [63:0] zext_ln708_61_fu_6234_p1;
wire   [63:0] zext_ln708_62_fu_6249_p1;
wire   [63:0] zext_ln708_63_fu_6264_p1;
wire   [63:0] zext_ln708_64_fu_6279_p1;
wire   [63:0] zext_ln708_65_fu_6294_p1;
wire   [63:0] zext_ln708_66_fu_6309_p1;
wire   [63:0] zext_ln708_67_fu_7146_p1;
wire   [63:0] zext_ln708_68_fu_7151_p1;
wire   [63:0] zext_ln708_69_fu_7156_p1;
wire   [63:0] zext_ln708_70_fu_7161_p1;
wire   [63:0] zext_ln708_71_fu_7166_p1;
wire   [63:0] zext_ln708_72_fu_7171_p1;
wire   [63:0] zext_ln708_73_fu_7176_p1;
wire   [63:0] zext_ln708_74_fu_7181_p1;
wire   [63:0] zext_ln708_75_fu_7186_p1;
wire   [63:0] zext_ln708_76_fu_7191_p1;
wire   [63:0] zext_ln708_77_fu_7196_p1;
wire   [63:0] zext_ln708_78_fu_7201_p1;
wire   [63:0] zext_ln708_79_fu_7206_p1;
wire   [63:0] zext_ln708_80_fu_7211_p1;
wire   [63:0] zext_ln708_81_fu_7216_p1;
wire   [63:0] zext_ln708_82_fu_7221_p1;
wire   [63:0] zext_ln708_83_fu_7271_p1;
wire   [63:0] zext_ln708_84_fu_7286_p1;
wire   [63:0] zext_ln708_85_fu_7301_p1;
wire   [63:0] zext_ln708_86_fu_7316_p1;
wire   [63:0] zext_ln708_87_fu_7331_p1;
wire   [63:0] zext_ln708_88_fu_7346_p1;
wire   [63:0] zext_ln708_89_fu_7361_p1;
wire   [63:0] zext_ln708_90_fu_7376_p1;
wire   [63:0] zext_ln708_91_fu_7391_p1;
wire   [63:0] zext_ln708_92_fu_7406_p1;
wire   [63:0] zext_ln708_93_fu_7421_p1;
wire   [63:0] zext_ln708_94_fu_7436_p1;
wire   [63:0] zext_ln708_95_fu_7451_p1;
wire   [63:0] zext_ln708_96_fu_7466_p1;
wire   [63:0] zext_ln708_97_fu_7481_p1;
wire   [63:0] zext_ln708_98_fu_7496_p1;
wire   [63:0] zext_ln708_99_fu_8333_p1;
wire   [63:0] zext_ln708_100_fu_8338_p1;
wire   [63:0] zext_ln708_101_fu_8343_p1;
wire   [63:0] zext_ln708_102_fu_8348_p1;
wire   [63:0] zext_ln708_103_fu_8353_p1;
wire   [63:0] zext_ln708_104_fu_8358_p1;
wire   [63:0] zext_ln708_105_fu_8363_p1;
wire   [63:0] zext_ln708_106_fu_8368_p1;
wire   [63:0] zext_ln708_107_fu_8373_p1;
wire   [63:0] zext_ln708_108_fu_8378_p1;
wire   [63:0] zext_ln708_109_fu_8383_p1;
wire   [63:0] zext_ln708_110_fu_8388_p1;
wire   [63:0] zext_ln708_111_fu_8393_p1;
wire   [63:0] zext_ln708_112_fu_8398_p1;
wire   [63:0] zext_ln708_113_fu_8403_p1;
wire   [63:0] zext_ln708_114_fu_8408_p1;
wire   [63:0] zext_ln708_115_fu_8458_p1;
wire   [63:0] zext_ln708_116_fu_8473_p1;
wire   [63:0] zext_ln708_117_fu_8488_p1;
wire   [63:0] zext_ln708_118_fu_8503_p1;
wire   [63:0] zext_ln708_119_fu_8518_p1;
wire   [63:0] zext_ln708_120_fu_8533_p1;
wire   [63:0] zext_ln708_121_fu_8548_p1;
wire   [63:0] zext_ln708_122_fu_8563_p1;
wire   [63:0] zext_ln708_123_fu_8578_p1;
wire   [63:0] zext_ln708_124_fu_8593_p1;
wire   [63:0] zext_ln708_125_fu_8608_p1;
wire   [63:0] zext_ln708_126_fu_8623_p1;
wire   [63:0] zext_ln708_127_fu_8638_p1;
wire   [63:0] zext_ln708_128_fu_8653_p1;
wire   [63:0] zext_ln708_129_fu_8668_p1;
wire   [63:0] zext_ln708_130_fu_8683_p1;
wire   [63:0] zext_ln708_131_fu_9520_p1;
wire   [63:0] zext_ln708_132_fu_9525_p1;
wire   [63:0] zext_ln708_133_fu_9530_p1;
wire   [63:0] zext_ln708_134_fu_9535_p1;
wire   [63:0] zext_ln708_135_fu_9540_p1;
wire   [63:0] zext_ln708_136_fu_9545_p1;
wire   [63:0] zext_ln708_137_fu_9550_p1;
wire   [63:0] zext_ln708_138_fu_9555_p1;
wire   [63:0] zext_ln708_139_fu_9560_p1;
wire   [63:0] zext_ln708_140_fu_9565_p1;
wire   [63:0] zext_ln708_141_fu_9570_p1;
wire   [63:0] zext_ln708_142_fu_9575_p1;
wire   [63:0] zext_ln708_143_fu_9580_p1;
wire   [63:0] zext_ln708_144_fu_9585_p1;
wire   [63:0] zext_ln708_145_fu_9590_p1;
wire   [63:0] zext_ln708_146_fu_9595_p1;
wire   [63:0] zext_ln708_147_fu_9645_p1;
wire   [63:0] zext_ln708_148_fu_9660_p1;
wire   [63:0] zext_ln708_149_fu_9675_p1;
wire   [63:0] zext_ln708_150_fu_9690_p1;
wire   [63:0] zext_ln708_151_fu_9705_p1;
wire   [63:0] zext_ln708_152_fu_9720_p1;
wire   [63:0] zext_ln708_153_fu_9735_p1;
wire   [63:0] zext_ln708_154_fu_9750_p1;
wire   [63:0] zext_ln708_155_fu_9765_p1;
wire   [63:0] zext_ln708_156_fu_9780_p1;
wire   [63:0] zext_ln708_157_fu_9795_p1;
wire   [63:0] zext_ln708_158_fu_9810_p1;
wire   [63:0] zext_ln708_159_fu_9825_p1;
wire   [63:0] zext_ln708_160_fu_9840_p1;
wire   [63:0] zext_ln708_161_fu_9855_p1;
wire   [63:0] zext_ln708_162_fu_9870_p1;
wire   [63:0] zext_ln708_163_fu_10707_p1;
wire   [63:0] zext_ln708_164_fu_10712_p1;
wire   [63:0] zext_ln708_165_fu_10717_p1;
wire   [63:0] zext_ln708_166_fu_10722_p1;
wire   [63:0] zext_ln708_167_fu_10727_p1;
wire   [63:0] zext_ln708_168_fu_10732_p1;
wire   [63:0] zext_ln708_169_fu_10737_p1;
wire   [63:0] zext_ln708_170_fu_10742_p1;
wire   [63:0] zext_ln708_171_fu_10747_p1;
wire   [63:0] zext_ln708_172_fu_10752_p1;
wire   [63:0] zext_ln708_173_fu_10757_p1;
wire   [63:0] zext_ln708_174_fu_10762_p1;
wire   [63:0] zext_ln708_175_fu_10767_p1;
wire   [63:0] zext_ln708_176_fu_10772_p1;
wire   [63:0] zext_ln708_177_fu_10777_p1;
wire   [63:0] zext_ln708_178_fu_10782_p1;
wire   [63:0] zext_ln708_179_fu_10832_p1;
wire   [63:0] zext_ln708_180_fu_10847_p1;
wire   [63:0] zext_ln708_181_fu_10862_p1;
wire   [63:0] zext_ln708_182_fu_10877_p1;
wire   [63:0] zext_ln708_183_fu_10892_p1;
wire   [63:0] zext_ln708_184_fu_10907_p1;
wire   [63:0] zext_ln708_185_fu_10922_p1;
wire   [63:0] zext_ln708_186_fu_10937_p1;
wire   [63:0] zext_ln708_187_fu_10952_p1;
wire   [63:0] zext_ln708_188_fu_10967_p1;
wire   [63:0] zext_ln708_189_fu_10982_p1;
wire   [63:0] zext_ln708_190_fu_10997_p1;
wire   [63:0] zext_ln708_191_fu_11012_p1;
wire   [63:0] zext_ln708_192_fu_11027_p1;
wire   [63:0] zext_ln708_193_fu_11042_p1;
wire   [63:0] zext_ln708_194_fu_11057_p1;
wire   [63:0] zext_ln708_195_fu_11894_p1;
wire   [63:0] zext_ln708_196_fu_11899_p1;
wire   [63:0] zext_ln708_197_fu_11904_p1;
wire   [63:0] zext_ln708_198_fu_11909_p1;
wire   [63:0] zext_ln708_199_fu_11914_p1;
wire   [63:0] zext_ln708_200_fu_11919_p1;
wire   [63:0] zext_ln708_201_fu_11924_p1;
wire   [63:0] zext_ln708_202_fu_11929_p1;
wire   [63:0] zext_ln708_203_fu_11934_p1;
wire   [63:0] zext_ln708_204_fu_11939_p1;
wire   [63:0] zext_ln708_205_fu_11944_p1;
wire   [63:0] zext_ln708_206_fu_11949_p1;
wire   [63:0] zext_ln708_207_fu_11954_p1;
wire   [63:0] zext_ln708_208_fu_11959_p1;
wire   [63:0] zext_ln708_209_fu_11964_p1;
wire   [63:0] zext_ln708_210_fu_11969_p1;
wire   [63:0] zext_ln708_211_fu_12019_p1;
wire   [63:0] zext_ln708_212_fu_12034_p1;
wire   [63:0] zext_ln708_213_fu_12049_p1;
wire   [63:0] zext_ln708_214_fu_12064_p1;
wire   [63:0] zext_ln708_215_fu_12079_p1;
wire   [63:0] zext_ln708_216_fu_12094_p1;
wire   [63:0] zext_ln708_217_fu_12109_p1;
wire   [63:0] zext_ln708_218_fu_12124_p1;
wire   [63:0] zext_ln708_219_fu_12139_p1;
wire   [63:0] zext_ln708_220_fu_12154_p1;
wire   [63:0] zext_ln708_221_fu_12169_p1;
wire   [63:0] zext_ln708_222_fu_12184_p1;
wire   [63:0] zext_ln708_223_fu_12199_p1;
wire   [63:0] zext_ln708_224_fu_12214_p1;
wire   [63:0] zext_ln708_225_fu_12229_p1;
wire   [63:0] zext_ln708_226_fu_12244_p1;
wire   [63:0] zext_ln708_227_fu_13081_p1;
wire   [63:0] zext_ln708_228_fu_13086_p1;
wire   [63:0] zext_ln708_229_fu_13091_p1;
wire   [63:0] zext_ln708_230_fu_13096_p1;
wire   [63:0] zext_ln708_231_fu_13101_p1;
wire   [63:0] zext_ln708_232_fu_13106_p1;
wire   [63:0] zext_ln708_233_fu_13111_p1;
wire   [63:0] zext_ln708_234_fu_13116_p1;
wire   [63:0] zext_ln708_235_fu_13121_p1;
wire   [63:0] zext_ln708_236_fu_13126_p1;
wire   [63:0] zext_ln708_237_fu_13131_p1;
wire   [63:0] zext_ln708_238_fu_13136_p1;
wire   [63:0] zext_ln708_239_fu_13141_p1;
wire   [63:0] zext_ln708_240_fu_13146_p1;
wire   [63:0] zext_ln708_241_fu_13151_p1;
wire   [63:0] zext_ln708_242_fu_13156_p1;
wire   [63:0] zext_ln708_243_fu_13206_p1;
wire   [63:0] zext_ln708_244_fu_13221_p1;
wire   [63:0] zext_ln708_245_fu_13236_p1;
wire   [63:0] zext_ln708_246_fu_13251_p1;
wire   [63:0] zext_ln708_247_fu_13266_p1;
wire   [63:0] zext_ln708_248_fu_13281_p1;
wire   [63:0] zext_ln708_249_fu_13296_p1;
wire   [63:0] zext_ln708_250_fu_13311_p1;
wire   [63:0] zext_ln708_251_fu_13326_p1;
wire   [63:0] zext_ln708_252_fu_13341_p1;
wire   [63:0] zext_ln708_253_fu_13356_p1;
wire   [63:0] zext_ln708_254_fu_13371_p1;
wire   [63:0] zext_ln708_255_fu_13386_p1;
wire   [63:0] zext_ln708_256_fu_13401_p1;
wire   [63:0] zext_ln708_257_fu_13416_p1;
wire   [63:0] zext_ln708_258_fu_13431_p1;
wire   [63:0] zext_ln708_259_fu_14268_p1;
wire   [63:0] zext_ln708_260_fu_14273_p1;
wire   [63:0] zext_ln708_261_fu_14278_p1;
wire   [63:0] zext_ln708_262_fu_14283_p1;
wire   [63:0] zext_ln708_263_fu_14288_p1;
wire   [63:0] zext_ln708_264_fu_14293_p1;
wire   [63:0] zext_ln708_265_fu_14298_p1;
wire   [63:0] zext_ln708_266_fu_14303_p1;
wire   [63:0] zext_ln708_267_fu_14308_p1;
wire   [63:0] zext_ln708_268_fu_14313_p1;
wire   [63:0] zext_ln708_269_fu_14318_p1;
wire   [63:0] zext_ln708_270_fu_14323_p1;
wire   [63:0] zext_ln708_271_fu_14328_p1;
wire   [63:0] zext_ln708_272_fu_14333_p1;
wire   [63:0] zext_ln708_273_fu_14338_p1;
wire   [63:0] zext_ln708_274_fu_14343_p1;
wire   [63:0] zext_ln708_275_fu_14393_p1;
wire   [63:0] zext_ln708_276_fu_14408_p1;
wire   [63:0] zext_ln708_277_fu_14423_p1;
wire   [63:0] zext_ln708_278_fu_14438_p1;
wire   [63:0] zext_ln708_279_fu_14453_p1;
wire   [63:0] zext_ln708_280_fu_14468_p1;
wire   [63:0] zext_ln708_281_fu_14483_p1;
wire   [63:0] zext_ln708_282_fu_14498_p1;
wire   [63:0] zext_ln708_283_fu_14513_p1;
wire   [63:0] zext_ln708_284_fu_14528_p1;
wire   [63:0] zext_ln708_285_fu_14543_p1;
wire   [63:0] zext_ln708_286_fu_14558_p1;
wire   [63:0] zext_ln708_287_fu_14573_p1;
wire   [63:0] zext_ln708_288_fu_14588_p1;
wire   [63:0] zext_ln708_289_fu_14603_p1;
wire   [63:0] zext_ln708_290_fu_14618_p1;
wire   [63:0] zext_ln708_291_fu_15455_p1;
wire   [63:0] zext_ln708_292_fu_15460_p1;
wire   [63:0] zext_ln708_293_fu_15465_p1;
wire   [63:0] zext_ln708_294_fu_15470_p1;
wire   [63:0] zext_ln708_295_fu_15475_p1;
wire   [63:0] zext_ln708_296_fu_15480_p1;
wire   [63:0] zext_ln708_297_fu_15485_p1;
wire   [63:0] zext_ln708_298_fu_15490_p1;
wire   [63:0] zext_ln708_299_fu_15495_p1;
wire   [63:0] zext_ln708_300_fu_15500_p1;
wire   [63:0] zext_ln708_301_fu_15505_p1;
wire   [63:0] zext_ln708_302_fu_15510_p1;
wire   [63:0] zext_ln708_303_fu_15515_p1;
wire   [63:0] zext_ln708_304_fu_15520_p1;
wire   [63:0] zext_ln708_305_fu_15525_p1;
wire   [63:0] zext_ln708_306_fu_15530_p1;
wire   [63:0] zext_ln708_307_fu_15580_p1;
wire   [63:0] zext_ln708_308_fu_15595_p1;
wire   [63:0] zext_ln708_309_fu_15610_p1;
wire   [63:0] zext_ln708_310_fu_15625_p1;
wire   [63:0] zext_ln708_311_fu_15640_p1;
wire   [63:0] zext_ln708_312_fu_15655_p1;
wire   [63:0] zext_ln708_313_fu_15670_p1;
wire   [63:0] zext_ln708_314_fu_15685_p1;
wire   [63:0] zext_ln708_315_fu_15700_p1;
wire   [63:0] zext_ln708_316_fu_15715_p1;
wire   [63:0] zext_ln708_317_fu_15730_p1;
wire   [63:0] zext_ln708_318_fu_15745_p1;
wire   [63:0] zext_ln708_319_fu_15760_p1;
wire   [63:0] zext_ln708_320_fu_15775_p1;
wire   [63:0] zext_ln708_321_fu_15790_p1;
wire   [63:0] zext_ln708_322_fu_15805_p1;
wire   [63:0] zext_ln708_323_fu_16642_p1;
wire   [63:0] zext_ln708_324_fu_16647_p1;
wire   [63:0] zext_ln708_325_fu_16652_p1;
wire   [63:0] zext_ln708_326_fu_16657_p1;
wire   [63:0] zext_ln708_327_fu_16662_p1;
wire   [63:0] zext_ln708_328_fu_16667_p1;
wire   [63:0] zext_ln708_329_fu_16672_p1;
wire   [63:0] zext_ln708_330_fu_16677_p1;
wire   [63:0] zext_ln708_331_fu_16682_p1;
wire   [63:0] zext_ln708_332_fu_16687_p1;
wire   [63:0] zext_ln708_333_fu_16692_p1;
wire   [63:0] zext_ln708_334_fu_16697_p1;
wire   [63:0] zext_ln708_335_fu_16702_p1;
wire   [63:0] zext_ln708_336_fu_16707_p1;
wire   [63:0] zext_ln708_337_fu_16712_p1;
wire   [63:0] zext_ln708_338_fu_16717_p1;
wire   [63:0] zext_ln708_339_fu_16767_p1;
wire   [63:0] zext_ln708_340_fu_16782_p1;
wire   [63:0] zext_ln708_341_fu_16797_p1;
wire   [63:0] zext_ln708_342_fu_16812_p1;
wire   [63:0] zext_ln708_343_fu_16827_p1;
wire   [63:0] zext_ln708_344_fu_16842_p1;
wire   [63:0] zext_ln708_345_fu_16857_p1;
wire   [63:0] zext_ln708_346_fu_16872_p1;
wire   [63:0] zext_ln708_347_fu_16887_p1;
wire   [63:0] zext_ln708_348_fu_16902_p1;
wire   [63:0] zext_ln708_349_fu_16917_p1;
wire   [63:0] zext_ln708_350_fu_16932_p1;
wire   [63:0] zext_ln708_351_fu_16947_p1;
wire   [63:0] zext_ln708_352_fu_16962_p1;
wire   [63:0] zext_ln708_353_fu_16977_p1;
wire   [63:0] zext_ln708_354_fu_16992_p1;
wire   [63:0] zext_ln708_355_fu_17829_p1;
wire   [63:0] zext_ln708_356_fu_17834_p1;
wire   [63:0] zext_ln708_357_fu_17839_p1;
wire   [63:0] zext_ln708_358_fu_17844_p1;
wire   [63:0] zext_ln708_359_fu_17849_p1;
wire   [63:0] zext_ln708_360_fu_17854_p1;
wire   [63:0] zext_ln708_361_fu_17859_p1;
wire   [63:0] zext_ln708_362_fu_17864_p1;
wire   [63:0] zext_ln708_363_fu_17869_p1;
wire   [63:0] zext_ln708_364_fu_17874_p1;
wire   [63:0] zext_ln708_365_fu_17879_p1;
wire   [63:0] zext_ln708_366_fu_17884_p1;
wire   [63:0] zext_ln708_367_fu_17889_p1;
wire   [63:0] zext_ln708_368_fu_17894_p1;
wire   [63:0] zext_ln708_369_fu_17899_p1;
wire   [63:0] zext_ln708_370_fu_17904_p1;
wire   [127:0] ret_V_fu_4612_p2;
wire   [7:0] trunc_ln708_fu_4618_p1;
wire   [7:0] tmp_s_fu_4627_p4;
wire   [7:0] tmp_14_fu_4642_p4;
wire   [7:0] tmp_15_fu_4657_p4;
wire   [7:0] tmp_16_fu_4672_p4;
wire   [7:0] tmp_17_fu_4687_p4;
wire   [7:0] tmp_18_fu_4702_p4;
wire   [7:0] tmp_19_fu_4717_p4;
wire   [7:0] tmp_20_fu_4732_p4;
wire   [7:0] tmp_21_fu_4747_p4;
wire   [7:0] tmp_22_fu_4762_p4;
wire   [7:0] tmp_23_fu_4777_p4;
wire   [7:0] tmp_24_fu_4792_p4;
wire   [7:0] tmp_25_fu_4807_p4;
wire   [7:0] tmp_26_fu_4822_p4;
wire   [7:0] tmp_27_fu_4837_p4;
wire   [127:0] p_Result_s_fu_4852_p17;
wire   [127:0] state_V_24_fu_4888_p2;
wire   [7:0] trunc_ln708_1_fu_4893_p1;
wire   [7:0] tmp_31_fu_4902_p4;
wire   [7:0] tmp_35_fu_4917_p4;
wire   [7:0] tmp_39_fu_4932_p4;
wire   [7:0] tmp_43_fu_4947_p4;
wire   [7:0] tmp_47_fu_4962_p4;
wire   [7:0] tmp_51_fu_4977_p4;
wire   [7:0] tmp_55_fu_4992_p4;
wire   [7:0] tmp_59_fu_5007_p4;
wire   [7:0] tmp_63_fu_5022_p4;
wire   [7:0] tmp_67_fu_5037_p4;
wire   [7:0] tmp_71_fu_5052_p4;
wire   [7:0] tmp_75_fu_5067_p4;
wire   [7:0] tmp_79_fu_5082_p4;
wire   [7:0] tmp_83_fu_5097_p4;
wire   [7:0] tmp_87_fu_5112_p4;
wire   [7:0] tmp_32_fu_5165_p4;
wire   [7:0] tmp_30_fu_5151_p4;
wire   [7:0] tmp_37_fu_5209_p4;
wire   [7:0] trunc_ln674_4_fu_5229_p1;
wire   [7:0] xor_ln1545_8_fu_5677_p2;
wire   [7:0] xor_ln1545_fu_5671_p2;
wire   [7:0] tmp_34_fu_5185_p4;
wire   [7:0] trunc_ln674_fu_5127_p1;
wire   [7:0] tmp_36_fu_5199_p4;
wire   [7:0] tmp_41_fu_5243_p4;
wire   [7:0] xor_ln1545_11_fu_5695_p2;
wire   [7:0] xor_ln1545_9_fu_5689_p2;
wire   [7:0] trunc_ln674_2_fu_5161_p1;
wire   [7:0] tmp_29_fu_5141_p4;
wire   [7:0] tmp_38_fu_5219_p4;
wire   [7:0] tmp_40_fu_5233_p4;
wire   [7:0] xor_ln1545_14_fu_5713_p2;
wire   [7:0] xor_ln1545_12_fu_5707_p2;
wire   [7:0] tmp_33_fu_5175_p4;
wire   [7:0] tmp_28_fu_5131_p4;
wire   [7:0] trunc_ln674_3_fu_5195_p1;
wire   [7:0] tmp_42_fu_5253_p4;
wire   [7:0] xor_ln1545_16_fu_5731_p2;
wire   [7:0] xor_ln1545_15_fu_5725_p2;
wire   [7:0] tmp_48_fu_5301_p4;
wire   [7:0] tmp_46_fu_5287_p4;
wire   [7:0] tmp_53_fu_5345_p4;
wire   [7:0] trunc_ln674_8_fu_5365_p1;
wire   [7:0] xor_ln1545_20_fu_5749_p2;
wire   [7:0] xor_ln1545_18_fu_5743_p2;
wire   [7:0] tmp_50_fu_5321_p4;
wire   [7:0] trunc_ln674_5_fu_5263_p1;
wire   [7:0] tmp_52_fu_5335_p4;
wire   [7:0] tmp_57_fu_5379_p4;
wire   [7:0] xor_ln1545_23_fu_5767_p2;
wire   [7:0] xor_ln1545_21_fu_5761_p2;
wire   [7:0] trunc_ln674_6_fu_5297_p1;
wire   [7:0] tmp_45_fu_5277_p4;
wire   [7:0] tmp_54_fu_5355_p4;
wire   [7:0] tmp_56_fu_5369_p4;
wire   [7:0] xor_ln1545_26_fu_5785_p2;
wire   [7:0] xor_ln1545_24_fu_5779_p2;
wire   [7:0] tmp_49_fu_5311_p4;
wire   [7:0] tmp_44_fu_5267_p4;
wire   [7:0] trunc_ln674_7_fu_5331_p1;
wire   [7:0] tmp_58_fu_5389_p4;
wire   [7:0] xor_ln1545_29_fu_5803_p2;
wire   [7:0] xor_ln1545_27_fu_5797_p2;
wire   [7:0] tmp_64_fu_5437_p4;
wire   [7:0] tmp_62_fu_5423_p4;
wire   [7:0] tmp_69_fu_5481_p4;
wire   [7:0] trunc_ln674_12_fu_5501_p1;
wire   [7:0] xor_ln1545_32_fu_5821_p2;
wire   [7:0] xor_ln1545_30_fu_5815_p2;
wire   [7:0] tmp_66_fu_5457_p4;
wire   [7:0] trunc_ln674_9_fu_5399_p1;
wire   [7:0] tmp_68_fu_5471_p4;
wire   [7:0] tmp_73_fu_5515_p4;
wire   [7:0] xor_ln1545_35_fu_5839_p2;
wire   [7:0] xor_ln1545_33_fu_5833_p2;
wire   [7:0] trunc_ln674_10_fu_5433_p1;
wire   [7:0] tmp_61_fu_5413_p4;
wire   [7:0] tmp_70_fu_5491_p4;
wire   [7:0] tmp_72_fu_5505_p4;
wire   [7:0] xor_ln1545_37_fu_5857_p2;
wire   [7:0] xor_ln1545_36_fu_5851_p2;
wire   [7:0] tmp_65_fu_5447_p4;
wire   [7:0] tmp_60_fu_5403_p4;
wire   [7:0] trunc_ln674_11_fu_5467_p1;
wire   [7:0] tmp_74_fu_5525_p4;
wire   [7:0] xor_ln1545_41_fu_5875_p2;
wire   [7:0] xor_ln1545_39_fu_5869_p2;
wire   [7:0] tmp_80_fu_5573_p4;
wire   [7:0] tmp_78_fu_5559_p4;
wire   [7:0] tmp_85_fu_5617_p4;
wire   [7:0] trunc_ln674_16_fu_5637_p1;
wire   [7:0] xor_ln1545_44_fu_5893_p2;
wire   [7:0] xor_ln1545_42_fu_5887_p2;
wire   [7:0] tmp_82_fu_5593_p4;
wire   [7:0] trunc_ln674_13_fu_5535_p1;
wire   [7:0] tmp_84_fu_5607_p4;
wire   [7:0] tmp_89_fu_5651_p4;
wire   [7:0] xor_ln1545_46_fu_5911_p2;
wire   [7:0] xor_ln1545_45_fu_5905_p2;
wire   [7:0] trunc_ln674_14_fu_5569_p1;
wire   [7:0] tmp_77_fu_5549_p4;
wire   [7:0] tmp_86_fu_5627_p4;
wire   [7:0] tmp_88_fu_5641_p4;
wire   [7:0] xor_ln1545_49_fu_5929_p2;
wire   [7:0] xor_ln1545_48_fu_5923_p2;
wire   [7:0] tmp_81_fu_5583_p4;
wire   [7:0] tmp_76_fu_5539_p4;
wire   [7:0] trunc_ln674_15_fu_5603_p1;
wire   [7:0] tmp_90_fu_5661_p4;
wire   [7:0] xor_ln1545_53_fu_5947_p2;
wire   [7:0] xor_ln1545_51_fu_5941_p2;
wire   [7:0] xor_ln1545_7_fu_5683_p2;
wire   [7:0] tmp_1_V_fu_5917_p2;
wire   [7:0] tmp_2_1_V_fu_5863_p2;
wire   [7:0] xor_ln1545_28_fu_5809_p2;
wire   [7:0] xor_ln1545_19_fu_5755_p2;
wire   [7:0] xor_ln1545_10_fu_5701_p2;
wire   [7:0] tmp_2_2_V_fu_5935_p2;
wire   [7:0] xor_ln1545_40_fu_5881_p2;
wire   [7:0] xor_ln1545_31_fu_5827_p2;
wire   [7:0] xor_ln1545_22_fu_5773_p2;
wire   [7:0] xor_ln1545_13_fu_5719_p2;
wire   [7:0] xor_ln1545_52_fu_5953_p2;
wire   [7:0] xor_ln1545_43_fu_5899_p2;
wire   [7:0] xor_ln1545_34_fu_5845_p2;
wire   [7:0] xor_ln1545_25_fu_5791_p2;
wire   [7:0] tmp_3_V_fu_5737_p2;
wire   [127:0] p_Result_25_fu_6039_p17;
wire   [127:0] state_V_25_fu_6075_p2;
wire   [7:0] trunc_ln708_2_fu_6080_p1;
wire   [7:0] tmp_94_fu_6089_p4;
wire   [7:0] tmp_98_fu_6104_p4;
wire   [7:0] tmp_102_fu_6119_p4;
wire   [7:0] tmp_106_fu_6134_p4;
wire   [7:0] tmp_110_fu_6149_p4;
wire   [7:0] tmp_114_fu_6164_p4;
wire   [7:0] tmp_118_fu_6179_p4;
wire   [7:0] tmp_122_fu_6194_p4;
wire   [7:0] tmp_126_fu_6209_p4;
wire   [7:0] tmp_130_fu_6224_p4;
wire   [7:0] tmp_134_fu_6239_p4;
wire   [7:0] tmp_138_fu_6254_p4;
wire   [7:0] tmp_142_fu_6269_p4;
wire   [7:0] tmp_146_fu_6284_p4;
wire   [7:0] tmp_150_fu_6299_p4;
wire   [7:0] tmp_95_fu_6352_p4;
wire   [7:0] tmp_93_fu_6338_p4;
wire   [7:0] tmp_100_fu_6396_p4;
wire   [7:0] trunc_ln674_20_fu_6416_p1;
wire   [7:0] xor_ln1545_56_fu_6864_p2;
wire   [7:0] xor_ln1545_54_fu_6858_p2;
wire   [7:0] tmp_97_fu_6372_p4;
wire   [7:0] trunc_ln674_17_fu_6314_p1;
wire   [7:0] tmp_99_fu_6386_p4;
wire   [7:0] tmp_104_fu_6430_p4;
wire   [7:0] xor_ln1545_59_fu_6882_p2;
wire   [7:0] xor_ln1545_57_fu_6876_p2;
wire   [7:0] trunc_ln674_18_fu_6348_p1;
wire   [7:0] tmp_92_fu_6328_p4;
wire   [7:0] tmp_101_fu_6406_p4;
wire   [7:0] tmp_103_fu_6420_p4;
wire   [7:0] xor_ln1545_62_fu_6900_p2;
wire   [7:0] xor_ln1545_60_fu_6894_p2;
wire   [7:0] tmp_96_fu_6362_p4;
wire   [7:0] tmp_91_fu_6318_p4;
wire   [7:0] trunc_ln674_19_fu_6382_p1;
wire   [7:0] tmp_105_fu_6440_p4;
wire   [7:0] xor_ln1545_64_fu_6918_p2;
wire   [7:0] xor_ln1545_63_fu_6912_p2;
wire   [7:0] tmp_111_fu_6488_p4;
wire   [7:0] tmp_109_fu_6474_p4;
wire   [7:0] tmp_116_fu_6532_p4;
wire   [7:0] trunc_ln674_24_fu_6552_p1;
wire   [7:0] xor_ln1545_68_fu_6936_p2;
wire   [7:0] xor_ln1545_66_fu_6930_p2;
wire   [7:0] tmp_113_fu_6508_p4;
wire   [7:0] trunc_ln674_21_fu_6450_p1;
wire   [7:0] tmp_115_fu_6522_p4;
wire   [7:0] tmp_120_fu_6566_p4;
wire   [7:0] xor_ln1545_71_fu_6954_p2;
wire   [7:0] xor_ln1545_69_fu_6948_p2;
wire   [7:0] trunc_ln674_22_fu_6484_p1;
wire   [7:0] tmp_108_fu_6464_p4;
wire   [7:0] tmp_117_fu_6542_p4;
wire   [7:0] tmp_119_fu_6556_p4;
wire   [7:0] xor_ln1545_74_fu_6972_p2;
wire   [7:0] xor_ln1545_72_fu_6966_p2;
wire   [7:0] tmp_112_fu_6498_p4;
wire   [7:0] tmp_107_fu_6454_p4;
wire   [7:0] trunc_ln674_23_fu_6518_p1;
wire   [7:0] tmp_121_fu_6576_p4;
wire   [7:0] xor_ln1545_77_fu_6990_p2;
wire   [7:0] xor_ln1545_75_fu_6984_p2;
wire   [7:0] tmp_127_fu_6624_p4;
wire   [7:0] tmp_125_fu_6610_p4;
wire   [7:0] tmp_132_fu_6668_p4;
wire   [7:0] trunc_ln674_28_fu_6688_p1;
wire   [7:0] xor_ln1545_80_fu_7008_p2;
wire   [7:0] xor_ln1545_78_fu_7002_p2;
wire   [7:0] tmp_129_fu_6644_p4;
wire   [7:0] trunc_ln674_25_fu_6586_p1;
wire   [7:0] tmp_131_fu_6658_p4;
wire   [7:0] tmp_136_fu_6702_p4;
wire   [7:0] xor_ln1545_83_fu_7026_p2;
wire   [7:0] xor_ln1545_81_fu_7020_p2;
wire   [7:0] trunc_ln674_26_fu_6620_p1;
wire   [7:0] tmp_124_fu_6600_p4;
wire   [7:0] tmp_133_fu_6678_p4;
wire   [7:0] tmp_135_fu_6692_p4;
wire   [7:0] xor_ln1545_85_fu_7044_p2;
wire   [7:0] xor_ln1545_84_fu_7038_p2;
wire   [7:0] tmp_128_fu_6634_p4;
wire   [7:0] tmp_123_fu_6590_p4;
wire   [7:0] trunc_ln674_27_fu_6654_p1;
wire   [7:0] tmp_137_fu_6712_p4;
wire   [7:0] xor_ln1545_89_fu_7062_p2;
wire   [7:0] xor_ln1545_87_fu_7056_p2;
wire   [7:0] tmp_143_fu_6760_p4;
wire   [7:0] tmp_141_fu_6746_p4;
wire   [7:0] tmp_148_fu_6804_p4;
wire   [7:0] trunc_ln674_32_fu_6824_p1;
wire   [7:0] xor_ln1545_92_fu_7080_p2;
wire   [7:0] xor_ln1545_90_fu_7074_p2;
wire   [7:0] tmp_145_fu_6780_p4;
wire   [7:0] trunc_ln674_29_fu_6722_p1;
wire   [7:0] tmp_147_fu_6794_p4;
wire   [7:0] tmp_152_fu_6838_p4;
wire   [7:0] xor_ln1545_94_fu_7098_p2;
wire   [7:0] xor_ln1545_93_fu_7092_p2;
wire   [7:0] trunc_ln674_30_fu_6756_p1;
wire   [7:0] tmp_140_fu_6736_p4;
wire   [7:0] tmp_149_fu_6814_p4;
wire   [7:0] tmp_151_fu_6828_p4;
wire   [7:0] xor_ln1545_97_fu_7116_p2;
wire   [7:0] xor_ln1545_96_fu_7110_p2;
wire   [7:0] tmp_144_fu_6770_p4;
wire   [7:0] tmp_139_fu_6726_p4;
wire   [7:0] trunc_ln674_31_fu_6790_p1;
wire   [7:0] tmp_153_fu_6848_p4;
wire   [7:0] xor_ln1545_101_fu_7134_p2;
wire   [7:0] xor_ln1545_99_fu_7128_p2;
wire   [7:0] xor_ln1545_55_fu_6870_p2;
wire   [7:0] tmp_1_V_1_fu_7104_p2;
wire   [7:0] tmp_2_1_V_1_fu_7050_p2;
wire   [7:0] xor_ln1545_76_fu_6996_p2;
wire   [7:0] xor_ln1545_67_fu_6942_p2;
wire   [7:0] xor_ln1545_58_fu_6888_p2;
wire   [7:0] tmp_2_2_V_1_fu_7122_p2;
wire   [7:0] xor_ln1545_88_fu_7068_p2;
wire   [7:0] xor_ln1545_79_fu_7014_p2;
wire   [7:0] xor_ln1545_70_fu_6960_p2;
wire   [7:0] xor_ln1545_61_fu_6906_p2;
wire   [7:0] xor_ln1545_100_fu_7140_p2;
wire   [7:0] xor_ln1545_91_fu_7086_p2;
wire   [7:0] xor_ln1545_82_fu_7032_p2;
wire   [7:0] xor_ln1545_73_fu_6978_p2;
wire   [7:0] tmp_3_V_1_fu_6924_p2;
wire   [127:0] p_Result_26_fu_7226_p17;
wire   [127:0] state_V_26_fu_7262_p2;
wire   [7:0] trunc_ln708_3_fu_7267_p1;
wire   [7:0] tmp_157_fu_7276_p4;
wire   [7:0] tmp_161_fu_7291_p4;
wire   [7:0] tmp_165_fu_7306_p4;
wire   [7:0] tmp_169_fu_7321_p4;
wire   [7:0] tmp_173_fu_7336_p4;
wire   [7:0] tmp_177_fu_7351_p4;
wire   [7:0] tmp_181_fu_7366_p4;
wire   [7:0] tmp_185_fu_7381_p4;
wire   [7:0] tmp_189_fu_7396_p4;
wire   [7:0] tmp_193_fu_7411_p4;
wire   [7:0] tmp_197_fu_7426_p4;
wire   [7:0] tmp_201_fu_7441_p4;
wire   [7:0] tmp_205_fu_7456_p4;
wire   [7:0] tmp_209_fu_7471_p4;
wire   [7:0] tmp_213_fu_7486_p4;
wire   [7:0] tmp_158_fu_7539_p4;
wire   [7:0] tmp_156_fu_7525_p4;
wire   [7:0] tmp_163_fu_7583_p4;
wire   [7:0] trunc_ln674_36_fu_7603_p1;
wire   [7:0] xor_ln1545_104_fu_8051_p2;
wire   [7:0] xor_ln1545_102_fu_8045_p2;
wire   [7:0] tmp_160_fu_7559_p4;
wire   [7:0] trunc_ln674_33_fu_7501_p1;
wire   [7:0] tmp_162_fu_7573_p4;
wire   [7:0] tmp_167_fu_7617_p4;
wire   [7:0] xor_ln1545_107_fu_8069_p2;
wire   [7:0] xor_ln1545_105_fu_8063_p2;
wire   [7:0] trunc_ln674_34_fu_7535_p1;
wire   [7:0] tmp_155_fu_7515_p4;
wire   [7:0] tmp_164_fu_7593_p4;
wire   [7:0] tmp_166_fu_7607_p4;
wire   [7:0] xor_ln1545_110_fu_8087_p2;
wire   [7:0] xor_ln1545_108_fu_8081_p2;
wire   [7:0] tmp_159_fu_7549_p4;
wire   [7:0] tmp_154_fu_7505_p4;
wire   [7:0] trunc_ln674_35_fu_7569_p1;
wire   [7:0] tmp_168_fu_7627_p4;
wire   [7:0] xor_ln1545_112_fu_8105_p2;
wire   [7:0] xor_ln1545_111_fu_8099_p2;
wire   [7:0] tmp_174_fu_7675_p4;
wire   [7:0] tmp_172_fu_7661_p4;
wire   [7:0] tmp_179_fu_7719_p4;
wire   [7:0] trunc_ln674_40_fu_7739_p1;
wire   [7:0] xor_ln1545_116_fu_8123_p2;
wire   [7:0] xor_ln1545_114_fu_8117_p2;
wire   [7:0] tmp_176_fu_7695_p4;
wire   [7:0] trunc_ln674_37_fu_7637_p1;
wire   [7:0] tmp_178_fu_7709_p4;
wire   [7:0] tmp_183_fu_7753_p4;
wire   [7:0] xor_ln1545_119_fu_8141_p2;
wire   [7:0] xor_ln1545_117_fu_8135_p2;
wire   [7:0] trunc_ln674_38_fu_7671_p1;
wire   [7:0] tmp_171_fu_7651_p4;
wire   [7:0] tmp_180_fu_7729_p4;
wire   [7:0] tmp_182_fu_7743_p4;
wire   [7:0] xor_ln1545_122_fu_8159_p2;
wire   [7:0] xor_ln1545_120_fu_8153_p2;
wire   [7:0] tmp_175_fu_7685_p4;
wire   [7:0] tmp_170_fu_7641_p4;
wire   [7:0] trunc_ln674_39_fu_7705_p1;
wire   [7:0] tmp_184_fu_7763_p4;
wire   [7:0] xor_ln1545_125_fu_8177_p2;
wire   [7:0] xor_ln1545_123_fu_8171_p2;
wire   [7:0] tmp_190_fu_7811_p4;
wire   [7:0] tmp_188_fu_7797_p4;
wire   [7:0] tmp_195_fu_7855_p4;
wire   [7:0] trunc_ln674_44_fu_7875_p1;
wire   [7:0] xor_ln1545_128_fu_8195_p2;
wire   [7:0] xor_ln1545_126_fu_8189_p2;
wire   [7:0] tmp_192_fu_7831_p4;
wire   [7:0] trunc_ln674_41_fu_7773_p1;
wire   [7:0] tmp_194_fu_7845_p4;
wire   [7:0] tmp_199_fu_7889_p4;
wire   [7:0] xor_ln1545_131_fu_8213_p2;
wire   [7:0] xor_ln1545_129_fu_8207_p2;
wire   [7:0] trunc_ln674_42_fu_7807_p1;
wire   [7:0] tmp_187_fu_7787_p4;
wire   [7:0] tmp_196_fu_7865_p4;
wire   [7:0] tmp_198_fu_7879_p4;
wire   [7:0] xor_ln1545_133_fu_8231_p2;
wire   [7:0] xor_ln1545_132_fu_8225_p2;
wire   [7:0] tmp_191_fu_7821_p4;
wire   [7:0] tmp_186_fu_7777_p4;
wire   [7:0] trunc_ln674_43_fu_7841_p1;
wire   [7:0] tmp_200_fu_7899_p4;
wire   [7:0] xor_ln1545_137_fu_8249_p2;
wire   [7:0] xor_ln1545_135_fu_8243_p2;
wire   [7:0] tmp_206_fu_7947_p4;
wire   [7:0] tmp_204_fu_7933_p4;
wire   [7:0] tmp_211_fu_7991_p4;
wire   [7:0] trunc_ln674_48_fu_8011_p1;
wire   [7:0] xor_ln1545_140_fu_8267_p2;
wire   [7:0] xor_ln1545_138_fu_8261_p2;
wire   [7:0] tmp_208_fu_7967_p4;
wire   [7:0] trunc_ln674_45_fu_7909_p1;
wire   [7:0] tmp_210_fu_7981_p4;
wire   [7:0] tmp_215_fu_8025_p4;
wire   [7:0] xor_ln1545_142_fu_8285_p2;
wire   [7:0] xor_ln1545_141_fu_8279_p2;
wire   [7:0] trunc_ln674_46_fu_7943_p1;
wire   [7:0] tmp_203_fu_7923_p4;
wire   [7:0] tmp_212_fu_8001_p4;
wire   [7:0] tmp_214_fu_8015_p4;
wire   [7:0] xor_ln1545_145_fu_8303_p2;
wire   [7:0] xor_ln1545_144_fu_8297_p2;
wire   [7:0] tmp_207_fu_7957_p4;
wire   [7:0] tmp_202_fu_7913_p4;
wire   [7:0] trunc_ln674_47_fu_7977_p1;
wire   [7:0] tmp_216_fu_8035_p4;
wire   [7:0] xor_ln1545_149_fu_8321_p2;
wire   [7:0] xor_ln1545_147_fu_8315_p2;
wire   [7:0] xor_ln1545_103_fu_8057_p2;
wire   [7:0] tmp_1_V_2_fu_8291_p2;
wire   [7:0] tmp_2_1_V_2_fu_8237_p2;
wire   [7:0] xor_ln1545_124_fu_8183_p2;
wire   [7:0] xor_ln1545_115_fu_8129_p2;
wire   [7:0] xor_ln1545_106_fu_8075_p2;
wire   [7:0] tmp_2_2_V_2_fu_8309_p2;
wire   [7:0] xor_ln1545_136_fu_8255_p2;
wire   [7:0] xor_ln1545_127_fu_8201_p2;
wire   [7:0] xor_ln1545_118_fu_8147_p2;
wire   [7:0] xor_ln1545_109_fu_8093_p2;
wire   [7:0] xor_ln1545_148_fu_8327_p2;
wire   [7:0] xor_ln1545_139_fu_8273_p2;
wire   [7:0] xor_ln1545_130_fu_8219_p2;
wire   [7:0] xor_ln1545_121_fu_8165_p2;
wire   [7:0] tmp_3_V_2_fu_8111_p2;
wire   [127:0] p_Result_27_fu_8413_p17;
wire   [127:0] state_V_27_fu_8449_p2;
wire   [7:0] trunc_ln708_4_fu_8454_p1;
wire   [7:0] tmp_220_fu_8463_p4;
wire   [7:0] tmp_224_fu_8478_p4;
wire   [7:0] tmp_228_fu_8493_p4;
wire   [7:0] tmp_232_fu_8508_p4;
wire   [7:0] tmp_236_fu_8523_p4;
wire   [7:0] tmp_240_fu_8538_p4;
wire   [7:0] tmp_244_fu_8553_p4;
wire   [7:0] tmp_248_fu_8568_p4;
wire   [7:0] tmp_252_fu_8583_p4;
wire   [7:0] tmp_256_fu_8598_p4;
wire   [7:0] tmp_260_fu_8613_p4;
wire   [7:0] tmp_264_fu_8628_p4;
wire   [7:0] tmp_268_fu_8643_p4;
wire   [7:0] tmp_272_fu_8658_p4;
wire   [7:0] tmp_276_fu_8673_p4;
wire   [7:0] tmp_221_fu_8726_p4;
wire   [7:0] tmp_219_fu_8712_p4;
wire   [7:0] tmp_226_fu_8770_p4;
wire   [7:0] trunc_ln674_52_fu_8790_p1;
wire   [7:0] xor_ln1545_152_fu_9238_p2;
wire   [7:0] xor_ln1545_150_fu_9232_p2;
wire   [7:0] tmp_223_fu_8746_p4;
wire   [7:0] trunc_ln674_49_fu_8688_p1;
wire   [7:0] tmp_225_fu_8760_p4;
wire   [7:0] tmp_230_fu_8804_p4;
wire   [7:0] xor_ln1545_155_fu_9256_p2;
wire   [7:0] xor_ln1545_153_fu_9250_p2;
wire   [7:0] trunc_ln674_50_fu_8722_p1;
wire   [7:0] tmp_218_fu_8702_p4;
wire   [7:0] tmp_227_fu_8780_p4;
wire   [7:0] tmp_229_fu_8794_p4;
wire   [7:0] xor_ln1545_158_fu_9274_p2;
wire   [7:0] xor_ln1545_156_fu_9268_p2;
wire   [7:0] tmp_222_fu_8736_p4;
wire   [7:0] tmp_217_fu_8692_p4;
wire   [7:0] trunc_ln674_51_fu_8756_p1;
wire   [7:0] tmp_231_fu_8814_p4;
wire   [7:0] xor_ln1545_160_fu_9292_p2;
wire   [7:0] xor_ln1545_159_fu_9286_p2;
wire   [7:0] tmp_237_fu_8862_p4;
wire   [7:0] tmp_235_fu_8848_p4;
wire   [7:0] tmp_242_fu_8906_p4;
wire   [7:0] trunc_ln674_56_fu_8926_p1;
wire   [7:0] xor_ln1545_164_fu_9310_p2;
wire   [7:0] xor_ln1545_162_fu_9304_p2;
wire   [7:0] tmp_239_fu_8882_p4;
wire   [7:0] trunc_ln674_53_fu_8824_p1;
wire   [7:0] tmp_241_fu_8896_p4;
wire   [7:0] tmp_246_fu_8940_p4;
wire   [7:0] xor_ln1545_167_fu_9328_p2;
wire   [7:0] xor_ln1545_165_fu_9322_p2;
wire   [7:0] trunc_ln674_54_fu_8858_p1;
wire   [7:0] tmp_234_fu_8838_p4;
wire   [7:0] tmp_243_fu_8916_p4;
wire   [7:0] tmp_245_fu_8930_p4;
wire   [7:0] xor_ln1545_170_fu_9346_p2;
wire   [7:0] xor_ln1545_168_fu_9340_p2;
wire   [7:0] tmp_238_fu_8872_p4;
wire   [7:0] tmp_233_fu_8828_p4;
wire   [7:0] trunc_ln674_55_fu_8892_p1;
wire   [7:0] tmp_247_fu_8950_p4;
wire   [7:0] xor_ln1545_173_fu_9364_p2;
wire   [7:0] xor_ln1545_171_fu_9358_p2;
wire   [7:0] tmp_253_fu_8998_p4;
wire   [7:0] tmp_251_fu_8984_p4;
wire   [7:0] tmp_258_fu_9042_p4;
wire   [7:0] trunc_ln674_60_fu_9062_p1;
wire   [7:0] xor_ln1545_176_fu_9382_p2;
wire   [7:0] xor_ln1545_174_fu_9376_p2;
wire   [7:0] tmp_255_fu_9018_p4;
wire   [7:0] trunc_ln674_57_fu_8960_p1;
wire   [7:0] tmp_257_fu_9032_p4;
wire   [7:0] tmp_262_fu_9076_p4;
wire   [7:0] xor_ln1545_179_fu_9400_p2;
wire   [7:0] xor_ln1545_177_fu_9394_p2;
wire   [7:0] trunc_ln674_58_fu_8994_p1;
wire   [7:0] tmp_250_fu_8974_p4;
wire   [7:0] tmp_259_fu_9052_p4;
wire   [7:0] tmp_261_fu_9066_p4;
wire   [7:0] xor_ln1545_181_fu_9418_p2;
wire   [7:0] xor_ln1545_180_fu_9412_p2;
wire   [7:0] tmp_254_fu_9008_p4;
wire   [7:0] tmp_249_fu_8964_p4;
wire   [7:0] trunc_ln674_59_fu_9028_p1;
wire   [7:0] tmp_263_fu_9086_p4;
wire   [7:0] xor_ln1545_185_fu_9436_p2;
wire   [7:0] xor_ln1545_183_fu_9430_p2;
wire   [7:0] tmp_269_fu_9134_p4;
wire   [7:0] tmp_267_fu_9120_p4;
wire   [7:0] tmp_274_fu_9178_p4;
wire   [7:0] trunc_ln674_64_fu_9198_p1;
wire   [7:0] xor_ln1545_188_fu_9454_p2;
wire   [7:0] xor_ln1545_186_fu_9448_p2;
wire   [7:0] tmp_271_fu_9154_p4;
wire   [7:0] trunc_ln674_61_fu_9096_p1;
wire   [7:0] tmp_273_fu_9168_p4;
wire   [7:0] tmp_278_fu_9212_p4;
wire   [7:0] xor_ln1545_190_fu_9472_p2;
wire   [7:0] xor_ln1545_189_fu_9466_p2;
wire   [7:0] trunc_ln674_62_fu_9130_p1;
wire   [7:0] tmp_266_fu_9110_p4;
wire   [7:0] tmp_275_fu_9188_p4;
wire   [7:0] tmp_277_fu_9202_p4;
wire   [7:0] xor_ln1545_193_fu_9490_p2;
wire   [7:0] xor_ln1545_192_fu_9484_p2;
wire   [7:0] tmp_270_fu_9144_p4;
wire   [7:0] tmp_265_fu_9100_p4;
wire   [7:0] trunc_ln674_63_fu_9164_p1;
wire   [7:0] tmp_279_fu_9222_p4;
wire   [7:0] xor_ln1545_197_fu_9508_p2;
wire   [7:0] xor_ln1545_195_fu_9502_p2;
wire   [7:0] xor_ln1545_151_fu_9244_p2;
wire   [7:0] tmp_1_V_3_fu_9478_p2;
wire   [7:0] tmp_2_1_V_3_fu_9424_p2;
wire   [7:0] xor_ln1545_172_fu_9370_p2;
wire   [7:0] xor_ln1545_163_fu_9316_p2;
wire   [7:0] xor_ln1545_154_fu_9262_p2;
wire   [7:0] tmp_2_2_V_3_fu_9496_p2;
wire   [7:0] xor_ln1545_184_fu_9442_p2;
wire   [7:0] xor_ln1545_175_fu_9388_p2;
wire   [7:0] xor_ln1545_166_fu_9334_p2;
wire   [7:0] xor_ln1545_157_fu_9280_p2;
wire   [7:0] xor_ln1545_196_fu_9514_p2;
wire   [7:0] xor_ln1545_187_fu_9460_p2;
wire   [7:0] xor_ln1545_178_fu_9406_p2;
wire   [7:0] xor_ln1545_169_fu_9352_p2;
wire   [7:0] tmp_3_V_3_fu_9298_p2;
wire   [127:0] p_Result_28_fu_9600_p17;
wire   [127:0] state_V_28_fu_9636_p2;
wire   [7:0] trunc_ln708_5_fu_9641_p1;
wire   [7:0] tmp_283_fu_9650_p4;
wire   [7:0] tmp_287_fu_9665_p4;
wire   [7:0] tmp_291_fu_9680_p4;
wire   [7:0] tmp_295_fu_9695_p4;
wire   [7:0] tmp_299_fu_9710_p4;
wire   [7:0] tmp_303_fu_9725_p4;
wire   [7:0] tmp_307_fu_9740_p4;
wire   [7:0] tmp_311_fu_9755_p4;
wire   [7:0] tmp_315_fu_9770_p4;
wire   [7:0] tmp_319_fu_9785_p4;
wire   [7:0] tmp_323_fu_9800_p4;
wire   [7:0] tmp_327_fu_9815_p4;
wire   [7:0] tmp_331_fu_9830_p4;
wire   [7:0] tmp_335_fu_9845_p4;
wire   [7:0] tmp_339_fu_9860_p4;
wire   [7:0] tmp_284_fu_9913_p4;
wire   [7:0] tmp_282_fu_9899_p4;
wire   [7:0] tmp_289_fu_9957_p4;
wire   [7:0] trunc_ln674_68_fu_9977_p1;
wire   [7:0] xor_ln1545_200_fu_10425_p2;
wire   [7:0] xor_ln1545_198_fu_10419_p2;
wire   [7:0] tmp_286_fu_9933_p4;
wire   [7:0] trunc_ln674_65_fu_9875_p1;
wire   [7:0] tmp_288_fu_9947_p4;
wire   [7:0] tmp_293_fu_9991_p4;
wire   [7:0] xor_ln1545_203_fu_10443_p2;
wire   [7:0] xor_ln1545_201_fu_10437_p2;
wire   [7:0] trunc_ln674_66_fu_9909_p1;
wire   [7:0] tmp_281_fu_9889_p4;
wire   [7:0] tmp_290_fu_9967_p4;
wire   [7:0] tmp_292_fu_9981_p4;
wire   [7:0] xor_ln1545_206_fu_10461_p2;
wire   [7:0] xor_ln1545_204_fu_10455_p2;
wire   [7:0] tmp_285_fu_9923_p4;
wire   [7:0] tmp_280_fu_9879_p4;
wire   [7:0] trunc_ln674_67_fu_9943_p1;
wire   [7:0] tmp_294_fu_10001_p4;
wire   [7:0] xor_ln1545_208_fu_10479_p2;
wire   [7:0] xor_ln1545_207_fu_10473_p2;
wire   [7:0] tmp_300_fu_10049_p4;
wire   [7:0] tmp_298_fu_10035_p4;
wire   [7:0] tmp_305_fu_10093_p4;
wire   [7:0] trunc_ln674_72_fu_10113_p1;
wire   [7:0] xor_ln1545_212_fu_10497_p2;
wire   [7:0] xor_ln1545_210_fu_10491_p2;
wire   [7:0] tmp_302_fu_10069_p4;
wire   [7:0] trunc_ln674_69_fu_10011_p1;
wire   [7:0] tmp_304_fu_10083_p4;
wire   [7:0] tmp_309_fu_10127_p4;
wire   [7:0] xor_ln1545_215_fu_10515_p2;
wire   [7:0] xor_ln1545_213_fu_10509_p2;
wire   [7:0] trunc_ln674_70_fu_10045_p1;
wire   [7:0] tmp_297_fu_10025_p4;
wire   [7:0] tmp_306_fu_10103_p4;
wire   [7:0] tmp_308_fu_10117_p4;
wire   [7:0] xor_ln1545_218_fu_10533_p2;
wire   [7:0] xor_ln1545_216_fu_10527_p2;
wire   [7:0] tmp_301_fu_10059_p4;
wire   [7:0] tmp_296_fu_10015_p4;
wire   [7:0] trunc_ln674_71_fu_10079_p1;
wire   [7:0] tmp_310_fu_10137_p4;
wire   [7:0] xor_ln1545_221_fu_10551_p2;
wire   [7:0] xor_ln1545_219_fu_10545_p2;
wire   [7:0] tmp_316_fu_10185_p4;
wire   [7:0] tmp_314_fu_10171_p4;
wire   [7:0] tmp_321_fu_10229_p4;
wire   [7:0] trunc_ln674_76_fu_10249_p1;
wire   [7:0] xor_ln1545_224_fu_10569_p2;
wire   [7:0] xor_ln1545_222_fu_10563_p2;
wire   [7:0] tmp_318_fu_10205_p4;
wire   [7:0] trunc_ln674_73_fu_10147_p1;
wire   [7:0] tmp_320_fu_10219_p4;
wire   [7:0] tmp_325_fu_10263_p4;
wire   [7:0] xor_ln1545_227_fu_10587_p2;
wire   [7:0] xor_ln1545_225_fu_10581_p2;
wire   [7:0] trunc_ln674_74_fu_10181_p1;
wire   [7:0] tmp_313_fu_10161_p4;
wire   [7:0] tmp_322_fu_10239_p4;
wire   [7:0] tmp_324_fu_10253_p4;
wire   [7:0] xor_ln1545_229_fu_10605_p2;
wire   [7:0] xor_ln1545_228_fu_10599_p2;
wire   [7:0] tmp_317_fu_10195_p4;
wire   [7:0] tmp_312_fu_10151_p4;
wire   [7:0] trunc_ln674_75_fu_10215_p1;
wire   [7:0] tmp_326_fu_10273_p4;
wire   [7:0] xor_ln1545_233_fu_10623_p2;
wire   [7:0] xor_ln1545_231_fu_10617_p2;
wire   [7:0] tmp_332_fu_10321_p4;
wire   [7:0] tmp_330_fu_10307_p4;
wire   [7:0] tmp_337_fu_10365_p4;
wire   [7:0] trunc_ln674_80_fu_10385_p1;
wire   [7:0] xor_ln1545_236_fu_10641_p2;
wire   [7:0] xor_ln1545_234_fu_10635_p2;
wire   [7:0] tmp_334_fu_10341_p4;
wire   [7:0] trunc_ln674_77_fu_10283_p1;
wire   [7:0] tmp_336_fu_10355_p4;
wire   [7:0] tmp_341_fu_10399_p4;
wire   [7:0] xor_ln1545_238_fu_10659_p2;
wire   [7:0] xor_ln1545_237_fu_10653_p2;
wire   [7:0] trunc_ln674_78_fu_10317_p1;
wire   [7:0] tmp_329_fu_10297_p4;
wire   [7:0] tmp_338_fu_10375_p4;
wire   [7:0] tmp_340_fu_10389_p4;
wire   [7:0] xor_ln1545_241_fu_10677_p2;
wire   [7:0] xor_ln1545_240_fu_10671_p2;
wire   [7:0] tmp_333_fu_10331_p4;
wire   [7:0] tmp_328_fu_10287_p4;
wire   [7:0] trunc_ln674_79_fu_10351_p1;
wire   [7:0] tmp_342_fu_10409_p4;
wire   [7:0] xor_ln1545_245_fu_10695_p2;
wire   [7:0] xor_ln1545_243_fu_10689_p2;
wire   [7:0] xor_ln1545_199_fu_10431_p2;
wire   [7:0] tmp_1_V_4_fu_10665_p2;
wire   [7:0] tmp_2_1_V_4_fu_10611_p2;
wire   [7:0] xor_ln1545_220_fu_10557_p2;
wire   [7:0] xor_ln1545_211_fu_10503_p2;
wire   [7:0] xor_ln1545_202_fu_10449_p2;
wire   [7:0] tmp_2_2_V_4_fu_10683_p2;
wire   [7:0] xor_ln1545_232_fu_10629_p2;
wire   [7:0] xor_ln1545_223_fu_10575_p2;
wire   [7:0] xor_ln1545_214_fu_10521_p2;
wire   [7:0] xor_ln1545_205_fu_10467_p2;
wire   [7:0] xor_ln1545_244_fu_10701_p2;
wire   [7:0] xor_ln1545_235_fu_10647_p2;
wire   [7:0] xor_ln1545_226_fu_10593_p2;
wire   [7:0] xor_ln1545_217_fu_10539_p2;
wire   [7:0] tmp_3_V_4_fu_10485_p2;
wire   [127:0] p_Result_29_fu_10787_p17;
wire   [127:0] state_V_29_fu_10823_p2;
wire   [7:0] trunc_ln708_6_fu_10828_p1;
wire   [7:0] tmp_346_fu_10837_p4;
wire   [7:0] tmp_350_fu_10852_p4;
wire   [7:0] tmp_354_fu_10867_p4;
wire   [7:0] tmp_358_fu_10882_p4;
wire   [7:0] tmp_362_fu_10897_p4;
wire   [7:0] tmp_366_fu_10912_p4;
wire   [7:0] tmp_370_fu_10927_p4;
wire   [7:0] tmp_374_fu_10942_p4;
wire   [7:0] tmp_378_fu_10957_p4;
wire   [7:0] tmp_382_fu_10972_p4;
wire   [7:0] tmp_386_fu_10987_p4;
wire   [7:0] tmp_390_fu_11002_p4;
wire   [7:0] tmp_394_fu_11017_p4;
wire   [7:0] tmp_398_fu_11032_p4;
wire   [7:0] tmp_402_fu_11047_p4;
wire   [7:0] tmp_347_fu_11100_p4;
wire   [7:0] tmp_345_fu_11086_p4;
wire   [7:0] tmp_352_fu_11144_p4;
wire   [7:0] trunc_ln674_84_fu_11164_p1;
wire   [7:0] xor_ln1545_248_fu_11612_p2;
wire   [7:0] xor_ln1545_246_fu_11606_p2;
wire   [7:0] tmp_349_fu_11120_p4;
wire   [7:0] trunc_ln674_81_fu_11062_p1;
wire   [7:0] tmp_351_fu_11134_p4;
wire   [7:0] tmp_356_fu_11178_p4;
wire   [7:0] xor_ln1545_251_fu_11630_p2;
wire   [7:0] xor_ln1545_249_fu_11624_p2;
wire   [7:0] trunc_ln674_82_fu_11096_p1;
wire   [7:0] tmp_344_fu_11076_p4;
wire   [7:0] tmp_353_fu_11154_p4;
wire   [7:0] tmp_355_fu_11168_p4;
wire   [7:0] xor_ln1545_254_fu_11648_p2;
wire   [7:0] xor_ln1545_252_fu_11642_p2;
wire   [7:0] tmp_348_fu_11110_p4;
wire   [7:0] tmp_343_fu_11066_p4;
wire   [7:0] trunc_ln674_83_fu_11130_p1;
wire   [7:0] tmp_357_fu_11188_p4;
wire   [7:0] xor_ln1545_256_fu_11666_p2;
wire   [7:0] xor_ln1545_255_fu_11660_p2;
wire   [7:0] tmp_363_fu_11236_p4;
wire   [7:0] tmp_361_fu_11222_p4;
wire   [7:0] tmp_368_fu_11280_p4;
wire   [7:0] trunc_ln674_88_fu_11300_p1;
wire   [7:0] xor_ln1545_260_fu_11684_p2;
wire   [7:0] xor_ln1545_258_fu_11678_p2;
wire   [7:0] tmp_365_fu_11256_p4;
wire   [7:0] trunc_ln674_85_fu_11198_p1;
wire   [7:0] tmp_367_fu_11270_p4;
wire   [7:0] tmp_372_fu_11314_p4;
wire   [7:0] xor_ln1545_263_fu_11702_p2;
wire   [7:0] xor_ln1545_261_fu_11696_p2;
wire   [7:0] trunc_ln674_86_fu_11232_p1;
wire   [7:0] tmp_360_fu_11212_p4;
wire   [7:0] tmp_369_fu_11290_p4;
wire   [7:0] tmp_371_fu_11304_p4;
wire   [7:0] xor_ln1545_266_fu_11720_p2;
wire   [7:0] xor_ln1545_264_fu_11714_p2;
wire   [7:0] tmp_364_fu_11246_p4;
wire   [7:0] tmp_359_fu_11202_p4;
wire   [7:0] trunc_ln674_87_fu_11266_p1;
wire   [7:0] tmp_373_fu_11324_p4;
wire   [7:0] xor_ln1545_269_fu_11738_p2;
wire   [7:0] xor_ln1545_267_fu_11732_p2;
wire   [7:0] tmp_379_fu_11372_p4;
wire   [7:0] tmp_377_fu_11358_p4;
wire   [7:0] tmp_384_fu_11416_p4;
wire   [7:0] trunc_ln674_92_fu_11436_p1;
wire   [7:0] xor_ln1545_272_fu_11756_p2;
wire   [7:0] xor_ln1545_270_fu_11750_p2;
wire   [7:0] tmp_381_fu_11392_p4;
wire   [7:0] trunc_ln674_89_fu_11334_p1;
wire   [7:0] tmp_383_fu_11406_p4;
wire   [7:0] tmp_388_fu_11450_p4;
wire   [7:0] xor_ln1545_275_fu_11774_p2;
wire   [7:0] xor_ln1545_273_fu_11768_p2;
wire   [7:0] trunc_ln674_90_fu_11368_p1;
wire   [7:0] tmp_376_fu_11348_p4;
wire   [7:0] tmp_385_fu_11426_p4;
wire   [7:0] tmp_387_fu_11440_p4;
wire   [7:0] xor_ln1545_277_fu_11792_p2;
wire   [7:0] xor_ln1545_276_fu_11786_p2;
wire   [7:0] tmp_380_fu_11382_p4;
wire   [7:0] tmp_375_fu_11338_p4;
wire   [7:0] trunc_ln674_91_fu_11402_p1;
wire   [7:0] tmp_389_fu_11460_p4;
wire   [7:0] xor_ln1545_281_fu_11810_p2;
wire   [7:0] xor_ln1545_279_fu_11804_p2;
wire   [7:0] tmp_395_fu_11508_p4;
wire   [7:0] tmp_393_fu_11494_p4;
wire   [7:0] tmp_400_fu_11552_p4;
wire   [7:0] trunc_ln674_96_fu_11572_p1;
wire   [7:0] xor_ln1545_284_fu_11828_p2;
wire   [7:0] xor_ln1545_282_fu_11822_p2;
wire   [7:0] tmp_397_fu_11528_p4;
wire   [7:0] trunc_ln674_93_fu_11470_p1;
wire   [7:0] tmp_399_fu_11542_p4;
wire   [7:0] tmp_404_fu_11586_p4;
wire   [7:0] xor_ln1545_286_fu_11846_p2;
wire   [7:0] xor_ln1545_285_fu_11840_p2;
wire   [7:0] trunc_ln674_94_fu_11504_p1;
wire   [7:0] tmp_392_fu_11484_p4;
wire   [7:0] tmp_401_fu_11562_p4;
wire   [7:0] tmp_403_fu_11576_p4;
wire   [7:0] xor_ln1545_289_fu_11864_p2;
wire   [7:0] xor_ln1545_288_fu_11858_p2;
wire   [7:0] tmp_396_fu_11518_p4;
wire   [7:0] tmp_391_fu_11474_p4;
wire   [7:0] trunc_ln674_95_fu_11538_p1;
wire   [7:0] tmp_405_fu_11596_p4;
wire   [7:0] xor_ln1545_293_fu_11882_p2;
wire   [7:0] xor_ln1545_291_fu_11876_p2;
wire   [7:0] xor_ln1545_247_fu_11618_p2;
wire   [7:0] tmp_1_V_5_fu_11852_p2;
wire   [7:0] tmp_2_1_V_5_fu_11798_p2;
wire   [7:0] xor_ln1545_268_fu_11744_p2;
wire   [7:0] xor_ln1545_259_fu_11690_p2;
wire   [7:0] xor_ln1545_250_fu_11636_p2;
wire   [7:0] tmp_2_2_V_5_fu_11870_p2;
wire   [7:0] xor_ln1545_280_fu_11816_p2;
wire   [7:0] xor_ln1545_271_fu_11762_p2;
wire   [7:0] xor_ln1545_262_fu_11708_p2;
wire   [7:0] xor_ln1545_253_fu_11654_p2;
wire   [7:0] xor_ln1545_292_fu_11888_p2;
wire   [7:0] xor_ln1545_283_fu_11834_p2;
wire   [7:0] xor_ln1545_274_fu_11780_p2;
wire   [7:0] xor_ln1545_265_fu_11726_p2;
wire   [7:0] tmp_3_V_5_fu_11672_p2;
wire   [127:0] p_Result_30_fu_11974_p17;
wire   [127:0] state_V_fu_12010_p2;
wire   [7:0] trunc_ln708_7_fu_12015_p1;
wire   [7:0] tmp_409_fu_12024_p4;
wire   [7:0] tmp_413_fu_12039_p4;
wire   [7:0] tmp_417_fu_12054_p4;
wire   [7:0] tmp_421_fu_12069_p4;
wire   [7:0] tmp_425_fu_12084_p4;
wire   [7:0] tmp_429_fu_12099_p4;
wire   [7:0] tmp_433_fu_12114_p4;
wire   [7:0] tmp_437_fu_12129_p4;
wire   [7:0] tmp_441_fu_12144_p4;
wire   [7:0] tmp_445_fu_12159_p4;
wire   [7:0] tmp_449_fu_12174_p4;
wire   [7:0] tmp_453_fu_12189_p4;
wire   [7:0] tmp_457_fu_12204_p4;
wire   [7:0] tmp_461_fu_12219_p4;
wire   [7:0] tmp_465_fu_12234_p4;
wire   [7:0] tmp_410_fu_12287_p4;
wire   [7:0] tmp_408_fu_12273_p4;
wire   [7:0] tmp_415_fu_12331_p4;
wire   [7:0] trunc_ln674_100_fu_12351_p1;
wire   [7:0] xor_ln1545_296_fu_12799_p2;
wire   [7:0] xor_ln1545_294_fu_12793_p2;
wire   [7:0] tmp_412_fu_12307_p4;
wire   [7:0] trunc_ln674_97_fu_12249_p1;
wire   [7:0] tmp_414_fu_12321_p4;
wire   [7:0] tmp_419_fu_12365_p4;
wire   [7:0] xor_ln1545_299_fu_12817_p2;
wire   [7:0] xor_ln1545_297_fu_12811_p2;
wire   [7:0] trunc_ln674_98_fu_12283_p1;
wire   [7:0] tmp_407_fu_12263_p4;
wire   [7:0] tmp_416_fu_12341_p4;
wire   [7:0] tmp_418_fu_12355_p4;
wire   [7:0] xor_ln1545_302_fu_12835_p2;
wire   [7:0] xor_ln1545_300_fu_12829_p2;
wire   [7:0] tmp_411_fu_12297_p4;
wire   [7:0] tmp_406_fu_12253_p4;
wire   [7:0] trunc_ln674_99_fu_12317_p1;
wire   [7:0] tmp_420_fu_12375_p4;
wire   [7:0] xor_ln1545_304_fu_12853_p2;
wire   [7:0] xor_ln1545_303_fu_12847_p2;
wire   [7:0] tmp_426_fu_12423_p4;
wire   [7:0] tmp_424_fu_12409_p4;
wire   [7:0] tmp_431_fu_12467_p4;
wire   [7:0] trunc_ln674_104_fu_12487_p1;
wire   [7:0] xor_ln1545_308_fu_12871_p2;
wire   [7:0] xor_ln1545_306_fu_12865_p2;
wire   [7:0] tmp_428_fu_12443_p4;
wire   [7:0] trunc_ln674_101_fu_12385_p1;
wire   [7:0] tmp_430_fu_12457_p4;
wire   [7:0] tmp_435_fu_12501_p4;
wire   [7:0] xor_ln1545_311_fu_12889_p2;
wire   [7:0] xor_ln1545_309_fu_12883_p2;
wire   [7:0] trunc_ln674_102_fu_12419_p1;
wire   [7:0] tmp_423_fu_12399_p4;
wire   [7:0] tmp_432_fu_12477_p4;
wire   [7:0] tmp_434_fu_12491_p4;
wire   [7:0] xor_ln1545_314_fu_12907_p2;
wire   [7:0] xor_ln1545_312_fu_12901_p2;
wire   [7:0] tmp_427_fu_12433_p4;
wire   [7:0] tmp_422_fu_12389_p4;
wire   [7:0] trunc_ln674_103_fu_12453_p1;
wire   [7:0] tmp_436_fu_12511_p4;
wire   [7:0] xor_ln1545_317_fu_12925_p2;
wire   [7:0] xor_ln1545_315_fu_12919_p2;
wire   [7:0] tmp_442_fu_12559_p4;
wire   [7:0] tmp_440_fu_12545_p4;
wire   [7:0] tmp_447_fu_12603_p4;
wire   [7:0] trunc_ln674_108_fu_12623_p1;
wire   [7:0] xor_ln1545_320_fu_12943_p2;
wire   [7:0] xor_ln1545_318_fu_12937_p2;
wire   [7:0] tmp_444_fu_12579_p4;
wire   [7:0] trunc_ln674_105_fu_12521_p1;
wire   [7:0] tmp_446_fu_12593_p4;
wire   [7:0] tmp_451_fu_12637_p4;
wire   [7:0] xor_ln1545_323_fu_12961_p2;
wire   [7:0] xor_ln1545_321_fu_12955_p2;
wire   [7:0] trunc_ln674_106_fu_12555_p1;
wire   [7:0] tmp_439_fu_12535_p4;
wire   [7:0] tmp_448_fu_12613_p4;
wire   [7:0] tmp_450_fu_12627_p4;
wire   [7:0] xor_ln1545_325_fu_12979_p2;
wire   [7:0] xor_ln1545_324_fu_12973_p2;
wire   [7:0] tmp_443_fu_12569_p4;
wire   [7:0] tmp_438_fu_12525_p4;
wire   [7:0] trunc_ln674_107_fu_12589_p1;
wire   [7:0] tmp_452_fu_12647_p4;
wire   [7:0] xor_ln1545_329_fu_12997_p2;
wire   [7:0] xor_ln1545_327_fu_12991_p2;
wire   [7:0] tmp_458_fu_12695_p4;
wire   [7:0] tmp_456_fu_12681_p4;
wire   [7:0] tmp_463_fu_12739_p4;
wire   [7:0] trunc_ln674_112_fu_12759_p1;
wire   [7:0] xor_ln1545_332_fu_13015_p2;
wire   [7:0] xor_ln1545_330_fu_13009_p2;
wire   [7:0] tmp_460_fu_12715_p4;
wire   [7:0] trunc_ln674_109_fu_12657_p1;
wire   [7:0] tmp_462_fu_12729_p4;
wire   [7:0] tmp_467_fu_12773_p4;
wire   [7:0] xor_ln1545_334_fu_13033_p2;
wire   [7:0] xor_ln1545_333_fu_13027_p2;
wire   [7:0] trunc_ln674_110_fu_12691_p1;
wire   [7:0] tmp_455_fu_12671_p4;
wire   [7:0] tmp_464_fu_12749_p4;
wire   [7:0] tmp_466_fu_12763_p4;
wire   [7:0] xor_ln1545_337_fu_13051_p2;
wire   [7:0] xor_ln1545_336_fu_13045_p2;
wire   [7:0] tmp_459_fu_12705_p4;
wire   [7:0] tmp_454_fu_12661_p4;
wire   [7:0] trunc_ln674_111_fu_12725_p1;
wire   [7:0] tmp_468_fu_12783_p4;
wire   [7:0] xor_ln1545_341_fu_13069_p2;
wire   [7:0] xor_ln1545_339_fu_13063_p2;
wire   [7:0] xor_ln1545_295_fu_12805_p2;
wire   [7:0] tmp_1_V_6_fu_13039_p2;
wire   [7:0] tmp_2_1_V_6_fu_12985_p2;
wire   [7:0] xor_ln1545_316_fu_12931_p2;
wire   [7:0] xor_ln1545_307_fu_12877_p2;
wire   [7:0] xor_ln1545_298_fu_12823_p2;
wire   [7:0] tmp_2_2_V_6_fu_13057_p2;
wire   [7:0] xor_ln1545_328_fu_13003_p2;
wire   [7:0] xor_ln1545_319_fu_12949_p2;
wire   [7:0] xor_ln1545_310_fu_12895_p2;
wire   [7:0] xor_ln1545_301_fu_12841_p2;
wire   [7:0] xor_ln1545_340_fu_13075_p2;
wire   [7:0] xor_ln1545_331_fu_13021_p2;
wire   [7:0] xor_ln1545_322_fu_12967_p2;
wire   [7:0] xor_ln1545_313_fu_12913_p2;
wire   [7:0] tmp_3_V_6_fu_12859_p2;
wire   [127:0] p_Result_31_fu_13161_p17;
wire   [127:0] state_V_30_fu_13197_p2;
wire   [7:0] trunc_ln708_8_fu_13202_p1;
wire   [7:0] tmp_472_fu_13211_p4;
wire   [7:0] tmp_476_fu_13226_p4;
wire   [7:0] tmp_480_fu_13241_p4;
wire   [7:0] tmp_484_fu_13256_p4;
wire   [7:0] tmp_488_fu_13271_p4;
wire   [7:0] tmp_492_fu_13286_p4;
wire   [7:0] tmp_496_fu_13301_p4;
wire   [7:0] tmp_500_fu_13316_p4;
wire   [7:0] tmp_504_fu_13331_p4;
wire   [7:0] tmp_508_fu_13346_p4;
wire   [7:0] tmp_512_fu_13361_p4;
wire   [7:0] tmp_516_fu_13376_p4;
wire   [7:0] tmp_520_fu_13391_p4;
wire   [7:0] tmp_524_fu_13406_p4;
wire   [7:0] tmp_528_fu_13421_p4;
wire   [7:0] tmp_473_fu_13474_p4;
wire   [7:0] tmp_471_fu_13460_p4;
wire   [7:0] tmp_478_fu_13518_p4;
wire   [7:0] trunc_ln674_116_fu_13538_p1;
wire   [7:0] xor_ln1545_344_fu_13986_p2;
wire   [7:0] xor_ln1545_342_fu_13980_p2;
wire   [7:0] tmp_475_fu_13494_p4;
wire   [7:0] trunc_ln674_113_fu_13436_p1;
wire   [7:0] tmp_477_fu_13508_p4;
wire   [7:0] tmp_482_fu_13552_p4;
wire   [7:0] xor_ln1545_347_fu_14004_p2;
wire   [7:0] xor_ln1545_345_fu_13998_p2;
wire   [7:0] trunc_ln674_114_fu_13470_p1;
wire   [7:0] tmp_470_fu_13450_p4;
wire   [7:0] tmp_479_fu_13528_p4;
wire   [7:0] tmp_481_fu_13542_p4;
wire   [7:0] xor_ln1545_350_fu_14022_p2;
wire   [7:0] xor_ln1545_348_fu_14016_p2;
wire   [7:0] tmp_474_fu_13484_p4;
wire   [7:0] tmp_469_fu_13440_p4;
wire   [7:0] trunc_ln674_115_fu_13504_p1;
wire   [7:0] tmp_483_fu_13562_p4;
wire   [7:0] xor_ln1545_352_fu_14040_p2;
wire   [7:0] xor_ln1545_351_fu_14034_p2;
wire   [7:0] tmp_489_fu_13610_p4;
wire   [7:0] tmp_487_fu_13596_p4;
wire   [7:0] tmp_494_fu_13654_p4;
wire   [7:0] trunc_ln674_120_fu_13674_p1;
wire   [7:0] xor_ln1545_356_fu_14058_p2;
wire   [7:0] xor_ln1545_354_fu_14052_p2;
wire   [7:0] tmp_491_fu_13630_p4;
wire   [7:0] trunc_ln674_117_fu_13572_p1;
wire   [7:0] tmp_493_fu_13644_p4;
wire   [7:0] tmp_498_fu_13688_p4;
wire   [7:0] xor_ln1545_359_fu_14076_p2;
wire   [7:0] xor_ln1545_357_fu_14070_p2;
wire   [7:0] trunc_ln674_118_fu_13606_p1;
wire   [7:0] tmp_486_fu_13586_p4;
wire   [7:0] tmp_495_fu_13664_p4;
wire   [7:0] tmp_497_fu_13678_p4;
wire   [7:0] xor_ln1545_362_fu_14094_p2;
wire   [7:0] xor_ln1545_360_fu_14088_p2;
wire   [7:0] tmp_490_fu_13620_p4;
wire   [7:0] tmp_485_fu_13576_p4;
wire   [7:0] trunc_ln674_119_fu_13640_p1;
wire   [7:0] tmp_499_fu_13698_p4;
wire   [7:0] xor_ln1545_365_fu_14112_p2;
wire   [7:0] xor_ln1545_363_fu_14106_p2;
wire   [7:0] tmp_505_fu_13746_p4;
wire   [7:0] tmp_503_fu_13732_p4;
wire   [7:0] tmp_510_fu_13790_p4;
wire   [7:0] trunc_ln674_124_fu_13810_p1;
wire   [7:0] xor_ln1545_368_fu_14130_p2;
wire   [7:0] xor_ln1545_366_fu_14124_p2;
wire   [7:0] tmp_507_fu_13766_p4;
wire   [7:0] trunc_ln674_121_fu_13708_p1;
wire   [7:0] tmp_509_fu_13780_p4;
wire   [7:0] tmp_514_fu_13824_p4;
wire   [7:0] xor_ln1545_371_fu_14148_p2;
wire   [7:0] xor_ln1545_369_fu_14142_p2;
wire   [7:0] trunc_ln674_122_fu_13742_p1;
wire   [7:0] tmp_502_fu_13722_p4;
wire   [7:0] tmp_511_fu_13800_p4;
wire   [7:0] tmp_513_fu_13814_p4;
wire   [7:0] xor_ln1545_373_fu_14166_p2;
wire   [7:0] xor_ln1545_372_fu_14160_p2;
wire   [7:0] tmp_506_fu_13756_p4;
wire   [7:0] tmp_501_fu_13712_p4;
wire   [7:0] trunc_ln674_123_fu_13776_p1;
wire   [7:0] tmp_515_fu_13834_p4;
wire   [7:0] xor_ln1545_377_fu_14184_p2;
wire   [7:0] xor_ln1545_375_fu_14178_p2;
wire   [7:0] tmp_521_fu_13882_p4;
wire   [7:0] tmp_519_fu_13868_p4;
wire   [7:0] tmp_526_fu_13926_p4;
wire   [7:0] trunc_ln674_128_fu_13946_p1;
wire   [7:0] xor_ln1545_380_fu_14202_p2;
wire   [7:0] xor_ln1545_378_fu_14196_p2;
wire   [7:0] tmp_523_fu_13902_p4;
wire   [7:0] trunc_ln674_125_fu_13844_p1;
wire   [7:0] tmp_525_fu_13916_p4;
wire   [7:0] tmp_530_fu_13960_p4;
wire   [7:0] xor_ln1545_382_fu_14220_p2;
wire   [7:0] xor_ln1545_381_fu_14214_p2;
wire   [7:0] trunc_ln674_126_fu_13878_p1;
wire   [7:0] tmp_518_fu_13858_p4;
wire   [7:0] tmp_527_fu_13936_p4;
wire   [7:0] tmp_529_fu_13950_p4;
wire   [7:0] xor_ln1545_385_fu_14238_p2;
wire   [7:0] xor_ln1545_384_fu_14232_p2;
wire   [7:0] tmp_522_fu_13892_p4;
wire   [7:0] tmp_517_fu_13848_p4;
wire   [7:0] trunc_ln674_127_fu_13912_p1;
wire   [7:0] tmp_531_fu_13970_p4;
wire   [7:0] xor_ln1545_389_fu_14256_p2;
wire   [7:0] xor_ln1545_387_fu_14250_p2;
wire   [7:0] xor_ln1545_343_fu_13992_p2;
wire   [7:0] tmp_1_V_7_fu_14226_p2;
wire   [7:0] tmp_2_1_V_7_fu_14172_p2;
wire   [7:0] xor_ln1545_364_fu_14118_p2;
wire   [7:0] xor_ln1545_355_fu_14064_p2;
wire   [7:0] xor_ln1545_346_fu_14010_p2;
wire   [7:0] tmp_2_2_V_7_fu_14244_p2;
wire   [7:0] xor_ln1545_376_fu_14190_p2;
wire   [7:0] xor_ln1545_367_fu_14136_p2;
wire   [7:0] xor_ln1545_358_fu_14082_p2;
wire   [7:0] xor_ln1545_349_fu_14028_p2;
wire   [7:0] xor_ln1545_388_fu_14262_p2;
wire   [7:0] xor_ln1545_379_fu_14208_p2;
wire   [7:0] xor_ln1545_370_fu_14154_p2;
wire   [7:0] xor_ln1545_361_fu_14100_p2;
wire   [7:0] tmp_3_V_7_fu_14046_p2;
wire   [127:0] p_Result_32_fu_14348_p17;
wire   [127:0] state_V_31_fu_14384_p2;
wire   [7:0] trunc_ln708_9_fu_14389_p1;
wire   [7:0] tmp_535_fu_14398_p4;
wire   [7:0] tmp_539_fu_14413_p4;
wire   [7:0] tmp_543_fu_14428_p4;
wire   [7:0] tmp_547_fu_14443_p4;
wire   [7:0] tmp_551_fu_14458_p4;
wire   [7:0] tmp_555_fu_14473_p4;
wire   [7:0] tmp_559_fu_14488_p4;
wire   [7:0] tmp_563_fu_14503_p4;
wire   [7:0] tmp_567_fu_14518_p4;
wire   [7:0] tmp_571_fu_14533_p4;
wire   [7:0] tmp_575_fu_14548_p4;
wire   [7:0] tmp_579_fu_14563_p4;
wire   [7:0] tmp_583_fu_14578_p4;
wire   [7:0] tmp_587_fu_14593_p4;
wire   [7:0] tmp_591_fu_14608_p4;
wire   [7:0] tmp_536_fu_14661_p4;
wire   [7:0] tmp_534_fu_14647_p4;
wire   [7:0] tmp_541_fu_14705_p4;
wire   [7:0] trunc_ln674_132_fu_14725_p1;
wire   [7:0] xor_ln1545_392_fu_15173_p2;
wire   [7:0] xor_ln1545_390_fu_15167_p2;
wire   [7:0] tmp_538_fu_14681_p4;
wire   [7:0] trunc_ln674_129_fu_14623_p1;
wire   [7:0] tmp_540_fu_14695_p4;
wire   [7:0] tmp_545_fu_14739_p4;
wire   [7:0] xor_ln1545_395_fu_15191_p2;
wire   [7:0] xor_ln1545_393_fu_15185_p2;
wire   [7:0] trunc_ln674_130_fu_14657_p1;
wire   [7:0] tmp_533_fu_14637_p4;
wire   [7:0] tmp_542_fu_14715_p4;
wire   [7:0] tmp_544_fu_14729_p4;
wire   [7:0] xor_ln1545_398_fu_15209_p2;
wire   [7:0] xor_ln1545_396_fu_15203_p2;
wire   [7:0] tmp_537_fu_14671_p4;
wire   [7:0] tmp_532_fu_14627_p4;
wire   [7:0] trunc_ln674_131_fu_14691_p1;
wire   [7:0] tmp_546_fu_14749_p4;
wire   [7:0] xor_ln1545_400_fu_15227_p2;
wire   [7:0] xor_ln1545_399_fu_15221_p2;
wire   [7:0] tmp_552_fu_14797_p4;
wire   [7:0] tmp_550_fu_14783_p4;
wire   [7:0] tmp_557_fu_14841_p4;
wire   [7:0] trunc_ln674_136_fu_14861_p1;
wire   [7:0] xor_ln1545_404_fu_15245_p2;
wire   [7:0] xor_ln1545_402_fu_15239_p2;
wire   [7:0] tmp_554_fu_14817_p4;
wire   [7:0] trunc_ln674_133_fu_14759_p1;
wire   [7:0] tmp_556_fu_14831_p4;
wire   [7:0] tmp_561_fu_14875_p4;
wire   [7:0] xor_ln1545_407_fu_15263_p2;
wire   [7:0] xor_ln1545_405_fu_15257_p2;
wire   [7:0] trunc_ln674_134_fu_14793_p1;
wire   [7:0] tmp_549_fu_14773_p4;
wire   [7:0] tmp_558_fu_14851_p4;
wire   [7:0] tmp_560_fu_14865_p4;
wire   [7:0] xor_ln1545_410_fu_15281_p2;
wire   [7:0] xor_ln1545_408_fu_15275_p2;
wire   [7:0] tmp_553_fu_14807_p4;
wire   [7:0] tmp_548_fu_14763_p4;
wire   [7:0] trunc_ln674_135_fu_14827_p1;
wire   [7:0] tmp_562_fu_14885_p4;
wire   [7:0] xor_ln1545_413_fu_15299_p2;
wire   [7:0] xor_ln1545_411_fu_15293_p2;
wire   [7:0] tmp_568_fu_14933_p4;
wire   [7:0] tmp_566_fu_14919_p4;
wire   [7:0] tmp_573_fu_14977_p4;
wire   [7:0] trunc_ln674_140_fu_14997_p1;
wire   [7:0] xor_ln1545_416_fu_15317_p2;
wire   [7:0] xor_ln1545_414_fu_15311_p2;
wire   [7:0] tmp_570_fu_14953_p4;
wire   [7:0] trunc_ln674_137_fu_14895_p1;
wire   [7:0] tmp_572_fu_14967_p4;
wire   [7:0] tmp_577_fu_15011_p4;
wire   [7:0] xor_ln1545_419_fu_15335_p2;
wire   [7:0] xor_ln1545_417_fu_15329_p2;
wire   [7:0] trunc_ln674_138_fu_14929_p1;
wire   [7:0] tmp_565_fu_14909_p4;
wire   [7:0] tmp_574_fu_14987_p4;
wire   [7:0] tmp_576_fu_15001_p4;
wire   [7:0] xor_ln1545_421_fu_15353_p2;
wire   [7:0] xor_ln1545_420_fu_15347_p2;
wire   [7:0] tmp_569_fu_14943_p4;
wire   [7:0] tmp_564_fu_14899_p4;
wire   [7:0] trunc_ln674_139_fu_14963_p1;
wire   [7:0] tmp_578_fu_15021_p4;
wire   [7:0] xor_ln1545_425_fu_15371_p2;
wire   [7:0] xor_ln1545_423_fu_15365_p2;
wire   [7:0] tmp_584_fu_15069_p4;
wire   [7:0] tmp_582_fu_15055_p4;
wire   [7:0] tmp_589_fu_15113_p4;
wire   [7:0] trunc_ln674_144_fu_15133_p1;
wire   [7:0] xor_ln1545_428_fu_15389_p2;
wire   [7:0] xor_ln1545_426_fu_15383_p2;
wire   [7:0] tmp_586_fu_15089_p4;
wire   [7:0] trunc_ln674_141_fu_15031_p1;
wire   [7:0] tmp_588_fu_15103_p4;
wire   [7:0] tmp_593_fu_15147_p4;
wire   [7:0] xor_ln1545_430_fu_15407_p2;
wire   [7:0] xor_ln1545_429_fu_15401_p2;
wire   [7:0] trunc_ln674_142_fu_15065_p1;
wire   [7:0] tmp_581_fu_15045_p4;
wire   [7:0] tmp_590_fu_15123_p4;
wire   [7:0] tmp_592_fu_15137_p4;
wire   [7:0] xor_ln1545_433_fu_15425_p2;
wire   [7:0] xor_ln1545_432_fu_15419_p2;
wire   [7:0] tmp_585_fu_15079_p4;
wire   [7:0] tmp_580_fu_15035_p4;
wire   [7:0] trunc_ln674_143_fu_15099_p1;
wire   [7:0] tmp_594_fu_15157_p4;
wire   [7:0] xor_ln1545_437_fu_15443_p2;
wire   [7:0] xor_ln1545_435_fu_15437_p2;
wire   [7:0] xor_ln1545_391_fu_15179_p2;
wire   [7:0] tmp_1_V_8_fu_15413_p2;
wire   [7:0] tmp_2_1_V_8_fu_15359_p2;
wire   [7:0] xor_ln1545_412_fu_15305_p2;
wire   [7:0] xor_ln1545_403_fu_15251_p2;
wire   [7:0] xor_ln1545_394_fu_15197_p2;
wire   [7:0] tmp_2_2_V_8_fu_15431_p2;
wire   [7:0] xor_ln1545_424_fu_15377_p2;
wire   [7:0] xor_ln1545_415_fu_15323_p2;
wire   [7:0] xor_ln1545_406_fu_15269_p2;
wire   [7:0] xor_ln1545_397_fu_15215_p2;
wire   [7:0] xor_ln1545_436_fu_15449_p2;
wire   [7:0] xor_ln1545_427_fu_15395_p2;
wire   [7:0] xor_ln1545_418_fu_15341_p2;
wire   [7:0] xor_ln1545_409_fu_15287_p2;
wire   [7:0] tmp_3_V_8_fu_15233_p2;
wire   [127:0] p_Result_33_fu_15535_p17;
wire   [127:0] state_V_32_fu_15571_p2;
wire   [7:0] trunc_ln708_10_fu_15576_p1;
wire   [7:0] tmp_598_fu_15585_p4;
wire   [7:0] tmp_602_fu_15600_p4;
wire   [7:0] tmp_606_fu_15615_p4;
wire   [7:0] tmp_610_fu_15630_p4;
wire   [7:0] tmp_614_fu_15645_p4;
wire   [7:0] tmp_618_fu_15660_p4;
wire   [7:0] tmp_622_fu_15675_p4;
wire   [7:0] tmp_626_fu_15690_p4;
wire   [7:0] tmp_630_fu_15705_p4;
wire   [7:0] tmp_634_fu_15720_p4;
wire   [7:0] tmp_638_fu_15735_p4;
wire   [7:0] tmp_642_fu_15750_p4;
wire   [7:0] tmp_646_fu_15765_p4;
wire   [7:0] tmp_650_fu_15780_p4;
wire   [7:0] tmp_654_fu_15795_p4;
wire   [7:0] tmp_599_fu_15848_p4;
wire   [7:0] tmp_597_fu_15834_p4;
wire   [7:0] tmp_604_fu_15892_p4;
wire   [7:0] trunc_ln674_148_fu_15912_p1;
wire   [7:0] xor_ln1545_440_fu_16360_p2;
wire   [7:0] xor_ln1545_438_fu_16354_p2;
wire   [7:0] tmp_601_fu_15868_p4;
wire   [7:0] trunc_ln674_145_fu_15810_p1;
wire   [7:0] tmp_603_fu_15882_p4;
wire   [7:0] tmp_608_fu_15926_p4;
wire   [7:0] xor_ln1545_443_fu_16378_p2;
wire   [7:0] xor_ln1545_441_fu_16372_p2;
wire   [7:0] trunc_ln674_146_fu_15844_p1;
wire   [7:0] tmp_596_fu_15824_p4;
wire   [7:0] tmp_605_fu_15902_p4;
wire   [7:0] tmp_607_fu_15916_p4;
wire   [7:0] xor_ln1545_446_fu_16396_p2;
wire   [7:0] xor_ln1545_444_fu_16390_p2;
wire   [7:0] tmp_600_fu_15858_p4;
wire   [7:0] tmp_595_fu_15814_p4;
wire   [7:0] trunc_ln674_147_fu_15878_p1;
wire   [7:0] tmp_609_fu_15936_p4;
wire   [7:0] xor_ln1545_448_fu_16414_p2;
wire   [7:0] xor_ln1545_447_fu_16408_p2;
wire   [7:0] tmp_615_fu_15984_p4;
wire   [7:0] tmp_613_fu_15970_p4;
wire   [7:0] tmp_620_fu_16028_p4;
wire   [7:0] trunc_ln674_152_fu_16048_p1;
wire   [7:0] xor_ln1545_452_fu_16432_p2;
wire   [7:0] xor_ln1545_450_fu_16426_p2;
wire   [7:0] tmp_617_fu_16004_p4;
wire   [7:0] trunc_ln674_149_fu_15946_p1;
wire   [7:0] tmp_619_fu_16018_p4;
wire   [7:0] tmp_624_fu_16062_p4;
wire   [7:0] xor_ln1545_455_fu_16450_p2;
wire   [7:0] xor_ln1545_453_fu_16444_p2;
wire   [7:0] trunc_ln674_150_fu_15980_p1;
wire   [7:0] tmp_612_fu_15960_p4;
wire   [7:0] tmp_621_fu_16038_p4;
wire   [7:0] tmp_623_fu_16052_p4;
wire   [7:0] xor_ln1545_458_fu_16468_p2;
wire   [7:0] xor_ln1545_456_fu_16462_p2;
wire   [7:0] tmp_616_fu_15994_p4;
wire   [7:0] tmp_611_fu_15950_p4;
wire   [7:0] trunc_ln674_151_fu_16014_p1;
wire   [7:0] tmp_625_fu_16072_p4;
wire   [7:0] xor_ln1545_461_fu_16486_p2;
wire   [7:0] xor_ln1545_459_fu_16480_p2;
wire   [7:0] tmp_631_fu_16120_p4;
wire   [7:0] tmp_629_fu_16106_p4;
wire   [7:0] tmp_636_fu_16164_p4;
wire   [7:0] trunc_ln674_156_fu_16184_p1;
wire   [7:0] xor_ln1545_464_fu_16504_p2;
wire   [7:0] xor_ln1545_462_fu_16498_p2;
wire   [7:0] tmp_633_fu_16140_p4;
wire   [7:0] trunc_ln674_153_fu_16082_p1;
wire   [7:0] tmp_635_fu_16154_p4;
wire   [7:0] tmp_640_fu_16198_p4;
wire   [7:0] xor_ln1545_467_fu_16522_p2;
wire   [7:0] xor_ln1545_465_fu_16516_p2;
wire   [7:0] trunc_ln674_154_fu_16116_p1;
wire   [7:0] tmp_628_fu_16096_p4;
wire   [7:0] tmp_637_fu_16174_p4;
wire   [7:0] tmp_639_fu_16188_p4;
wire   [7:0] xor_ln1545_469_fu_16540_p2;
wire   [7:0] xor_ln1545_468_fu_16534_p2;
wire   [7:0] tmp_632_fu_16130_p4;
wire   [7:0] tmp_627_fu_16086_p4;
wire   [7:0] trunc_ln674_155_fu_16150_p1;
wire   [7:0] tmp_641_fu_16208_p4;
wire   [7:0] xor_ln1545_473_fu_16558_p2;
wire   [7:0] xor_ln1545_471_fu_16552_p2;
wire   [7:0] tmp_647_fu_16256_p4;
wire   [7:0] tmp_645_fu_16242_p4;
wire   [7:0] tmp_652_fu_16300_p4;
wire   [7:0] trunc_ln674_160_fu_16320_p1;
wire   [7:0] xor_ln1545_476_fu_16576_p2;
wire   [7:0] xor_ln1545_474_fu_16570_p2;
wire   [7:0] tmp_649_fu_16276_p4;
wire   [7:0] trunc_ln674_157_fu_16218_p1;
wire   [7:0] tmp_651_fu_16290_p4;
wire   [7:0] tmp_656_fu_16334_p4;
wire   [7:0] xor_ln1545_478_fu_16594_p2;
wire   [7:0] xor_ln1545_477_fu_16588_p2;
wire   [7:0] trunc_ln674_158_fu_16252_p1;
wire   [7:0] tmp_644_fu_16232_p4;
wire   [7:0] tmp_653_fu_16310_p4;
wire   [7:0] tmp_655_fu_16324_p4;
wire   [7:0] xor_ln1545_481_fu_16612_p2;
wire   [7:0] xor_ln1545_480_fu_16606_p2;
wire   [7:0] tmp_648_fu_16266_p4;
wire   [7:0] tmp_643_fu_16222_p4;
wire   [7:0] trunc_ln674_159_fu_16286_p1;
wire   [7:0] tmp_657_fu_16344_p4;
wire   [7:0] xor_ln1545_485_fu_16630_p2;
wire   [7:0] xor_ln1545_483_fu_16624_p2;
wire   [7:0] xor_ln1545_439_fu_16366_p2;
wire   [7:0] tmp_1_V_9_fu_16600_p2;
wire   [7:0] tmp_2_1_V_9_fu_16546_p2;
wire   [7:0] xor_ln1545_460_fu_16492_p2;
wire   [7:0] xor_ln1545_451_fu_16438_p2;
wire   [7:0] xor_ln1545_442_fu_16384_p2;
wire   [7:0] tmp_2_2_V_9_fu_16618_p2;
wire   [7:0] xor_ln1545_472_fu_16564_p2;
wire   [7:0] xor_ln1545_463_fu_16510_p2;
wire   [7:0] xor_ln1545_454_fu_16456_p2;
wire   [7:0] xor_ln1545_445_fu_16402_p2;
wire   [7:0] xor_ln1545_484_fu_16636_p2;
wire   [7:0] xor_ln1545_475_fu_16582_p2;
wire   [7:0] xor_ln1545_466_fu_16528_p2;
wire   [7:0] xor_ln1545_457_fu_16474_p2;
wire   [7:0] tmp_3_V_9_fu_16420_p2;
wire   [127:0] p_Result_34_fu_16722_p17;
wire   [127:0] state_V_33_fu_16758_p2;
wire   [7:0] trunc_ln708_11_fu_16763_p1;
wire   [7:0] tmp_661_fu_16772_p4;
wire   [7:0] tmp_665_fu_16787_p4;
wire   [7:0] tmp_669_fu_16802_p4;
wire   [7:0] tmp_673_fu_16817_p4;
wire   [7:0] tmp_677_fu_16832_p4;
wire   [7:0] tmp_681_fu_16847_p4;
wire   [7:0] tmp_685_fu_16862_p4;
wire   [7:0] tmp_689_fu_16877_p4;
wire   [7:0] tmp_693_fu_16892_p4;
wire   [7:0] tmp_697_fu_16907_p4;
wire   [7:0] tmp_701_fu_16922_p4;
wire   [7:0] tmp_705_fu_16937_p4;
wire   [7:0] tmp_709_fu_16952_p4;
wire   [7:0] tmp_713_fu_16967_p4;
wire   [7:0] tmp_717_fu_16982_p4;
wire   [7:0] tmp_662_fu_17035_p4;
wire   [7:0] tmp_660_fu_17021_p4;
wire   [7:0] tmp_667_fu_17079_p4;
wire   [7:0] trunc_ln674_164_fu_17099_p1;
wire   [7:0] xor_ln1545_488_fu_17547_p2;
wire   [7:0] xor_ln1545_486_fu_17541_p2;
wire   [7:0] tmp_664_fu_17055_p4;
wire   [7:0] trunc_ln674_161_fu_16997_p1;
wire   [7:0] tmp_666_fu_17069_p4;
wire   [7:0] tmp_671_fu_17113_p4;
wire   [7:0] xor_ln1545_491_fu_17565_p2;
wire   [7:0] xor_ln1545_489_fu_17559_p2;
wire   [7:0] trunc_ln674_162_fu_17031_p1;
wire   [7:0] tmp_659_fu_17011_p4;
wire   [7:0] tmp_668_fu_17089_p4;
wire   [7:0] tmp_670_fu_17103_p4;
wire   [7:0] xor_ln1545_494_fu_17583_p2;
wire   [7:0] xor_ln1545_492_fu_17577_p2;
wire   [7:0] tmp_663_fu_17045_p4;
wire   [7:0] tmp_658_fu_17001_p4;
wire   [7:0] trunc_ln674_163_fu_17065_p1;
wire   [7:0] tmp_672_fu_17123_p4;
wire   [7:0] xor_ln1545_496_fu_17601_p2;
wire   [7:0] xor_ln1545_495_fu_17595_p2;
wire   [7:0] tmp_678_fu_17171_p4;
wire   [7:0] tmp_676_fu_17157_p4;
wire   [7:0] tmp_683_fu_17215_p4;
wire   [7:0] trunc_ln674_168_fu_17235_p1;
wire   [7:0] xor_ln1545_500_fu_17619_p2;
wire   [7:0] xor_ln1545_498_fu_17613_p2;
wire   [7:0] tmp_680_fu_17191_p4;
wire   [7:0] trunc_ln674_165_fu_17133_p1;
wire   [7:0] tmp_682_fu_17205_p4;
wire   [7:0] tmp_687_fu_17249_p4;
wire   [7:0] xor_ln1545_503_fu_17637_p2;
wire   [7:0] xor_ln1545_501_fu_17631_p2;
wire   [7:0] trunc_ln674_166_fu_17167_p1;
wire   [7:0] tmp_675_fu_17147_p4;
wire   [7:0] tmp_684_fu_17225_p4;
wire   [7:0] tmp_686_fu_17239_p4;
wire   [7:0] xor_ln1545_506_fu_17655_p2;
wire   [7:0] xor_ln1545_504_fu_17649_p2;
wire   [7:0] tmp_679_fu_17181_p4;
wire   [7:0] tmp_674_fu_17137_p4;
wire   [7:0] trunc_ln674_167_fu_17201_p1;
wire   [7:0] tmp_688_fu_17259_p4;
wire   [7:0] xor_ln1545_509_fu_17673_p2;
wire   [7:0] xor_ln1545_507_fu_17667_p2;
wire   [7:0] tmp_694_fu_17307_p4;
wire   [7:0] tmp_692_fu_17293_p4;
wire   [7:0] tmp_699_fu_17351_p4;
wire   [7:0] trunc_ln674_172_fu_17371_p1;
wire   [7:0] xor_ln1545_512_fu_17691_p2;
wire   [7:0] xor_ln1545_510_fu_17685_p2;
wire   [7:0] tmp_696_fu_17327_p4;
wire   [7:0] trunc_ln674_169_fu_17269_p1;
wire   [7:0] tmp_698_fu_17341_p4;
wire   [7:0] tmp_703_fu_17385_p4;
wire   [7:0] xor_ln1545_515_fu_17709_p2;
wire   [7:0] xor_ln1545_513_fu_17703_p2;
wire   [7:0] trunc_ln674_170_fu_17303_p1;
wire   [7:0] tmp_691_fu_17283_p4;
wire   [7:0] tmp_700_fu_17361_p4;
wire   [7:0] tmp_702_fu_17375_p4;
wire   [7:0] xor_ln1545_517_fu_17727_p2;
wire   [7:0] xor_ln1545_516_fu_17721_p2;
wire   [7:0] tmp_695_fu_17317_p4;
wire   [7:0] tmp_690_fu_17273_p4;
wire   [7:0] trunc_ln674_171_fu_17337_p1;
wire   [7:0] tmp_704_fu_17395_p4;
wire   [7:0] xor_ln1545_521_fu_17745_p2;
wire   [7:0] xor_ln1545_519_fu_17739_p2;
wire   [7:0] tmp_710_fu_17443_p4;
wire   [7:0] tmp_708_fu_17429_p4;
wire   [7:0] tmp_715_fu_17487_p4;
wire   [7:0] trunc_ln674_176_fu_17507_p1;
wire   [7:0] xor_ln1545_524_fu_17763_p2;
wire   [7:0] xor_ln1545_522_fu_17757_p2;
wire   [7:0] tmp_712_fu_17463_p4;
wire   [7:0] trunc_ln674_173_fu_17405_p1;
wire   [7:0] tmp_714_fu_17477_p4;
wire   [7:0] tmp_719_fu_17521_p4;
wire   [7:0] xor_ln1545_526_fu_17781_p2;
wire   [7:0] xor_ln1545_525_fu_17775_p2;
wire   [7:0] trunc_ln674_174_fu_17439_p1;
wire   [7:0] tmp_707_fu_17419_p4;
wire   [7:0] tmp_716_fu_17497_p4;
wire   [7:0] tmp_718_fu_17511_p4;
wire   [7:0] xor_ln1545_529_fu_17799_p2;
wire   [7:0] xor_ln1545_528_fu_17793_p2;
wire   [7:0] tmp_711_fu_17453_p4;
wire   [7:0] tmp_706_fu_17409_p4;
wire   [7:0] trunc_ln674_175_fu_17473_p1;
wire   [7:0] tmp_720_fu_17531_p4;
wire   [7:0] xor_ln1545_533_fu_17817_p2;
wire   [7:0] xor_ln1545_531_fu_17811_p2;
wire   [7:0] xor_ln1545_487_fu_17553_p2;
wire   [7:0] tmp_1_V_10_fu_17787_p2;
wire   [7:0] tmp_2_1_V_10_fu_17733_p2;
wire   [7:0] xor_ln1545_508_fu_17679_p2;
wire   [7:0] xor_ln1545_499_fu_17625_p2;
wire   [7:0] xor_ln1545_490_fu_17571_p2;
wire   [7:0] tmp_2_2_V_10_fu_17805_p2;
wire   [7:0] xor_ln1545_520_fu_17751_p2;
wire   [7:0] xor_ln1545_511_fu_17697_p2;
wire   [7:0] xor_ln1545_502_fu_17643_p2;
wire   [7:0] xor_ln1545_493_fu_17589_p2;
wire   [7:0] xor_ln1545_532_fu_17823_p2;
wire   [7:0] xor_ln1545_523_fu_17769_p2;
wire   [7:0] xor_ln1545_514_fu_17715_p2;
wire   [7:0] xor_ln1545_505_fu_17661_p2;
wire   [7:0] tmp_3_V_10_fu_17607_p2;
wire   [127:0] p_Result_35_fu_17909_p17;
reg   [0:0] ap_NS_fsm;
reg    ap_idle_pp0_0to22;
reg    ap_reset_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 1'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter5 = 1'b0;
#0 ap_enable_reg_pp0_iter6 = 1'b0;
#0 ap_enable_reg_pp0_iter7 = 1'b0;
#0 ap_enable_reg_pp0_iter8 = 1'b0;
#0 ap_enable_reg_pp0_iter9 = 1'b0;
#0 ap_enable_reg_pp0_iter10 = 1'b0;
#0 ap_enable_reg_pp0_iter11 = 1'b0;
#0 ap_enable_reg_pp0_iter12 = 1'b0;
#0 ap_enable_reg_pp0_iter13 = 1'b0;
#0 ap_enable_reg_pp0_iter14 = 1'b0;
#0 ap_enable_reg_pp0_iter15 = 1'b0;
#0 ap_enable_reg_pp0_iter16 = 1'b0;
#0 ap_enable_reg_pp0_iter17 = 1'b0;
#0 ap_enable_reg_pp0_iter18 = 1'b0;
#0 ap_enable_reg_pp0_iter19 = 1'b0;
#0 ap_enable_reg_pp0_iter20 = 1'b0;
#0 ap_enable_reg_pp0_iter21 = 1'b0;
#0 ap_enable_reg_pp0_iter22 = 1'b0;
#0 ap_enable_reg_pp0_iter23 = 1'b0;
end

testDec_process_r_decipher_0_iibox_ROM_NP_LUTRAM_1R #(
    .DataWidth( 8 ),
    .AddressRange( 256 ),
    .AddressWidth( 8 ))
decipher_0_iibox_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(decipher_0_iibox_address0),
    .ce0(decipher_0_iibox_ce0),
    .q0(decipher_0_iibox_q0),
    .address1(decipher_0_iibox_address1),
    .ce1(decipher_0_iibox_ce1),
    .q1(decipher_0_iibox_q1),
    .address2(decipher_0_iibox_address2),
    .ce2(decipher_0_iibox_ce2),
    .q2(decipher_0_iibox_q2),
    .address3(decipher_0_iibox_address3),
    .ce3(decipher_0_iibox_ce3),
    .q3(decipher_0_iibox_q3),
    .address4(decipher_0_iibox_address4),
    .ce4(decipher_0_iibox_ce4),
    .q4(decipher_0_iibox_q4),
    .address5(decipher_0_iibox_address5),
    .ce5(decipher_0_iibox_ce5),
    .q5(decipher_0_iibox_q5),
    .address6(decipher_0_iibox_address6),
    .ce6(decipher_0_iibox_ce6),
    .q6(decipher_0_iibox_q6),
    .address7(decipher_0_iibox_address7),
    .ce7(decipher_0_iibox_ce7),
    .q7(decipher_0_iibox_q7),
    .address8(decipher_0_iibox_address8),
    .ce8(decipher_0_iibox_ce8),
    .q8(decipher_0_iibox_q8),
    .address9(decipher_0_iibox_address9),
    .ce9(decipher_0_iibox_ce9),
    .q9(decipher_0_iibox_q9),
    .address10(decipher_0_iibox_address10),
    .ce10(decipher_0_iibox_ce10),
    .q10(decipher_0_iibox_q10),
    .address11(decipher_0_iibox_address11),
    .ce11(decipher_0_iibox_ce11),
    .q11(decipher_0_iibox_q11),
    .address12(decipher_0_iibox_address12),
    .ce12(decipher_0_iibox_ce12),
    .q12(decipher_0_iibox_q12),
    .address13(decipher_0_iibox_address13),
    .ce13(decipher_0_iibox_ce13),
    .q13(decipher_0_iibox_q13),
    .address14(decipher_0_iibox_address14),
    .ce14(decipher_0_iibox_ce14),
    .q14(decipher_0_iibox_q14),
    .address15(decipher_0_iibox_address15),
    .ce15(decipher_0_iibox_ce15),
    .q15(decipher_0_iibox_q15),
    .address16(decipher_0_iibox_address16),
    .ce16(decipher_0_iibox_ce16),
    .q16(decipher_0_iibox_q16),
    .address17(decipher_0_iibox_address17),
    .ce17(decipher_0_iibox_ce17),
    .q17(decipher_0_iibox_q17),
    .address18(decipher_0_iibox_address18),
    .ce18(decipher_0_iibox_ce18),
    .q18(decipher_0_iibox_q18),
    .address19(decipher_0_iibox_address19),
    .ce19(decipher_0_iibox_ce19),
    .q19(decipher_0_iibox_q19),
    .address20(decipher_0_iibox_address20),
    .ce20(decipher_0_iibox_ce20),
    .q20(decipher_0_iibox_q20),
    .address21(decipher_0_iibox_address21),
    .ce21(decipher_0_iibox_ce21),
    .q21(decipher_0_iibox_q21),
    .address22(decipher_0_iibox_address22),
    .ce22(decipher_0_iibox_ce22),
    .q22(decipher_0_iibox_q22),
    .address23(decipher_0_iibox_address23),
    .ce23(decipher_0_iibox_ce23),
    .q23(decipher_0_iibox_q23),
    .address24(decipher_0_iibox_address24),
    .ce24(decipher_0_iibox_ce24),
    .q24(decipher_0_iibox_q24),
    .address25(decipher_0_iibox_address25),
    .ce25(decipher_0_iibox_ce25),
    .q25(decipher_0_iibox_q25),
    .address26(decipher_0_iibox_address26),
    .ce26(decipher_0_iibox_ce26),
    .q26(decipher_0_iibox_q26),
    .address27(decipher_0_iibox_address27),
    .ce27(decipher_0_iibox_ce27),
    .q27(decipher_0_iibox_q27),
    .address28(decipher_0_iibox_address28),
    .ce28(decipher_0_iibox_ce28),
    .q28(decipher_0_iibox_q28),
    .address29(decipher_0_iibox_address29),
    .ce29(decipher_0_iibox_ce29),
    .q29(decipher_0_iibox_q29),
    .address30(decipher_0_iibox_address30),
    .ce30(decipher_0_iibox_ce30),
    .q30(decipher_0_iibox_q30),
    .address31(decipher_0_iibox_address31),
    .ce31(decipher_0_iibox_ce31),
    .q31(decipher_0_iibox_q31),
    .address32(decipher_0_iibox_address32),
    .ce32(decipher_0_iibox_ce32),
    .q32(decipher_0_iibox_q32),
    .address33(decipher_0_iibox_address33),
    .ce33(decipher_0_iibox_ce33),
    .q33(decipher_0_iibox_q33),
    .address34(decipher_0_iibox_address34),
    .ce34(decipher_0_iibox_ce34),
    .q34(decipher_0_iibox_q34),
    .address35(decipher_0_iibox_address35),
    .ce35(decipher_0_iibox_ce35),
    .q35(decipher_0_iibox_q35),
    .address36(decipher_0_iibox_address36),
    .ce36(decipher_0_iibox_ce36),
    .q36(decipher_0_iibox_q36),
    .address37(decipher_0_iibox_address37),
    .ce37(decipher_0_iibox_ce37),
    .q37(decipher_0_iibox_q37),
    .address38(decipher_0_iibox_address38),
    .ce38(decipher_0_iibox_ce38),
    .q38(decipher_0_iibox_q38),
    .address39(decipher_0_iibox_address39),
    .ce39(decipher_0_iibox_ce39),
    .q39(decipher_0_iibox_q39),
    .address40(decipher_0_iibox_address40),
    .ce40(decipher_0_iibox_ce40),
    .q40(decipher_0_iibox_q40),
    .address41(decipher_0_iibox_address41),
    .ce41(decipher_0_iibox_ce41),
    .q41(decipher_0_iibox_q41),
    .address42(decipher_0_iibox_address42),
    .ce42(decipher_0_iibox_ce42),
    .q42(decipher_0_iibox_q42),
    .address43(decipher_0_iibox_address43),
    .ce43(decipher_0_iibox_ce43),
    .q43(decipher_0_iibox_q43),
    .address44(decipher_0_iibox_address44),
    .ce44(decipher_0_iibox_ce44),
    .q44(decipher_0_iibox_q44),
    .address45(decipher_0_iibox_address45),
    .ce45(decipher_0_iibox_ce45),
    .q45(decipher_0_iibox_q45),
    .address46(decipher_0_iibox_address46),
    .ce46(decipher_0_iibox_ce46),
    .q46(decipher_0_iibox_q46),
    .address47(decipher_0_iibox_address47),
    .ce47(decipher_0_iibox_ce47),
    .q47(decipher_0_iibox_q47),
    .address48(decipher_0_iibox_address48),
    .ce48(decipher_0_iibox_ce48),
    .q48(decipher_0_iibox_q48),
    .address49(decipher_0_iibox_address49),
    .ce49(decipher_0_iibox_ce49),
    .q49(decipher_0_iibox_q49),
    .address50(decipher_0_iibox_address50),
    .ce50(decipher_0_iibox_ce50),
    .q50(decipher_0_iibox_q50),
    .address51(decipher_0_iibox_address51),
    .ce51(decipher_0_iibox_ce51),
    .q51(decipher_0_iibox_q51),
    .address52(decipher_0_iibox_address52),
    .ce52(decipher_0_iibox_ce52),
    .q52(decipher_0_iibox_q52),
    .address53(decipher_0_iibox_address53),
    .ce53(decipher_0_iibox_ce53),
    .q53(decipher_0_iibox_q53),
    .address54(decipher_0_iibox_address54),
    .ce54(decipher_0_iibox_ce54),
    .q54(decipher_0_iibox_q54),
    .address55(decipher_0_iibox_address55),
    .ce55(decipher_0_iibox_ce55),
    .q55(decipher_0_iibox_q55),
    .address56(decipher_0_iibox_address56),
    .ce56(decipher_0_iibox_ce56),
    .q56(decipher_0_iibox_q56),
    .address57(decipher_0_iibox_address57),
    .ce57(decipher_0_iibox_ce57),
    .q57(decipher_0_iibox_q57),
    .address58(decipher_0_iibox_address58),
    .ce58(decipher_0_iibox_ce58),
    .q58(decipher_0_iibox_q58),
    .address59(decipher_0_iibox_address59),
    .ce59(decipher_0_iibox_ce59),
    .q59(decipher_0_iibox_q59),
    .address60(decipher_0_iibox_address60),
    .ce60(decipher_0_iibox_ce60),
    .q60(decipher_0_iibox_q60),
    .address61(decipher_0_iibox_address61),
    .ce61(decipher_0_iibox_ce61),
    .q61(decipher_0_iibox_q61),
    .address62(decipher_0_iibox_address62),
    .ce62(decipher_0_iibox_ce62),
    .q62(decipher_0_iibox_q62),
    .address63(decipher_0_iibox_address63),
    .ce63(decipher_0_iibox_ce63),
    .q63(decipher_0_iibox_q63),
    .address64(decipher_0_iibox_address64),
    .ce64(decipher_0_iibox_ce64),
    .q64(decipher_0_iibox_q64),
    .address65(decipher_0_iibox_address65),
    .ce65(decipher_0_iibox_ce65),
    .q65(decipher_0_iibox_q65),
    .address66(decipher_0_iibox_address66),
    .ce66(decipher_0_iibox_ce66),
    .q66(decipher_0_iibox_q66),
    .address67(decipher_0_iibox_address67),
    .ce67(decipher_0_iibox_ce67),
    .q67(decipher_0_iibox_q67),
    .address68(decipher_0_iibox_address68),
    .ce68(decipher_0_iibox_ce68),
    .q68(decipher_0_iibox_q68),
    .address69(decipher_0_iibox_address69),
    .ce69(decipher_0_iibox_ce69),
    .q69(decipher_0_iibox_q69),
    .address70(decipher_0_iibox_address70),
    .ce70(decipher_0_iibox_ce70),
    .q70(decipher_0_iibox_q70),
    .address71(decipher_0_iibox_address71),
    .ce71(decipher_0_iibox_ce71),
    .q71(decipher_0_iibox_q71),
    .address72(decipher_0_iibox_address72),
    .ce72(decipher_0_iibox_ce72),
    .q72(decipher_0_iibox_q72),
    .address73(decipher_0_iibox_address73),
    .ce73(decipher_0_iibox_ce73),
    .q73(decipher_0_iibox_q73),
    .address74(decipher_0_iibox_address74),
    .ce74(decipher_0_iibox_ce74),
    .q74(decipher_0_iibox_q74),
    .address75(decipher_0_iibox_address75),
    .ce75(decipher_0_iibox_ce75),
    .q75(decipher_0_iibox_q75),
    .address76(decipher_0_iibox_address76),
    .ce76(decipher_0_iibox_ce76),
    .q76(decipher_0_iibox_q76),
    .address77(decipher_0_iibox_address77),
    .ce77(decipher_0_iibox_ce77),
    .q77(decipher_0_iibox_q77),
    .address78(decipher_0_iibox_address78),
    .ce78(decipher_0_iibox_ce78),
    .q78(decipher_0_iibox_q78),
    .address79(decipher_0_iibox_address79),
    .ce79(decipher_0_iibox_ce79),
    .q79(decipher_0_iibox_q79),
    .address80(decipher_0_iibox_address80),
    .ce80(decipher_0_iibox_ce80),
    .q80(decipher_0_iibox_q80),
    .address81(decipher_0_iibox_address81),
    .ce81(decipher_0_iibox_ce81),
    .q81(decipher_0_iibox_q81),
    .address82(decipher_0_iibox_address82),
    .ce82(decipher_0_iibox_ce82),
    .q82(decipher_0_iibox_q82),
    .address83(decipher_0_iibox_address83),
    .ce83(decipher_0_iibox_ce83),
    .q83(decipher_0_iibox_q83),
    .address84(decipher_0_iibox_address84),
    .ce84(decipher_0_iibox_ce84),
    .q84(decipher_0_iibox_q84),
    .address85(decipher_0_iibox_address85),
    .ce85(decipher_0_iibox_ce85),
    .q85(decipher_0_iibox_q85),
    .address86(decipher_0_iibox_address86),
    .ce86(decipher_0_iibox_ce86),
    .q86(decipher_0_iibox_q86),
    .address87(decipher_0_iibox_address87),
    .ce87(decipher_0_iibox_ce87),
    .q87(decipher_0_iibox_q87),
    .address88(decipher_0_iibox_address88),
    .ce88(decipher_0_iibox_ce88),
    .q88(decipher_0_iibox_q88),
    .address89(decipher_0_iibox_address89),
    .ce89(decipher_0_iibox_ce89),
    .q89(decipher_0_iibox_q89),
    .address90(decipher_0_iibox_address90),
    .ce90(decipher_0_iibox_ce90),
    .q90(decipher_0_iibox_q90),
    .address91(decipher_0_iibox_address91),
    .ce91(decipher_0_iibox_ce91),
    .q91(decipher_0_iibox_q91),
    .address92(decipher_0_iibox_address92),
    .ce92(decipher_0_iibox_ce92),
    .q92(decipher_0_iibox_q92),
    .address93(decipher_0_iibox_address93),
    .ce93(decipher_0_iibox_ce93),
    .q93(decipher_0_iibox_q93),
    .address94(decipher_0_iibox_address94),
    .ce94(decipher_0_iibox_ce94),
    .q94(decipher_0_iibox_q94),
    .address95(decipher_0_iibox_address95),
    .ce95(decipher_0_iibox_ce95),
    .q95(decipher_0_iibox_q95),
    .address96(decipher_0_iibox_address96),
    .ce96(decipher_0_iibox_ce96),
    .q96(decipher_0_iibox_q96),
    .address97(decipher_0_iibox_address97),
    .ce97(decipher_0_iibox_ce97),
    .q97(decipher_0_iibox_q97),
    .address98(decipher_0_iibox_address98),
    .ce98(decipher_0_iibox_ce98),
    .q98(decipher_0_iibox_q98),
    .address99(decipher_0_iibox_address99),
    .ce99(decipher_0_iibox_ce99),
    .q99(decipher_0_iibox_q99),
    .address100(decipher_0_iibox_address100),
    .ce100(decipher_0_iibox_ce100),
    .q100(decipher_0_iibox_q100),
    .address101(decipher_0_iibox_address101),
    .ce101(decipher_0_iibox_ce101),
    .q101(decipher_0_iibox_q101),
    .address102(decipher_0_iibox_address102),
    .ce102(decipher_0_iibox_ce102),
    .q102(decipher_0_iibox_q102),
    .address103(decipher_0_iibox_address103),
    .ce103(decipher_0_iibox_ce103),
    .q103(decipher_0_iibox_q103),
    .address104(decipher_0_iibox_address104),
    .ce104(decipher_0_iibox_ce104),
    .q104(decipher_0_iibox_q104),
    .address105(decipher_0_iibox_address105),
    .ce105(decipher_0_iibox_ce105),
    .q105(decipher_0_iibox_q105),
    .address106(decipher_0_iibox_address106),
    .ce106(decipher_0_iibox_ce106),
    .q106(decipher_0_iibox_q106),
    .address107(decipher_0_iibox_address107),
    .ce107(decipher_0_iibox_ce107),
    .q107(decipher_0_iibox_q107),
    .address108(decipher_0_iibox_address108),
    .ce108(decipher_0_iibox_ce108),
    .q108(decipher_0_iibox_q108),
    .address109(decipher_0_iibox_address109),
    .ce109(decipher_0_iibox_ce109),
    .q109(decipher_0_iibox_q109),
    .address110(decipher_0_iibox_address110),
    .ce110(decipher_0_iibox_ce110),
    .q110(decipher_0_iibox_q110),
    .address111(decipher_0_iibox_address111),
    .ce111(decipher_0_iibox_ce111),
    .q111(decipher_0_iibox_q111),
    .address112(decipher_0_iibox_address112),
    .ce112(decipher_0_iibox_ce112),
    .q112(decipher_0_iibox_q112),
    .address113(decipher_0_iibox_address113),
    .ce113(decipher_0_iibox_ce113),
    .q113(decipher_0_iibox_q113),
    .address114(decipher_0_iibox_address114),
    .ce114(decipher_0_iibox_ce114),
    .q114(decipher_0_iibox_q114),
    .address115(decipher_0_iibox_address115),
    .ce115(decipher_0_iibox_ce115),
    .q115(decipher_0_iibox_q115),
    .address116(decipher_0_iibox_address116),
    .ce116(decipher_0_iibox_ce116),
    .q116(decipher_0_iibox_q116),
    .address117(decipher_0_iibox_address117),
    .ce117(decipher_0_iibox_ce117),
    .q117(decipher_0_iibox_q117),
    .address118(decipher_0_iibox_address118),
    .ce118(decipher_0_iibox_ce118),
    .q118(decipher_0_iibox_q118),
    .address119(decipher_0_iibox_address119),
    .ce119(decipher_0_iibox_ce119),
    .q119(decipher_0_iibox_q119),
    .address120(decipher_0_iibox_address120),
    .ce120(decipher_0_iibox_ce120),
    .q120(decipher_0_iibox_q120),
    .address121(decipher_0_iibox_address121),
    .ce121(decipher_0_iibox_ce121),
    .q121(decipher_0_iibox_q121),
    .address122(decipher_0_iibox_address122),
    .ce122(decipher_0_iibox_ce122),
    .q122(decipher_0_iibox_q122),
    .address123(decipher_0_iibox_address123),
    .ce123(decipher_0_iibox_ce123),
    .q123(decipher_0_iibox_q123),
    .address124(decipher_0_iibox_address124),
    .ce124(decipher_0_iibox_ce124),
    .q124(decipher_0_iibox_q124),
    .address125(decipher_0_iibox_address125),
    .ce125(decipher_0_iibox_ce125),
    .q125(decipher_0_iibox_q125),
    .address126(decipher_0_iibox_address126),
    .ce126(decipher_0_iibox_ce126),
    .q126(decipher_0_iibox_q126),
    .address127(decipher_0_iibox_address127),
    .ce127(decipher_0_iibox_ce127),
    .q127(decipher_0_iibox_q127),
    .address128(decipher_0_iibox_address128),
    .ce128(decipher_0_iibox_ce128),
    .q128(decipher_0_iibox_q128),
    .address129(decipher_0_iibox_address129),
    .ce129(decipher_0_iibox_ce129),
    .q129(decipher_0_iibox_q129),
    .address130(decipher_0_iibox_address130),
    .ce130(decipher_0_iibox_ce130),
    .q130(decipher_0_iibox_q130),
    .address131(decipher_0_iibox_address131),
    .ce131(decipher_0_iibox_ce131),
    .q131(decipher_0_iibox_q131),
    .address132(decipher_0_iibox_address132),
    .ce132(decipher_0_iibox_ce132),
    .q132(decipher_0_iibox_q132),
    .address133(decipher_0_iibox_address133),
    .ce133(decipher_0_iibox_ce133),
    .q133(decipher_0_iibox_q133),
    .address134(decipher_0_iibox_address134),
    .ce134(decipher_0_iibox_ce134),
    .q134(decipher_0_iibox_q134),
    .address135(decipher_0_iibox_address135),
    .ce135(decipher_0_iibox_ce135),
    .q135(decipher_0_iibox_q135),
    .address136(decipher_0_iibox_address136),
    .ce136(decipher_0_iibox_ce136),
    .q136(decipher_0_iibox_q136),
    .address137(decipher_0_iibox_address137),
    .ce137(decipher_0_iibox_ce137),
    .q137(decipher_0_iibox_q137),
    .address138(decipher_0_iibox_address138),
    .ce138(decipher_0_iibox_ce138),
    .q138(decipher_0_iibox_q138),
    .address139(decipher_0_iibox_address139),
    .ce139(decipher_0_iibox_ce139),
    .q139(decipher_0_iibox_q139),
    .address140(decipher_0_iibox_address140),
    .ce140(decipher_0_iibox_ce140),
    .q140(decipher_0_iibox_q140),
    .address141(decipher_0_iibox_address141),
    .ce141(decipher_0_iibox_ce141),
    .q141(decipher_0_iibox_q141),
    .address142(decipher_0_iibox_address142),
    .ce142(decipher_0_iibox_ce142),
    .q142(decipher_0_iibox_q142),
    .address143(decipher_0_iibox_address143),
    .ce143(decipher_0_iibox_ce143),
    .q143(decipher_0_iibox_q143),
    .address144(decipher_0_iibox_address144),
    .ce144(decipher_0_iibox_ce144),
    .q144(decipher_0_iibox_q144),
    .address145(decipher_0_iibox_address145),
    .ce145(decipher_0_iibox_ce145),
    .q145(decipher_0_iibox_q145),
    .address146(decipher_0_iibox_address146),
    .ce146(decipher_0_iibox_ce146),
    .q146(decipher_0_iibox_q146),
    .address147(decipher_0_iibox_address147),
    .ce147(decipher_0_iibox_ce147),
    .q147(decipher_0_iibox_q147),
    .address148(decipher_0_iibox_address148),
    .ce148(decipher_0_iibox_ce148),
    .q148(decipher_0_iibox_q148),
    .address149(decipher_0_iibox_address149),
    .ce149(decipher_0_iibox_ce149),
    .q149(decipher_0_iibox_q149),
    .address150(decipher_0_iibox_address150),
    .ce150(decipher_0_iibox_ce150),
    .q150(decipher_0_iibox_q150),
    .address151(decipher_0_iibox_address151),
    .ce151(decipher_0_iibox_ce151),
    .q151(decipher_0_iibox_q151),
    .address152(decipher_0_iibox_address152),
    .ce152(decipher_0_iibox_ce152),
    .q152(decipher_0_iibox_q152),
    .address153(decipher_0_iibox_address153),
    .ce153(decipher_0_iibox_ce153),
    .q153(decipher_0_iibox_q153),
    .address154(decipher_0_iibox_address154),
    .ce154(decipher_0_iibox_ce154),
    .q154(decipher_0_iibox_q154),
    .address155(decipher_0_iibox_address155),
    .ce155(decipher_0_iibox_ce155),
    .q155(decipher_0_iibox_q155),
    .address156(decipher_0_iibox_address156),
    .ce156(decipher_0_iibox_ce156),
    .q156(decipher_0_iibox_q156),
    .address157(decipher_0_iibox_address157),
    .ce157(decipher_0_iibox_ce157),
    .q157(decipher_0_iibox_q157),
    .address158(decipher_0_iibox_address158),
    .ce158(decipher_0_iibox_ce158),
    .q158(decipher_0_iibox_q158),
    .address159(decipher_0_iibox_address159),
    .ce159(decipher_0_iibox_ce159),
    .q159(decipher_0_iibox_q159),
    .address160(decipher_0_iibox_address160),
    .ce160(decipher_0_iibox_ce160),
    .q160(decipher_0_iibox_q160),
    .address161(decipher_0_iibox_address161),
    .ce161(decipher_0_iibox_ce161),
    .q161(decipher_0_iibox_q161),
    .address162(decipher_0_iibox_address162),
    .ce162(decipher_0_iibox_ce162),
    .q162(decipher_0_iibox_q162),
    .address163(decipher_0_iibox_address163),
    .ce163(decipher_0_iibox_ce163),
    .q163(decipher_0_iibox_q163),
    .address164(decipher_0_iibox_address164),
    .ce164(decipher_0_iibox_ce164),
    .q164(decipher_0_iibox_q164),
    .address165(decipher_0_iibox_address165),
    .ce165(decipher_0_iibox_ce165),
    .q165(decipher_0_iibox_q165),
    .address166(decipher_0_iibox_address166),
    .ce166(decipher_0_iibox_ce166),
    .q166(decipher_0_iibox_q166),
    .address167(decipher_0_iibox_address167),
    .ce167(decipher_0_iibox_ce167),
    .q167(decipher_0_iibox_q167),
    .address168(decipher_0_iibox_address168),
    .ce168(decipher_0_iibox_ce168),
    .q168(decipher_0_iibox_q168),
    .address169(decipher_0_iibox_address169),
    .ce169(decipher_0_iibox_ce169),
    .q169(decipher_0_iibox_q169),
    .address170(decipher_0_iibox_address170),
    .ce170(decipher_0_iibox_ce170),
    .q170(decipher_0_iibox_q170),
    .address171(decipher_0_iibox_address171),
    .ce171(decipher_0_iibox_ce171),
    .q171(decipher_0_iibox_q171),
    .address172(decipher_0_iibox_address172),
    .ce172(decipher_0_iibox_ce172),
    .q172(decipher_0_iibox_q172),
    .address173(decipher_0_iibox_address173),
    .ce173(decipher_0_iibox_ce173),
    .q173(decipher_0_iibox_q173),
    .address174(decipher_0_iibox_address174),
    .ce174(decipher_0_iibox_ce174),
    .q174(decipher_0_iibox_q174),
    .address175(decipher_0_iibox_address175),
    .ce175(decipher_0_iibox_ce175),
    .q175(decipher_0_iibox_q175),
    .address176(decipher_0_iibox_address176),
    .ce176(decipher_0_iibox_ce176),
    .q176(decipher_0_iibox_q176),
    .address177(decipher_0_iibox_address177),
    .ce177(decipher_0_iibox_ce177),
    .q177(decipher_0_iibox_q177),
    .address178(decipher_0_iibox_address178),
    .ce178(decipher_0_iibox_ce178),
    .q178(decipher_0_iibox_q178),
    .address179(decipher_0_iibox_address179),
    .ce179(decipher_0_iibox_ce179),
    .q179(decipher_0_iibox_q179),
    .address180(decipher_0_iibox_address180),
    .ce180(decipher_0_iibox_ce180),
    .q180(decipher_0_iibox_q180),
    .address181(decipher_0_iibox_address181),
    .ce181(decipher_0_iibox_ce181),
    .q181(decipher_0_iibox_q181),
    .address182(decipher_0_iibox_address182),
    .ce182(decipher_0_iibox_ce182),
    .q182(decipher_0_iibox_q182),
    .address183(decipher_0_iibox_address183),
    .ce183(decipher_0_iibox_ce183),
    .q183(decipher_0_iibox_q183),
    .address184(decipher_0_iibox_address184),
    .ce184(decipher_0_iibox_ce184),
    .q184(decipher_0_iibox_q184),
    .address185(decipher_0_iibox_address185),
    .ce185(decipher_0_iibox_ce185),
    .q185(decipher_0_iibox_q185),
    .address186(decipher_0_iibox_address186),
    .ce186(decipher_0_iibox_ce186),
    .q186(decipher_0_iibox_q186),
    .address187(decipher_0_iibox_address187),
    .ce187(decipher_0_iibox_ce187),
    .q187(decipher_0_iibox_q187),
    .address188(decipher_0_iibox_address188),
    .ce188(decipher_0_iibox_ce188),
    .q188(decipher_0_iibox_q188),
    .address189(decipher_0_iibox_address189),
    .ce189(decipher_0_iibox_ce189),
    .q189(decipher_0_iibox_q189),
    .address190(decipher_0_iibox_address190),
    .ce190(decipher_0_iibox_ce190),
    .q190(decipher_0_iibox_q190),
    .address191(decipher_0_iibox_address191),
    .ce191(decipher_0_iibox_ce191),
    .q191(decipher_0_iibox_q191)
);

testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R #(
    .DataWidth( 32 ),
    .AddressRange( 256 ),
    .AddressWidth( 8 ))
decipher_0_i32box_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(decipher_0_i32box_address0),
    .ce0(decipher_0_i32box_ce0),
    .q0(decipher_0_i32box_q0),
    .address1(decipher_0_i32box_address1),
    .ce1(decipher_0_i32box_ce1),
    .q1(decipher_0_i32box_q1),
    .address2(decipher_0_i32box_address2),
    .ce2(decipher_0_i32box_ce2),
    .q2(decipher_0_i32box_q2),
    .address3(decipher_0_i32box_address3),
    .ce3(decipher_0_i32box_ce3),
    .q3(decipher_0_i32box_q3),
    .address4(decipher_0_i32box_address4),
    .ce4(decipher_0_i32box_ce4),
    .q4(decipher_0_i32box_q4),
    .address5(decipher_0_i32box_address5),
    .ce5(decipher_0_i32box_ce5),
    .q5(decipher_0_i32box_q5),
    .address6(decipher_0_i32box_address6),
    .ce6(decipher_0_i32box_ce6),
    .q6(decipher_0_i32box_q6),
    .address7(decipher_0_i32box_address7),
    .ce7(decipher_0_i32box_ce7),
    .q7(decipher_0_i32box_q7),
    .address8(decipher_0_i32box_address8),
    .ce8(decipher_0_i32box_ce8),
    .q8(decipher_0_i32box_q8),
    .address9(decipher_0_i32box_address9),
    .ce9(decipher_0_i32box_ce9),
    .q9(decipher_0_i32box_q9),
    .address10(decipher_0_i32box_address10),
    .ce10(decipher_0_i32box_ce10),
    .q10(decipher_0_i32box_q10),
    .address11(decipher_0_i32box_address11),
    .ce11(decipher_0_i32box_ce11),
    .q11(decipher_0_i32box_q11),
    .address12(decipher_0_i32box_address12),
    .ce12(decipher_0_i32box_ce12),
    .q12(decipher_0_i32box_q12),
    .address13(decipher_0_i32box_address13),
    .ce13(decipher_0_i32box_ce13),
    .q13(decipher_0_i32box_q13),
    .address14(decipher_0_i32box_address14),
    .ce14(decipher_0_i32box_ce14),
    .q14(decipher_0_i32box_q14),
    .address15(decipher_0_i32box_address15),
    .ce15(decipher_0_i32box_ce15),
    .q15(decipher_0_i32box_q15),
    .address16(decipher_0_i32box_address16),
    .ce16(decipher_0_i32box_ce16),
    .q16(decipher_0_i32box_q16),
    .address17(decipher_0_i32box_address17),
    .ce17(decipher_0_i32box_ce17),
    .q17(decipher_0_i32box_q17),
    .address18(decipher_0_i32box_address18),
    .ce18(decipher_0_i32box_ce18),
    .q18(decipher_0_i32box_q18),
    .address19(decipher_0_i32box_address19),
    .ce19(decipher_0_i32box_ce19),
    .q19(decipher_0_i32box_q19),
    .address20(decipher_0_i32box_address20),
    .ce20(decipher_0_i32box_ce20),
    .q20(decipher_0_i32box_q20),
    .address21(decipher_0_i32box_address21),
    .ce21(decipher_0_i32box_ce21),
    .q21(decipher_0_i32box_q21),
    .address22(decipher_0_i32box_address22),
    .ce22(decipher_0_i32box_ce22),
    .q22(decipher_0_i32box_q22),
    .address23(decipher_0_i32box_address23),
    .ce23(decipher_0_i32box_ce23),
    .q23(decipher_0_i32box_q23),
    .address24(decipher_0_i32box_address24),
    .ce24(decipher_0_i32box_ce24),
    .q24(decipher_0_i32box_q24),
    .address25(decipher_0_i32box_address25),
    .ce25(decipher_0_i32box_ce25),
    .q25(decipher_0_i32box_q25),
    .address26(decipher_0_i32box_address26),
    .ce26(decipher_0_i32box_ce26),
    .q26(decipher_0_i32box_q26),
    .address27(decipher_0_i32box_address27),
    .ce27(decipher_0_i32box_ce27),
    .q27(decipher_0_i32box_q27),
    .address28(decipher_0_i32box_address28),
    .ce28(decipher_0_i32box_ce28),
    .q28(decipher_0_i32box_q28),
    .address29(decipher_0_i32box_address29),
    .ce29(decipher_0_i32box_ce29),
    .q29(decipher_0_i32box_q29),
    .address30(decipher_0_i32box_address30),
    .ce30(decipher_0_i32box_ce30),
    .q30(decipher_0_i32box_q30),
    .address31(decipher_0_i32box_address31),
    .ce31(decipher_0_i32box_ce31),
    .q31(decipher_0_i32box_q31),
    .address32(decipher_0_i32box_address32),
    .ce32(decipher_0_i32box_ce32),
    .q32(decipher_0_i32box_q32),
    .address33(decipher_0_i32box_address33),
    .ce33(decipher_0_i32box_ce33),
    .q33(decipher_0_i32box_q33),
    .address34(decipher_0_i32box_address34),
    .ce34(decipher_0_i32box_ce34),
    .q34(decipher_0_i32box_q34),
    .address35(decipher_0_i32box_address35),
    .ce35(decipher_0_i32box_ce35),
    .q35(decipher_0_i32box_q35),
    .address36(decipher_0_i32box_address36),
    .ce36(decipher_0_i32box_ce36),
    .q36(decipher_0_i32box_q36),
    .address37(decipher_0_i32box_address37),
    .ce37(decipher_0_i32box_ce37),
    .q37(decipher_0_i32box_q37),
    .address38(decipher_0_i32box_address38),
    .ce38(decipher_0_i32box_ce38),
    .q38(decipher_0_i32box_q38),
    .address39(decipher_0_i32box_address39),
    .ce39(decipher_0_i32box_ce39),
    .q39(decipher_0_i32box_q39),
    .address40(decipher_0_i32box_address40),
    .ce40(decipher_0_i32box_ce40),
    .q40(decipher_0_i32box_q40),
    .address41(decipher_0_i32box_address41),
    .ce41(decipher_0_i32box_ce41),
    .q41(decipher_0_i32box_q41),
    .address42(decipher_0_i32box_address42),
    .ce42(decipher_0_i32box_ce42),
    .q42(decipher_0_i32box_q42),
    .address43(decipher_0_i32box_address43),
    .ce43(decipher_0_i32box_ce43),
    .q43(decipher_0_i32box_q43),
    .address44(decipher_0_i32box_address44),
    .ce44(decipher_0_i32box_ce44),
    .q44(decipher_0_i32box_q44),
    .address45(decipher_0_i32box_address45),
    .ce45(decipher_0_i32box_ce45),
    .q45(decipher_0_i32box_q45),
    .address46(decipher_0_i32box_address46),
    .ce46(decipher_0_i32box_ce46),
    .q46(decipher_0_i32box_q46),
    .address47(decipher_0_i32box_address47),
    .ce47(decipher_0_i32box_ce47),
    .q47(decipher_0_i32box_q47),
    .address48(decipher_0_i32box_address48),
    .ce48(decipher_0_i32box_ce48),
    .q48(decipher_0_i32box_q48),
    .address49(decipher_0_i32box_address49),
    .ce49(decipher_0_i32box_ce49),
    .q49(decipher_0_i32box_q49),
    .address50(decipher_0_i32box_address50),
    .ce50(decipher_0_i32box_ce50),
    .q50(decipher_0_i32box_q50),
    .address51(decipher_0_i32box_address51),
    .ce51(decipher_0_i32box_ce51),
    .q51(decipher_0_i32box_q51),
    .address52(decipher_0_i32box_address52),
    .ce52(decipher_0_i32box_ce52),
    .q52(decipher_0_i32box_q52),
    .address53(decipher_0_i32box_address53),
    .ce53(decipher_0_i32box_ce53),
    .q53(decipher_0_i32box_q53),
    .address54(decipher_0_i32box_address54),
    .ce54(decipher_0_i32box_ce54),
    .q54(decipher_0_i32box_q54),
    .address55(decipher_0_i32box_address55),
    .ce55(decipher_0_i32box_ce55),
    .q55(decipher_0_i32box_q55),
    .address56(decipher_0_i32box_address56),
    .ce56(decipher_0_i32box_ce56),
    .q56(decipher_0_i32box_q56),
    .address57(decipher_0_i32box_address57),
    .ce57(decipher_0_i32box_ce57),
    .q57(decipher_0_i32box_q57),
    .address58(decipher_0_i32box_address58),
    .ce58(decipher_0_i32box_ce58),
    .q58(decipher_0_i32box_q58),
    .address59(decipher_0_i32box_address59),
    .ce59(decipher_0_i32box_ce59),
    .q59(decipher_0_i32box_q59),
    .address60(decipher_0_i32box_address60),
    .ce60(decipher_0_i32box_ce60),
    .q60(decipher_0_i32box_q60),
    .address61(decipher_0_i32box_address61),
    .ce61(decipher_0_i32box_ce61),
    .q61(decipher_0_i32box_q61),
    .address62(decipher_0_i32box_address62),
    .ce62(decipher_0_i32box_ce62),
    .q62(decipher_0_i32box_q62),
    .address63(decipher_0_i32box_address63),
    .ce63(decipher_0_i32box_ce63),
    .q63(decipher_0_i32box_q63),
    .address64(decipher_0_i32box_address64),
    .ce64(decipher_0_i32box_ce64),
    .q64(decipher_0_i32box_q64),
    .address65(decipher_0_i32box_address65),
    .ce65(decipher_0_i32box_ce65),
    .q65(decipher_0_i32box_q65),
    .address66(decipher_0_i32box_address66),
    .ce66(decipher_0_i32box_ce66),
    .q66(decipher_0_i32box_q66),
    .address67(decipher_0_i32box_address67),
    .ce67(decipher_0_i32box_ce67),
    .q67(decipher_0_i32box_q67),
    .address68(decipher_0_i32box_address68),
    .ce68(decipher_0_i32box_ce68),
    .q68(decipher_0_i32box_q68),
    .address69(decipher_0_i32box_address69),
    .ce69(decipher_0_i32box_ce69),
    .q69(decipher_0_i32box_q69),
    .address70(decipher_0_i32box_address70),
    .ce70(decipher_0_i32box_ce70),
    .q70(decipher_0_i32box_q70),
    .address71(decipher_0_i32box_address71),
    .ce71(decipher_0_i32box_ce71),
    .q71(decipher_0_i32box_q71),
    .address72(decipher_0_i32box_address72),
    .ce72(decipher_0_i32box_ce72),
    .q72(decipher_0_i32box_q72),
    .address73(decipher_0_i32box_address73),
    .ce73(decipher_0_i32box_ce73),
    .q73(decipher_0_i32box_q73),
    .address74(decipher_0_i32box_address74),
    .ce74(decipher_0_i32box_ce74),
    .q74(decipher_0_i32box_q74),
    .address75(decipher_0_i32box_address75),
    .ce75(decipher_0_i32box_ce75),
    .q75(decipher_0_i32box_q75),
    .address76(decipher_0_i32box_address76),
    .ce76(decipher_0_i32box_ce76),
    .q76(decipher_0_i32box_q76),
    .address77(decipher_0_i32box_address77),
    .ce77(decipher_0_i32box_ce77),
    .q77(decipher_0_i32box_q77),
    .address78(decipher_0_i32box_address78),
    .ce78(decipher_0_i32box_ce78),
    .q78(decipher_0_i32box_q78),
    .address79(decipher_0_i32box_address79),
    .ce79(decipher_0_i32box_ce79),
    .q79(decipher_0_i32box_q79),
    .address80(decipher_0_i32box_address80),
    .ce80(decipher_0_i32box_ce80),
    .q80(decipher_0_i32box_q80),
    .address81(decipher_0_i32box_address81),
    .ce81(decipher_0_i32box_ce81),
    .q81(decipher_0_i32box_q81),
    .address82(decipher_0_i32box_address82),
    .ce82(decipher_0_i32box_ce82),
    .q82(decipher_0_i32box_q82),
    .address83(decipher_0_i32box_address83),
    .ce83(decipher_0_i32box_ce83),
    .q83(decipher_0_i32box_q83),
    .address84(decipher_0_i32box_address84),
    .ce84(decipher_0_i32box_ce84),
    .q84(decipher_0_i32box_q84),
    .address85(decipher_0_i32box_address85),
    .ce85(decipher_0_i32box_ce85),
    .q85(decipher_0_i32box_q85),
    .address86(decipher_0_i32box_address86),
    .ce86(decipher_0_i32box_ce86),
    .q86(decipher_0_i32box_q86),
    .address87(decipher_0_i32box_address87),
    .ce87(decipher_0_i32box_ce87),
    .q87(decipher_0_i32box_q87),
    .address88(decipher_0_i32box_address88),
    .ce88(decipher_0_i32box_ce88),
    .q88(decipher_0_i32box_q88),
    .address89(decipher_0_i32box_address89),
    .ce89(decipher_0_i32box_ce89),
    .q89(decipher_0_i32box_q89),
    .address90(decipher_0_i32box_address90),
    .ce90(decipher_0_i32box_ce90),
    .q90(decipher_0_i32box_q90),
    .address91(decipher_0_i32box_address91),
    .ce91(decipher_0_i32box_ce91),
    .q91(decipher_0_i32box_q91),
    .address92(decipher_0_i32box_address92),
    .ce92(decipher_0_i32box_ce92),
    .q92(decipher_0_i32box_q92),
    .address93(decipher_0_i32box_address93),
    .ce93(decipher_0_i32box_ce93),
    .q93(decipher_0_i32box_q93),
    .address94(decipher_0_i32box_address94),
    .ce94(decipher_0_i32box_ce94),
    .q94(decipher_0_i32box_q94),
    .address95(decipher_0_i32box_address95),
    .ce95(decipher_0_i32box_ce95),
    .q95(decipher_0_i32box_q95),
    .address96(decipher_0_i32box_address96),
    .ce96(decipher_0_i32box_ce96),
    .q96(decipher_0_i32box_q96),
    .address97(decipher_0_i32box_address97),
    .ce97(decipher_0_i32box_ce97),
    .q97(decipher_0_i32box_q97),
    .address98(decipher_0_i32box_address98),
    .ce98(decipher_0_i32box_ce98),
    .q98(decipher_0_i32box_q98),
    .address99(decipher_0_i32box_address99),
    .ce99(decipher_0_i32box_ce99),
    .q99(decipher_0_i32box_q99),
    .address100(decipher_0_i32box_address100),
    .ce100(decipher_0_i32box_ce100),
    .q100(decipher_0_i32box_q100),
    .address101(decipher_0_i32box_address101),
    .ce101(decipher_0_i32box_ce101),
    .q101(decipher_0_i32box_q101),
    .address102(decipher_0_i32box_address102),
    .ce102(decipher_0_i32box_ce102),
    .q102(decipher_0_i32box_q102),
    .address103(decipher_0_i32box_address103),
    .ce103(decipher_0_i32box_ce103),
    .q103(decipher_0_i32box_q103),
    .address104(decipher_0_i32box_address104),
    .ce104(decipher_0_i32box_ce104),
    .q104(decipher_0_i32box_q104),
    .address105(decipher_0_i32box_address105),
    .ce105(decipher_0_i32box_ce105),
    .q105(decipher_0_i32box_q105),
    .address106(decipher_0_i32box_address106),
    .ce106(decipher_0_i32box_ce106),
    .q106(decipher_0_i32box_q106),
    .address107(decipher_0_i32box_address107),
    .ce107(decipher_0_i32box_ce107),
    .q107(decipher_0_i32box_q107),
    .address108(decipher_0_i32box_address108),
    .ce108(decipher_0_i32box_ce108),
    .q108(decipher_0_i32box_q108),
    .address109(decipher_0_i32box_address109),
    .ce109(decipher_0_i32box_ce109),
    .q109(decipher_0_i32box_q109),
    .address110(decipher_0_i32box_address110),
    .ce110(decipher_0_i32box_ce110),
    .q110(decipher_0_i32box_q110),
    .address111(decipher_0_i32box_address111),
    .ce111(decipher_0_i32box_ce111),
    .q111(decipher_0_i32box_q111),
    .address112(decipher_0_i32box_address112),
    .ce112(decipher_0_i32box_ce112),
    .q112(decipher_0_i32box_q112),
    .address113(decipher_0_i32box_address113),
    .ce113(decipher_0_i32box_ce113),
    .q113(decipher_0_i32box_q113),
    .address114(decipher_0_i32box_address114),
    .ce114(decipher_0_i32box_ce114),
    .q114(decipher_0_i32box_q114),
    .address115(decipher_0_i32box_address115),
    .ce115(decipher_0_i32box_ce115),
    .q115(decipher_0_i32box_q115),
    .address116(decipher_0_i32box_address116),
    .ce116(decipher_0_i32box_ce116),
    .q116(decipher_0_i32box_q116),
    .address117(decipher_0_i32box_address117),
    .ce117(decipher_0_i32box_ce117),
    .q117(decipher_0_i32box_q117),
    .address118(decipher_0_i32box_address118),
    .ce118(decipher_0_i32box_ce118),
    .q118(decipher_0_i32box_q118),
    .address119(decipher_0_i32box_address119),
    .ce119(decipher_0_i32box_ce119),
    .q119(decipher_0_i32box_q119),
    .address120(decipher_0_i32box_address120),
    .ce120(decipher_0_i32box_ce120),
    .q120(decipher_0_i32box_q120),
    .address121(decipher_0_i32box_address121),
    .ce121(decipher_0_i32box_ce121),
    .q121(decipher_0_i32box_q121),
    .address122(decipher_0_i32box_address122),
    .ce122(decipher_0_i32box_ce122),
    .q122(decipher_0_i32box_q122),
    .address123(decipher_0_i32box_address123),
    .ce123(decipher_0_i32box_ce123),
    .q123(decipher_0_i32box_q123),
    .address124(decipher_0_i32box_address124),
    .ce124(decipher_0_i32box_ce124),
    .q124(decipher_0_i32box_q124),
    .address125(decipher_0_i32box_address125),
    .ce125(decipher_0_i32box_ce125),
    .q125(decipher_0_i32box_q125),
    .address126(decipher_0_i32box_address126),
    .ce126(decipher_0_i32box_ce126),
    .q126(decipher_0_i32box_q126),
    .address127(decipher_0_i32box_address127),
    .ce127(decipher_0_i32box_ce127),
    .q127(decipher_0_i32box_q127),
    .address128(decipher_0_i32box_address128),
    .ce128(decipher_0_i32box_ce128),
    .q128(decipher_0_i32box_q128),
    .address129(decipher_0_i32box_address129),
    .ce129(decipher_0_i32box_ce129),
    .q129(decipher_0_i32box_q129),
    .address130(decipher_0_i32box_address130),
    .ce130(decipher_0_i32box_ce130),
    .q130(decipher_0_i32box_q130),
    .address131(decipher_0_i32box_address131),
    .ce131(decipher_0_i32box_ce131),
    .q131(decipher_0_i32box_q131),
    .address132(decipher_0_i32box_address132),
    .ce132(decipher_0_i32box_ce132),
    .q132(decipher_0_i32box_q132),
    .address133(decipher_0_i32box_address133),
    .ce133(decipher_0_i32box_ce133),
    .q133(decipher_0_i32box_q133),
    .address134(decipher_0_i32box_address134),
    .ce134(decipher_0_i32box_ce134),
    .q134(decipher_0_i32box_q134),
    .address135(decipher_0_i32box_address135),
    .ce135(decipher_0_i32box_ce135),
    .q135(decipher_0_i32box_q135),
    .address136(decipher_0_i32box_address136),
    .ce136(decipher_0_i32box_ce136),
    .q136(decipher_0_i32box_q136),
    .address137(decipher_0_i32box_address137),
    .ce137(decipher_0_i32box_ce137),
    .q137(decipher_0_i32box_q137),
    .address138(decipher_0_i32box_address138),
    .ce138(decipher_0_i32box_ce138),
    .q138(decipher_0_i32box_q138),
    .address139(decipher_0_i32box_address139),
    .ce139(decipher_0_i32box_ce139),
    .q139(decipher_0_i32box_q139),
    .address140(decipher_0_i32box_address140),
    .ce140(decipher_0_i32box_ce140),
    .q140(decipher_0_i32box_q140),
    .address141(decipher_0_i32box_address141),
    .ce141(decipher_0_i32box_ce141),
    .q141(decipher_0_i32box_q141),
    .address142(decipher_0_i32box_address142),
    .ce142(decipher_0_i32box_ce142),
    .q142(decipher_0_i32box_q142),
    .address143(decipher_0_i32box_address143),
    .ce143(decipher_0_i32box_ce143),
    .q143(decipher_0_i32box_q143),
    .address144(decipher_0_i32box_address144),
    .ce144(decipher_0_i32box_ce144),
    .q144(decipher_0_i32box_q144),
    .address145(decipher_0_i32box_address145),
    .ce145(decipher_0_i32box_ce145),
    .q145(decipher_0_i32box_q145),
    .address146(decipher_0_i32box_address146),
    .ce146(decipher_0_i32box_ce146),
    .q146(decipher_0_i32box_q146),
    .address147(decipher_0_i32box_address147),
    .ce147(decipher_0_i32box_ce147),
    .q147(decipher_0_i32box_q147),
    .address148(decipher_0_i32box_address148),
    .ce148(decipher_0_i32box_ce148),
    .q148(decipher_0_i32box_q148),
    .address149(decipher_0_i32box_address149),
    .ce149(decipher_0_i32box_ce149),
    .q149(decipher_0_i32box_q149),
    .address150(decipher_0_i32box_address150),
    .ce150(decipher_0_i32box_ce150),
    .q150(decipher_0_i32box_q150),
    .address151(decipher_0_i32box_address151),
    .ce151(decipher_0_i32box_ce151),
    .q151(decipher_0_i32box_q151),
    .address152(decipher_0_i32box_address152),
    .ce152(decipher_0_i32box_ce152),
    .q152(decipher_0_i32box_q152),
    .address153(decipher_0_i32box_address153),
    .ce153(decipher_0_i32box_ce153),
    .q153(decipher_0_i32box_q153),
    .address154(decipher_0_i32box_address154),
    .ce154(decipher_0_i32box_ce154),
    .q154(decipher_0_i32box_q154),
    .address155(decipher_0_i32box_address155),
    .ce155(decipher_0_i32box_ce155),
    .q155(decipher_0_i32box_q155),
    .address156(decipher_0_i32box_address156),
    .ce156(decipher_0_i32box_ce156),
    .q156(decipher_0_i32box_q156),
    .address157(decipher_0_i32box_address157),
    .ce157(decipher_0_i32box_ce157),
    .q157(decipher_0_i32box_q157),
    .address158(decipher_0_i32box_address158),
    .ce158(decipher_0_i32box_ce158),
    .q158(decipher_0_i32box_q158),
    .address159(decipher_0_i32box_address159),
    .ce159(decipher_0_i32box_ce159),
    .q159(decipher_0_i32box_q159),
    .address160(decipher_0_i32box_address160),
    .ce160(decipher_0_i32box_ce160),
    .q160(decipher_0_i32box_q160),
    .address161(decipher_0_i32box_address161),
    .ce161(decipher_0_i32box_ce161),
    .q161(decipher_0_i32box_q161),
    .address162(decipher_0_i32box_address162),
    .ce162(decipher_0_i32box_ce162),
    .q162(decipher_0_i32box_q162),
    .address163(decipher_0_i32box_address163),
    .ce163(decipher_0_i32box_ce163),
    .q163(decipher_0_i32box_q163),
    .address164(decipher_0_i32box_address164),
    .ce164(decipher_0_i32box_ce164),
    .q164(decipher_0_i32box_q164),
    .address165(decipher_0_i32box_address165),
    .ce165(decipher_0_i32box_ce165),
    .q165(decipher_0_i32box_q165),
    .address166(decipher_0_i32box_address166),
    .ce166(decipher_0_i32box_ce166),
    .q166(decipher_0_i32box_q166),
    .address167(decipher_0_i32box_address167),
    .ce167(decipher_0_i32box_ce167),
    .q167(decipher_0_i32box_q167),
    .address168(decipher_0_i32box_address168),
    .ce168(decipher_0_i32box_ce168),
    .q168(decipher_0_i32box_q168),
    .address169(decipher_0_i32box_address169),
    .ce169(decipher_0_i32box_ce169),
    .q169(decipher_0_i32box_q169),
    .address170(decipher_0_i32box_address170),
    .ce170(decipher_0_i32box_ce170),
    .q170(decipher_0_i32box_q170),
    .address171(decipher_0_i32box_address171),
    .ce171(decipher_0_i32box_ce171),
    .q171(decipher_0_i32box_q171),
    .address172(decipher_0_i32box_address172),
    .ce172(decipher_0_i32box_ce172),
    .q172(decipher_0_i32box_q172),
    .address173(decipher_0_i32box_address173),
    .ce173(decipher_0_i32box_ce173),
    .q173(decipher_0_i32box_q173),
    .address174(decipher_0_i32box_address174),
    .ce174(decipher_0_i32box_ce174),
    .q174(decipher_0_i32box_q174),
    .address175(decipher_0_i32box_address175),
    .ce175(decipher_0_i32box_ce175),
    .q175(decipher_0_i32box_q175)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_enable_reg_pp0_iter1 <= ap_start;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter10 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter10 <= ap_enable_reg_pp0_iter9;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter11 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter11 <= ap_enable_reg_pp0_iter10;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter12 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter12 <= ap_enable_reg_pp0_iter11;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter13 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter13 <= ap_enable_reg_pp0_iter12;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter14 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter14 <= ap_enable_reg_pp0_iter13;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter15 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter15 <= ap_enable_reg_pp0_iter14;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter16 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter16 <= ap_enable_reg_pp0_iter15;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter17 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter17 <= ap_enable_reg_pp0_iter16;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter18 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter18 <= ap_enable_reg_pp0_iter17;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter19 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter19 <= ap_enable_reg_pp0_iter18;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter20 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter20 <= ap_enable_reg_pp0_iter19;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter21 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter21 <= ap_enable_reg_pp0_iter20;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter22 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter22 <= ap_enable_reg_pp0_iter21;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter23 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter23 <= ap_enable_reg_pp0_iter22;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter5 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter6 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter7 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter8 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter8 <= ap_enable_reg_pp0_iter7;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter9 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter9 <= ap_enable_reg_pp0_iter8;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        p_read13_reg_18005 <= p_read;
        p_read13_reg_18005_pp0_iter1_reg <= p_read13_reg_18005;
        p_read_10_reg_17990 <= p_read3;
        p_read_10_reg_17990_pp0_iter1_reg <= p_read_10_reg_17990;
        p_read_11_reg_17995 <= p_read2;
        p_read_11_reg_17995_pp0_iter1_reg <= p_read_11_reg_17995;
        p_read_12_reg_18000 <= p_read1;
        p_read_12_reg_18000_pp0_iter1_reg <= p_read_12_reg_18000;
        p_read_2_reg_17950 <= p_read11;
        p_read_3_reg_17955 <= p_read10;
        p_read_3_reg_17955_pp0_iter1_reg <= p_read_3_reg_17955;
        p_read_4_reg_17960 <= p_read9;
        p_read_4_reg_17960_pp0_iter1_reg <= p_read_4_reg_17960;
        p_read_5_reg_17965 <= p_read8;
        p_read_5_reg_17965_pp0_iter1_reg <= p_read_5_reg_17965;
        p_read_6_reg_17970 <= p_read7;
        p_read_6_reg_17970_pp0_iter1_reg <= p_read_6_reg_17970;
        p_read_7_reg_17975 <= p_read6;
        p_read_7_reg_17975_pp0_iter1_reg <= p_read_7_reg_17975;
        p_read_8_reg_17980 <= p_read5;
        p_read_8_reg_17980_pp0_iter1_reg <= p_read_8_reg_17980;
        p_read_9_reg_17985 <= p_read4;
        p_read_9_reg_17985_pp0_iter1_reg <= p_read_9_reg_17985;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        p_read13_reg_18005_pp0_iter10_reg <= p_read13_reg_18005_pp0_iter9_reg;
        p_read13_reg_18005_pp0_iter11_reg <= p_read13_reg_18005_pp0_iter10_reg;
        p_read13_reg_18005_pp0_iter12_reg <= p_read13_reg_18005_pp0_iter11_reg;
        p_read13_reg_18005_pp0_iter13_reg <= p_read13_reg_18005_pp0_iter12_reg;
        p_read13_reg_18005_pp0_iter14_reg <= p_read13_reg_18005_pp0_iter13_reg;
        p_read13_reg_18005_pp0_iter15_reg <= p_read13_reg_18005_pp0_iter14_reg;
        p_read13_reg_18005_pp0_iter16_reg <= p_read13_reg_18005_pp0_iter15_reg;
        p_read13_reg_18005_pp0_iter17_reg <= p_read13_reg_18005_pp0_iter16_reg;
        p_read13_reg_18005_pp0_iter18_reg <= p_read13_reg_18005_pp0_iter17_reg;
        p_read13_reg_18005_pp0_iter19_reg <= p_read13_reg_18005_pp0_iter18_reg;
        p_read13_reg_18005_pp0_iter20_reg <= p_read13_reg_18005_pp0_iter19_reg;
        p_read13_reg_18005_pp0_iter21_reg <= p_read13_reg_18005_pp0_iter20_reg;
        p_read13_reg_18005_pp0_iter22_reg <= p_read13_reg_18005_pp0_iter21_reg;
        p_read13_reg_18005_pp0_iter2_reg <= p_read13_reg_18005_pp0_iter1_reg;
        p_read13_reg_18005_pp0_iter3_reg <= p_read13_reg_18005_pp0_iter2_reg;
        p_read13_reg_18005_pp0_iter4_reg <= p_read13_reg_18005_pp0_iter3_reg;
        p_read13_reg_18005_pp0_iter5_reg <= p_read13_reg_18005_pp0_iter4_reg;
        p_read13_reg_18005_pp0_iter6_reg <= p_read13_reg_18005_pp0_iter5_reg;
        p_read13_reg_18005_pp0_iter7_reg <= p_read13_reg_18005_pp0_iter6_reg;
        p_read13_reg_18005_pp0_iter8_reg <= p_read13_reg_18005_pp0_iter7_reg;
        p_read13_reg_18005_pp0_iter9_reg <= p_read13_reg_18005_pp0_iter8_reg;
        p_read_10_reg_17990_pp0_iter10_reg <= p_read_10_reg_17990_pp0_iter9_reg;
        p_read_10_reg_17990_pp0_iter11_reg <= p_read_10_reg_17990_pp0_iter10_reg;
        p_read_10_reg_17990_pp0_iter12_reg <= p_read_10_reg_17990_pp0_iter11_reg;
        p_read_10_reg_17990_pp0_iter13_reg <= p_read_10_reg_17990_pp0_iter12_reg;
        p_read_10_reg_17990_pp0_iter14_reg <= p_read_10_reg_17990_pp0_iter13_reg;
        p_read_10_reg_17990_pp0_iter15_reg <= p_read_10_reg_17990_pp0_iter14_reg;
        p_read_10_reg_17990_pp0_iter16_reg <= p_read_10_reg_17990_pp0_iter15_reg;
        p_read_10_reg_17990_pp0_iter2_reg <= p_read_10_reg_17990_pp0_iter1_reg;
        p_read_10_reg_17990_pp0_iter3_reg <= p_read_10_reg_17990_pp0_iter2_reg;
        p_read_10_reg_17990_pp0_iter4_reg <= p_read_10_reg_17990_pp0_iter3_reg;
        p_read_10_reg_17990_pp0_iter5_reg <= p_read_10_reg_17990_pp0_iter4_reg;
        p_read_10_reg_17990_pp0_iter6_reg <= p_read_10_reg_17990_pp0_iter5_reg;
        p_read_10_reg_17990_pp0_iter7_reg <= p_read_10_reg_17990_pp0_iter6_reg;
        p_read_10_reg_17990_pp0_iter8_reg <= p_read_10_reg_17990_pp0_iter7_reg;
        p_read_10_reg_17990_pp0_iter9_reg <= p_read_10_reg_17990_pp0_iter8_reg;
        p_read_11_reg_17995_pp0_iter10_reg <= p_read_11_reg_17995_pp0_iter9_reg;
        p_read_11_reg_17995_pp0_iter11_reg <= p_read_11_reg_17995_pp0_iter10_reg;
        p_read_11_reg_17995_pp0_iter12_reg <= p_read_11_reg_17995_pp0_iter11_reg;
        p_read_11_reg_17995_pp0_iter13_reg <= p_read_11_reg_17995_pp0_iter12_reg;
        p_read_11_reg_17995_pp0_iter14_reg <= p_read_11_reg_17995_pp0_iter13_reg;
        p_read_11_reg_17995_pp0_iter15_reg <= p_read_11_reg_17995_pp0_iter14_reg;
        p_read_11_reg_17995_pp0_iter16_reg <= p_read_11_reg_17995_pp0_iter15_reg;
        p_read_11_reg_17995_pp0_iter17_reg <= p_read_11_reg_17995_pp0_iter16_reg;
        p_read_11_reg_17995_pp0_iter18_reg <= p_read_11_reg_17995_pp0_iter17_reg;
        p_read_11_reg_17995_pp0_iter2_reg <= p_read_11_reg_17995_pp0_iter1_reg;
        p_read_11_reg_17995_pp0_iter3_reg <= p_read_11_reg_17995_pp0_iter2_reg;
        p_read_11_reg_17995_pp0_iter4_reg <= p_read_11_reg_17995_pp0_iter3_reg;
        p_read_11_reg_17995_pp0_iter5_reg <= p_read_11_reg_17995_pp0_iter4_reg;
        p_read_11_reg_17995_pp0_iter6_reg <= p_read_11_reg_17995_pp0_iter5_reg;
        p_read_11_reg_17995_pp0_iter7_reg <= p_read_11_reg_17995_pp0_iter6_reg;
        p_read_11_reg_17995_pp0_iter8_reg <= p_read_11_reg_17995_pp0_iter7_reg;
        p_read_11_reg_17995_pp0_iter9_reg <= p_read_11_reg_17995_pp0_iter8_reg;
        p_read_12_reg_18000_pp0_iter10_reg <= p_read_12_reg_18000_pp0_iter9_reg;
        p_read_12_reg_18000_pp0_iter11_reg <= p_read_12_reg_18000_pp0_iter10_reg;
        p_read_12_reg_18000_pp0_iter12_reg <= p_read_12_reg_18000_pp0_iter11_reg;
        p_read_12_reg_18000_pp0_iter13_reg <= p_read_12_reg_18000_pp0_iter12_reg;
        p_read_12_reg_18000_pp0_iter14_reg <= p_read_12_reg_18000_pp0_iter13_reg;
        p_read_12_reg_18000_pp0_iter15_reg <= p_read_12_reg_18000_pp0_iter14_reg;
        p_read_12_reg_18000_pp0_iter16_reg <= p_read_12_reg_18000_pp0_iter15_reg;
        p_read_12_reg_18000_pp0_iter17_reg <= p_read_12_reg_18000_pp0_iter16_reg;
        p_read_12_reg_18000_pp0_iter18_reg <= p_read_12_reg_18000_pp0_iter17_reg;
        p_read_12_reg_18000_pp0_iter19_reg <= p_read_12_reg_18000_pp0_iter18_reg;
        p_read_12_reg_18000_pp0_iter20_reg <= p_read_12_reg_18000_pp0_iter19_reg;
        p_read_12_reg_18000_pp0_iter2_reg <= p_read_12_reg_18000_pp0_iter1_reg;
        p_read_12_reg_18000_pp0_iter3_reg <= p_read_12_reg_18000_pp0_iter2_reg;
        p_read_12_reg_18000_pp0_iter4_reg <= p_read_12_reg_18000_pp0_iter3_reg;
        p_read_12_reg_18000_pp0_iter5_reg <= p_read_12_reg_18000_pp0_iter4_reg;
        p_read_12_reg_18000_pp0_iter6_reg <= p_read_12_reg_18000_pp0_iter5_reg;
        p_read_12_reg_18000_pp0_iter7_reg <= p_read_12_reg_18000_pp0_iter6_reg;
        p_read_12_reg_18000_pp0_iter8_reg <= p_read_12_reg_18000_pp0_iter7_reg;
        p_read_12_reg_18000_pp0_iter9_reg <= p_read_12_reg_18000_pp0_iter8_reg;
        p_read_3_reg_17955_pp0_iter2_reg <= p_read_3_reg_17955_pp0_iter1_reg;
        p_read_4_reg_17960_pp0_iter2_reg <= p_read_4_reg_17960_pp0_iter1_reg;
        p_read_4_reg_17960_pp0_iter3_reg <= p_read_4_reg_17960_pp0_iter2_reg;
        p_read_4_reg_17960_pp0_iter4_reg <= p_read_4_reg_17960_pp0_iter3_reg;
        p_read_5_reg_17965_pp0_iter2_reg <= p_read_5_reg_17965_pp0_iter1_reg;
        p_read_5_reg_17965_pp0_iter3_reg <= p_read_5_reg_17965_pp0_iter2_reg;
        p_read_5_reg_17965_pp0_iter4_reg <= p_read_5_reg_17965_pp0_iter3_reg;
        p_read_5_reg_17965_pp0_iter5_reg <= p_read_5_reg_17965_pp0_iter4_reg;
        p_read_5_reg_17965_pp0_iter6_reg <= p_read_5_reg_17965_pp0_iter5_reg;
        p_read_6_reg_17970_pp0_iter2_reg <= p_read_6_reg_17970_pp0_iter1_reg;
        p_read_6_reg_17970_pp0_iter3_reg <= p_read_6_reg_17970_pp0_iter2_reg;
        p_read_6_reg_17970_pp0_iter4_reg <= p_read_6_reg_17970_pp0_iter3_reg;
        p_read_6_reg_17970_pp0_iter5_reg <= p_read_6_reg_17970_pp0_iter4_reg;
        p_read_6_reg_17970_pp0_iter6_reg <= p_read_6_reg_17970_pp0_iter5_reg;
        p_read_6_reg_17970_pp0_iter7_reg <= p_read_6_reg_17970_pp0_iter6_reg;
        p_read_6_reg_17970_pp0_iter8_reg <= p_read_6_reg_17970_pp0_iter7_reg;
        p_read_7_reg_17975_pp0_iter10_reg <= p_read_7_reg_17975_pp0_iter9_reg;
        p_read_7_reg_17975_pp0_iter2_reg <= p_read_7_reg_17975_pp0_iter1_reg;
        p_read_7_reg_17975_pp0_iter3_reg <= p_read_7_reg_17975_pp0_iter2_reg;
        p_read_7_reg_17975_pp0_iter4_reg <= p_read_7_reg_17975_pp0_iter3_reg;
        p_read_7_reg_17975_pp0_iter5_reg <= p_read_7_reg_17975_pp0_iter4_reg;
        p_read_7_reg_17975_pp0_iter6_reg <= p_read_7_reg_17975_pp0_iter5_reg;
        p_read_7_reg_17975_pp0_iter7_reg <= p_read_7_reg_17975_pp0_iter6_reg;
        p_read_7_reg_17975_pp0_iter8_reg <= p_read_7_reg_17975_pp0_iter7_reg;
        p_read_7_reg_17975_pp0_iter9_reg <= p_read_7_reg_17975_pp0_iter8_reg;
        p_read_8_reg_17980_pp0_iter10_reg <= p_read_8_reg_17980_pp0_iter9_reg;
        p_read_8_reg_17980_pp0_iter11_reg <= p_read_8_reg_17980_pp0_iter10_reg;
        p_read_8_reg_17980_pp0_iter12_reg <= p_read_8_reg_17980_pp0_iter11_reg;
        p_read_8_reg_17980_pp0_iter2_reg <= p_read_8_reg_17980_pp0_iter1_reg;
        p_read_8_reg_17980_pp0_iter3_reg <= p_read_8_reg_17980_pp0_iter2_reg;
        p_read_8_reg_17980_pp0_iter4_reg <= p_read_8_reg_17980_pp0_iter3_reg;
        p_read_8_reg_17980_pp0_iter5_reg <= p_read_8_reg_17980_pp0_iter4_reg;
        p_read_8_reg_17980_pp0_iter6_reg <= p_read_8_reg_17980_pp0_iter5_reg;
        p_read_8_reg_17980_pp0_iter7_reg <= p_read_8_reg_17980_pp0_iter6_reg;
        p_read_8_reg_17980_pp0_iter8_reg <= p_read_8_reg_17980_pp0_iter7_reg;
        p_read_8_reg_17980_pp0_iter9_reg <= p_read_8_reg_17980_pp0_iter8_reg;
        p_read_9_reg_17985_pp0_iter10_reg <= p_read_9_reg_17985_pp0_iter9_reg;
        p_read_9_reg_17985_pp0_iter11_reg <= p_read_9_reg_17985_pp0_iter10_reg;
        p_read_9_reg_17985_pp0_iter12_reg <= p_read_9_reg_17985_pp0_iter11_reg;
        p_read_9_reg_17985_pp0_iter13_reg <= p_read_9_reg_17985_pp0_iter12_reg;
        p_read_9_reg_17985_pp0_iter14_reg <= p_read_9_reg_17985_pp0_iter13_reg;
        p_read_9_reg_17985_pp0_iter2_reg <= p_read_9_reg_17985_pp0_iter1_reg;
        p_read_9_reg_17985_pp0_iter3_reg <= p_read_9_reg_17985_pp0_iter2_reg;
        p_read_9_reg_17985_pp0_iter4_reg <= p_read_9_reg_17985_pp0_iter3_reg;
        p_read_9_reg_17985_pp0_iter5_reg <= p_read_9_reg_17985_pp0_iter4_reg;
        p_read_9_reg_17985_pp0_iter6_reg <= p_read_9_reg_17985_pp0_iter5_reg;
        p_read_9_reg_17985_pp0_iter7_reg <= p_read_9_reg_17985_pp0_iter6_reg;
        p_read_9_reg_17985_pp0_iter8_reg <= p_read_9_reg_17985_pp0_iter7_reg;
        p_read_9_reg_17985_pp0_iter9_reg <= p_read_9_reg_17985_pp0_iter8_reg;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter23 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_idle_pp0 == 1'b1) & (ap_start == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter23 == 1'b0) & (ap_enable_reg_pp0_iter22 == 1'b0) & (ap_enable_reg_pp0_iter21 == 1'b0) & (ap_enable_reg_pp0_iter20 == 1'b0) & (ap_enable_reg_pp0_iter19 == 1'b0) & (ap_enable_reg_pp0_iter18 == 1'b0) & (ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b0) & (ap_enable_reg_pp0_iter21 == 1'b0) & (ap_enable_reg_pp0_iter20 == 1'b0) & (ap_enable_reg_pp0_iter19 == 1'b0) & (ap_enable_reg_pp0_iter18 == 1'b0) & (ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0_0to22 = 1'b1;
    end else begin
        ap_idle_pp0_0to22 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (ap_idle_pp0_0to22 == 1'b1))) begin
        ap_reset_idle_pp0 = 1'b1;
    end else begin
        ap_reset_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce0 = 1'b1;
    end else begin
        decipher_0_i32box_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce1 = 1'b1;
    end else begin
        decipher_0_i32box_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce10 = 1'b1;
    end else begin
        decipher_0_i32box_ce10 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce100 = 1'b1;
    end else begin
        decipher_0_i32box_ce100 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce101 = 1'b1;
    end else begin
        decipher_0_i32box_ce101 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce102 = 1'b1;
    end else begin
        decipher_0_i32box_ce102 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce103 = 1'b1;
    end else begin
        decipher_0_i32box_ce103 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce104 = 1'b1;
    end else begin
        decipher_0_i32box_ce104 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce105 = 1'b1;
    end else begin
        decipher_0_i32box_ce105 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce106 = 1'b1;
    end else begin
        decipher_0_i32box_ce106 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce107 = 1'b1;
    end else begin
        decipher_0_i32box_ce107 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce108 = 1'b1;
    end else begin
        decipher_0_i32box_ce108 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce109 = 1'b1;
    end else begin
        decipher_0_i32box_ce109 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce11 = 1'b1;
    end else begin
        decipher_0_i32box_ce11 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce110 = 1'b1;
    end else begin
        decipher_0_i32box_ce110 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce111 = 1'b1;
    end else begin
        decipher_0_i32box_ce111 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce112 = 1'b1;
    end else begin
        decipher_0_i32box_ce112 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce113 = 1'b1;
    end else begin
        decipher_0_i32box_ce113 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce114 = 1'b1;
    end else begin
        decipher_0_i32box_ce114 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce115 = 1'b1;
    end else begin
        decipher_0_i32box_ce115 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce116 = 1'b1;
    end else begin
        decipher_0_i32box_ce116 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce117 = 1'b1;
    end else begin
        decipher_0_i32box_ce117 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce118 = 1'b1;
    end else begin
        decipher_0_i32box_ce118 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce119 = 1'b1;
    end else begin
        decipher_0_i32box_ce119 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce12 = 1'b1;
    end else begin
        decipher_0_i32box_ce12 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce120 = 1'b1;
    end else begin
        decipher_0_i32box_ce120 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce121 = 1'b1;
    end else begin
        decipher_0_i32box_ce121 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce122 = 1'b1;
    end else begin
        decipher_0_i32box_ce122 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce123 = 1'b1;
    end else begin
        decipher_0_i32box_ce123 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce124 = 1'b1;
    end else begin
        decipher_0_i32box_ce124 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce125 = 1'b1;
    end else begin
        decipher_0_i32box_ce125 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce126 = 1'b1;
    end else begin
        decipher_0_i32box_ce126 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce127 = 1'b1;
    end else begin
        decipher_0_i32box_ce127 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce128 = 1'b1;
    end else begin
        decipher_0_i32box_ce128 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce129 = 1'b1;
    end else begin
        decipher_0_i32box_ce129 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce13 = 1'b1;
    end else begin
        decipher_0_i32box_ce13 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce130 = 1'b1;
    end else begin
        decipher_0_i32box_ce130 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce131 = 1'b1;
    end else begin
        decipher_0_i32box_ce131 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce132 = 1'b1;
    end else begin
        decipher_0_i32box_ce132 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce133 = 1'b1;
    end else begin
        decipher_0_i32box_ce133 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce134 = 1'b1;
    end else begin
        decipher_0_i32box_ce134 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce135 = 1'b1;
    end else begin
        decipher_0_i32box_ce135 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce136 = 1'b1;
    end else begin
        decipher_0_i32box_ce136 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce137 = 1'b1;
    end else begin
        decipher_0_i32box_ce137 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce138 = 1'b1;
    end else begin
        decipher_0_i32box_ce138 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce139 = 1'b1;
    end else begin
        decipher_0_i32box_ce139 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce14 = 1'b1;
    end else begin
        decipher_0_i32box_ce14 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce140 = 1'b1;
    end else begin
        decipher_0_i32box_ce140 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce141 = 1'b1;
    end else begin
        decipher_0_i32box_ce141 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce142 = 1'b1;
    end else begin
        decipher_0_i32box_ce142 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce143 = 1'b1;
    end else begin
        decipher_0_i32box_ce143 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce144 = 1'b1;
    end else begin
        decipher_0_i32box_ce144 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce145 = 1'b1;
    end else begin
        decipher_0_i32box_ce145 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce146 = 1'b1;
    end else begin
        decipher_0_i32box_ce146 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce147 = 1'b1;
    end else begin
        decipher_0_i32box_ce147 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce148 = 1'b1;
    end else begin
        decipher_0_i32box_ce148 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce149 = 1'b1;
    end else begin
        decipher_0_i32box_ce149 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce15 = 1'b1;
    end else begin
        decipher_0_i32box_ce15 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce150 = 1'b1;
    end else begin
        decipher_0_i32box_ce150 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce151 = 1'b1;
    end else begin
        decipher_0_i32box_ce151 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce152 = 1'b1;
    end else begin
        decipher_0_i32box_ce152 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce153 = 1'b1;
    end else begin
        decipher_0_i32box_ce153 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce154 = 1'b1;
    end else begin
        decipher_0_i32box_ce154 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce155 = 1'b1;
    end else begin
        decipher_0_i32box_ce155 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce156 = 1'b1;
    end else begin
        decipher_0_i32box_ce156 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce157 = 1'b1;
    end else begin
        decipher_0_i32box_ce157 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce158 = 1'b1;
    end else begin
        decipher_0_i32box_ce158 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce159 = 1'b1;
    end else begin
        decipher_0_i32box_ce159 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce16 = 1'b1;
    end else begin
        decipher_0_i32box_ce16 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce160 = 1'b1;
    end else begin
        decipher_0_i32box_ce160 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce161 = 1'b1;
    end else begin
        decipher_0_i32box_ce161 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce162 = 1'b1;
    end else begin
        decipher_0_i32box_ce162 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce163 = 1'b1;
    end else begin
        decipher_0_i32box_ce163 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce164 = 1'b1;
    end else begin
        decipher_0_i32box_ce164 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce165 = 1'b1;
    end else begin
        decipher_0_i32box_ce165 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce166 = 1'b1;
    end else begin
        decipher_0_i32box_ce166 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce167 = 1'b1;
    end else begin
        decipher_0_i32box_ce167 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce168 = 1'b1;
    end else begin
        decipher_0_i32box_ce168 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce169 = 1'b1;
    end else begin
        decipher_0_i32box_ce169 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce17 = 1'b1;
    end else begin
        decipher_0_i32box_ce17 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce170 = 1'b1;
    end else begin
        decipher_0_i32box_ce170 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce171 = 1'b1;
    end else begin
        decipher_0_i32box_ce171 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce172 = 1'b1;
    end else begin
        decipher_0_i32box_ce172 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce173 = 1'b1;
    end else begin
        decipher_0_i32box_ce173 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce174 = 1'b1;
    end else begin
        decipher_0_i32box_ce174 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce175 = 1'b1;
    end else begin
        decipher_0_i32box_ce175 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce18 = 1'b1;
    end else begin
        decipher_0_i32box_ce18 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce19 = 1'b1;
    end else begin
        decipher_0_i32box_ce19 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce2 = 1'b1;
    end else begin
        decipher_0_i32box_ce2 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce20 = 1'b1;
    end else begin
        decipher_0_i32box_ce20 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce21 = 1'b1;
    end else begin
        decipher_0_i32box_ce21 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce22 = 1'b1;
    end else begin
        decipher_0_i32box_ce22 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce23 = 1'b1;
    end else begin
        decipher_0_i32box_ce23 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce24 = 1'b1;
    end else begin
        decipher_0_i32box_ce24 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce25 = 1'b1;
    end else begin
        decipher_0_i32box_ce25 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce26 = 1'b1;
    end else begin
        decipher_0_i32box_ce26 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce27 = 1'b1;
    end else begin
        decipher_0_i32box_ce27 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce28 = 1'b1;
    end else begin
        decipher_0_i32box_ce28 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce29 = 1'b1;
    end else begin
        decipher_0_i32box_ce29 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce3 = 1'b1;
    end else begin
        decipher_0_i32box_ce3 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce30 = 1'b1;
    end else begin
        decipher_0_i32box_ce30 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce31 = 1'b1;
    end else begin
        decipher_0_i32box_ce31 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce32 = 1'b1;
    end else begin
        decipher_0_i32box_ce32 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce33 = 1'b1;
    end else begin
        decipher_0_i32box_ce33 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce34 = 1'b1;
    end else begin
        decipher_0_i32box_ce34 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce35 = 1'b1;
    end else begin
        decipher_0_i32box_ce35 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce36 = 1'b1;
    end else begin
        decipher_0_i32box_ce36 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce37 = 1'b1;
    end else begin
        decipher_0_i32box_ce37 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce38 = 1'b1;
    end else begin
        decipher_0_i32box_ce38 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce39 = 1'b1;
    end else begin
        decipher_0_i32box_ce39 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce4 = 1'b1;
    end else begin
        decipher_0_i32box_ce4 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce40 = 1'b1;
    end else begin
        decipher_0_i32box_ce40 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce41 = 1'b1;
    end else begin
        decipher_0_i32box_ce41 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce42 = 1'b1;
    end else begin
        decipher_0_i32box_ce42 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce43 = 1'b1;
    end else begin
        decipher_0_i32box_ce43 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce44 = 1'b1;
    end else begin
        decipher_0_i32box_ce44 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce45 = 1'b1;
    end else begin
        decipher_0_i32box_ce45 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce46 = 1'b1;
    end else begin
        decipher_0_i32box_ce46 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce47 = 1'b1;
    end else begin
        decipher_0_i32box_ce47 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce48 = 1'b1;
    end else begin
        decipher_0_i32box_ce48 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce49 = 1'b1;
    end else begin
        decipher_0_i32box_ce49 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce5 = 1'b1;
    end else begin
        decipher_0_i32box_ce5 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce50 = 1'b1;
    end else begin
        decipher_0_i32box_ce50 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce51 = 1'b1;
    end else begin
        decipher_0_i32box_ce51 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce52 = 1'b1;
    end else begin
        decipher_0_i32box_ce52 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce53 = 1'b1;
    end else begin
        decipher_0_i32box_ce53 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce54 = 1'b1;
    end else begin
        decipher_0_i32box_ce54 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce55 = 1'b1;
    end else begin
        decipher_0_i32box_ce55 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce56 = 1'b1;
    end else begin
        decipher_0_i32box_ce56 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce57 = 1'b1;
    end else begin
        decipher_0_i32box_ce57 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce58 = 1'b1;
    end else begin
        decipher_0_i32box_ce58 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce59 = 1'b1;
    end else begin
        decipher_0_i32box_ce59 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce6 = 1'b1;
    end else begin
        decipher_0_i32box_ce6 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce60 = 1'b1;
    end else begin
        decipher_0_i32box_ce60 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce61 = 1'b1;
    end else begin
        decipher_0_i32box_ce61 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce62 = 1'b1;
    end else begin
        decipher_0_i32box_ce62 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce63 = 1'b1;
    end else begin
        decipher_0_i32box_ce63 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce64 = 1'b1;
    end else begin
        decipher_0_i32box_ce64 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce65 = 1'b1;
    end else begin
        decipher_0_i32box_ce65 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce66 = 1'b1;
    end else begin
        decipher_0_i32box_ce66 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce67 = 1'b1;
    end else begin
        decipher_0_i32box_ce67 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce68 = 1'b1;
    end else begin
        decipher_0_i32box_ce68 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce69 = 1'b1;
    end else begin
        decipher_0_i32box_ce69 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce7 = 1'b1;
    end else begin
        decipher_0_i32box_ce7 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce70 = 1'b1;
    end else begin
        decipher_0_i32box_ce70 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce71 = 1'b1;
    end else begin
        decipher_0_i32box_ce71 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce72 = 1'b1;
    end else begin
        decipher_0_i32box_ce72 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce73 = 1'b1;
    end else begin
        decipher_0_i32box_ce73 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce74 = 1'b1;
    end else begin
        decipher_0_i32box_ce74 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce75 = 1'b1;
    end else begin
        decipher_0_i32box_ce75 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce76 = 1'b1;
    end else begin
        decipher_0_i32box_ce76 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce77 = 1'b1;
    end else begin
        decipher_0_i32box_ce77 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce78 = 1'b1;
    end else begin
        decipher_0_i32box_ce78 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce79 = 1'b1;
    end else begin
        decipher_0_i32box_ce79 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce8 = 1'b1;
    end else begin
        decipher_0_i32box_ce8 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce80 = 1'b1;
    end else begin
        decipher_0_i32box_ce80 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce81 = 1'b1;
    end else begin
        decipher_0_i32box_ce81 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce82 = 1'b1;
    end else begin
        decipher_0_i32box_ce82 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce83 = 1'b1;
    end else begin
        decipher_0_i32box_ce83 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce84 = 1'b1;
    end else begin
        decipher_0_i32box_ce84 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce85 = 1'b1;
    end else begin
        decipher_0_i32box_ce85 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce86 = 1'b1;
    end else begin
        decipher_0_i32box_ce86 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce87 = 1'b1;
    end else begin
        decipher_0_i32box_ce87 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce88 = 1'b1;
    end else begin
        decipher_0_i32box_ce88 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce89 = 1'b1;
    end else begin
        decipher_0_i32box_ce89 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce9 = 1'b1;
    end else begin
        decipher_0_i32box_ce9 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce90 = 1'b1;
    end else begin
        decipher_0_i32box_ce90 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce91 = 1'b1;
    end else begin
        decipher_0_i32box_ce91 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce92 = 1'b1;
    end else begin
        decipher_0_i32box_ce92 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce93 = 1'b1;
    end else begin
        decipher_0_i32box_ce93 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce94 = 1'b1;
    end else begin
        decipher_0_i32box_ce94 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce95 = 1'b1;
    end else begin
        decipher_0_i32box_ce95 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce96 = 1'b1;
    end else begin
        decipher_0_i32box_ce96 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce97 = 1'b1;
    end else begin
        decipher_0_i32box_ce97 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce98 = 1'b1;
    end else begin
        decipher_0_i32box_ce98 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce99 = 1'b1;
    end else begin
        decipher_0_i32box_ce99 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce0 = 1'b1;
    end else begin
        decipher_0_iibox_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce1 = 1'b1;
    end else begin
        decipher_0_iibox_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce10 = 1'b1;
    end else begin
        decipher_0_iibox_ce10 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce100 = 1'b1;
    end else begin
        decipher_0_iibox_ce100 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce101 = 1'b1;
    end else begin
        decipher_0_iibox_ce101 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce102 = 1'b1;
    end else begin
        decipher_0_iibox_ce102 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce103 = 1'b1;
    end else begin
        decipher_0_iibox_ce103 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce104 = 1'b1;
    end else begin
        decipher_0_iibox_ce104 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce105 = 1'b1;
    end else begin
        decipher_0_iibox_ce105 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce106 = 1'b1;
    end else begin
        decipher_0_iibox_ce106 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce107 = 1'b1;
    end else begin
        decipher_0_iibox_ce107 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce108 = 1'b1;
    end else begin
        decipher_0_iibox_ce108 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce109 = 1'b1;
    end else begin
        decipher_0_iibox_ce109 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce11 = 1'b1;
    end else begin
        decipher_0_iibox_ce11 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce110 = 1'b1;
    end else begin
        decipher_0_iibox_ce110 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce111 = 1'b1;
    end else begin
        decipher_0_iibox_ce111 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce112 = 1'b1;
    end else begin
        decipher_0_iibox_ce112 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce113 = 1'b1;
    end else begin
        decipher_0_iibox_ce113 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce114 = 1'b1;
    end else begin
        decipher_0_iibox_ce114 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce115 = 1'b1;
    end else begin
        decipher_0_iibox_ce115 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce116 = 1'b1;
    end else begin
        decipher_0_iibox_ce116 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce117 = 1'b1;
    end else begin
        decipher_0_iibox_ce117 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce118 = 1'b1;
    end else begin
        decipher_0_iibox_ce118 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce119 = 1'b1;
    end else begin
        decipher_0_iibox_ce119 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce12 = 1'b1;
    end else begin
        decipher_0_iibox_ce12 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce120 = 1'b1;
    end else begin
        decipher_0_iibox_ce120 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce121 = 1'b1;
    end else begin
        decipher_0_iibox_ce121 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce122 = 1'b1;
    end else begin
        decipher_0_iibox_ce122 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce123 = 1'b1;
    end else begin
        decipher_0_iibox_ce123 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce124 = 1'b1;
    end else begin
        decipher_0_iibox_ce124 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce125 = 1'b1;
    end else begin
        decipher_0_iibox_ce125 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce126 = 1'b1;
    end else begin
        decipher_0_iibox_ce126 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce127 = 1'b1;
    end else begin
        decipher_0_iibox_ce127 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce128 = 1'b1;
    end else begin
        decipher_0_iibox_ce128 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce129 = 1'b1;
    end else begin
        decipher_0_iibox_ce129 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce13 = 1'b1;
    end else begin
        decipher_0_iibox_ce13 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce130 = 1'b1;
    end else begin
        decipher_0_iibox_ce130 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce131 = 1'b1;
    end else begin
        decipher_0_iibox_ce131 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce132 = 1'b1;
    end else begin
        decipher_0_iibox_ce132 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce133 = 1'b1;
    end else begin
        decipher_0_iibox_ce133 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce134 = 1'b1;
    end else begin
        decipher_0_iibox_ce134 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce135 = 1'b1;
    end else begin
        decipher_0_iibox_ce135 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce136 = 1'b1;
    end else begin
        decipher_0_iibox_ce136 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce137 = 1'b1;
    end else begin
        decipher_0_iibox_ce137 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce138 = 1'b1;
    end else begin
        decipher_0_iibox_ce138 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce139 = 1'b1;
    end else begin
        decipher_0_iibox_ce139 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce14 = 1'b1;
    end else begin
        decipher_0_iibox_ce14 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce140 = 1'b1;
    end else begin
        decipher_0_iibox_ce140 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce141 = 1'b1;
    end else begin
        decipher_0_iibox_ce141 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce142 = 1'b1;
    end else begin
        decipher_0_iibox_ce142 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce143 = 1'b1;
    end else begin
        decipher_0_iibox_ce143 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce144 = 1'b1;
    end else begin
        decipher_0_iibox_ce144 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce145 = 1'b1;
    end else begin
        decipher_0_iibox_ce145 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce146 = 1'b1;
    end else begin
        decipher_0_iibox_ce146 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce147 = 1'b1;
    end else begin
        decipher_0_iibox_ce147 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce148 = 1'b1;
    end else begin
        decipher_0_iibox_ce148 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce149 = 1'b1;
    end else begin
        decipher_0_iibox_ce149 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce15 = 1'b1;
    end else begin
        decipher_0_iibox_ce15 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce150 = 1'b1;
    end else begin
        decipher_0_iibox_ce150 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce151 = 1'b1;
    end else begin
        decipher_0_iibox_ce151 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce152 = 1'b1;
    end else begin
        decipher_0_iibox_ce152 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce153 = 1'b1;
    end else begin
        decipher_0_iibox_ce153 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce154 = 1'b1;
    end else begin
        decipher_0_iibox_ce154 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce155 = 1'b1;
    end else begin
        decipher_0_iibox_ce155 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce156 = 1'b1;
    end else begin
        decipher_0_iibox_ce156 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce157 = 1'b1;
    end else begin
        decipher_0_iibox_ce157 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce158 = 1'b1;
    end else begin
        decipher_0_iibox_ce158 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce159 = 1'b1;
    end else begin
        decipher_0_iibox_ce159 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce16 = 1'b1;
    end else begin
        decipher_0_iibox_ce16 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce160 = 1'b1;
    end else begin
        decipher_0_iibox_ce160 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce161 = 1'b1;
    end else begin
        decipher_0_iibox_ce161 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce162 = 1'b1;
    end else begin
        decipher_0_iibox_ce162 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce163 = 1'b1;
    end else begin
        decipher_0_iibox_ce163 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce164 = 1'b1;
    end else begin
        decipher_0_iibox_ce164 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce165 = 1'b1;
    end else begin
        decipher_0_iibox_ce165 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce166 = 1'b1;
    end else begin
        decipher_0_iibox_ce166 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce167 = 1'b1;
    end else begin
        decipher_0_iibox_ce167 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce168 = 1'b1;
    end else begin
        decipher_0_iibox_ce168 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce169 = 1'b1;
    end else begin
        decipher_0_iibox_ce169 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce17 = 1'b1;
    end else begin
        decipher_0_iibox_ce17 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce170 = 1'b1;
    end else begin
        decipher_0_iibox_ce170 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce171 = 1'b1;
    end else begin
        decipher_0_iibox_ce171 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce172 = 1'b1;
    end else begin
        decipher_0_iibox_ce172 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce173 = 1'b1;
    end else begin
        decipher_0_iibox_ce173 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce174 = 1'b1;
    end else begin
        decipher_0_iibox_ce174 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce175 = 1'b1;
    end else begin
        decipher_0_iibox_ce175 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce176 = 1'b1;
    end else begin
        decipher_0_iibox_ce176 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce177 = 1'b1;
    end else begin
        decipher_0_iibox_ce177 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce178 = 1'b1;
    end else begin
        decipher_0_iibox_ce178 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce179 = 1'b1;
    end else begin
        decipher_0_iibox_ce179 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce18 = 1'b1;
    end else begin
        decipher_0_iibox_ce18 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce180 = 1'b1;
    end else begin
        decipher_0_iibox_ce180 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce181 = 1'b1;
    end else begin
        decipher_0_iibox_ce181 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce182 = 1'b1;
    end else begin
        decipher_0_iibox_ce182 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce183 = 1'b1;
    end else begin
        decipher_0_iibox_ce183 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce184 = 1'b1;
    end else begin
        decipher_0_iibox_ce184 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce185 = 1'b1;
    end else begin
        decipher_0_iibox_ce185 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce186 = 1'b1;
    end else begin
        decipher_0_iibox_ce186 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce187 = 1'b1;
    end else begin
        decipher_0_iibox_ce187 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce188 = 1'b1;
    end else begin
        decipher_0_iibox_ce188 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce189 = 1'b1;
    end else begin
        decipher_0_iibox_ce189 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce19 = 1'b1;
    end else begin
        decipher_0_iibox_ce19 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce190 = 1'b1;
    end else begin
        decipher_0_iibox_ce190 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce191 = 1'b1;
    end else begin
        decipher_0_iibox_ce191 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce2 = 1'b1;
    end else begin
        decipher_0_iibox_ce2 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce20 = 1'b1;
    end else begin
        decipher_0_iibox_ce20 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce21 = 1'b1;
    end else begin
        decipher_0_iibox_ce21 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce22 = 1'b1;
    end else begin
        decipher_0_iibox_ce22 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce23 = 1'b1;
    end else begin
        decipher_0_iibox_ce23 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce24 = 1'b1;
    end else begin
        decipher_0_iibox_ce24 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce25 = 1'b1;
    end else begin
        decipher_0_iibox_ce25 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce26 = 1'b1;
    end else begin
        decipher_0_iibox_ce26 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce27 = 1'b1;
    end else begin
        decipher_0_iibox_ce27 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce28 = 1'b1;
    end else begin
        decipher_0_iibox_ce28 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce29 = 1'b1;
    end else begin
        decipher_0_iibox_ce29 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce3 = 1'b1;
    end else begin
        decipher_0_iibox_ce3 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce30 = 1'b1;
    end else begin
        decipher_0_iibox_ce30 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce31 = 1'b1;
    end else begin
        decipher_0_iibox_ce31 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce32 = 1'b1;
    end else begin
        decipher_0_iibox_ce32 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce33 = 1'b1;
    end else begin
        decipher_0_iibox_ce33 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce34 = 1'b1;
    end else begin
        decipher_0_iibox_ce34 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce35 = 1'b1;
    end else begin
        decipher_0_iibox_ce35 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce36 = 1'b1;
    end else begin
        decipher_0_iibox_ce36 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce37 = 1'b1;
    end else begin
        decipher_0_iibox_ce37 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce38 = 1'b1;
    end else begin
        decipher_0_iibox_ce38 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce39 = 1'b1;
    end else begin
        decipher_0_iibox_ce39 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce4 = 1'b1;
    end else begin
        decipher_0_iibox_ce4 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce40 = 1'b1;
    end else begin
        decipher_0_iibox_ce40 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce41 = 1'b1;
    end else begin
        decipher_0_iibox_ce41 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce42 = 1'b1;
    end else begin
        decipher_0_iibox_ce42 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce43 = 1'b1;
    end else begin
        decipher_0_iibox_ce43 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce44 = 1'b1;
    end else begin
        decipher_0_iibox_ce44 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce45 = 1'b1;
    end else begin
        decipher_0_iibox_ce45 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce46 = 1'b1;
    end else begin
        decipher_0_iibox_ce46 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce47 = 1'b1;
    end else begin
        decipher_0_iibox_ce47 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce48 = 1'b1;
    end else begin
        decipher_0_iibox_ce48 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce49 = 1'b1;
    end else begin
        decipher_0_iibox_ce49 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce5 = 1'b1;
    end else begin
        decipher_0_iibox_ce5 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce50 = 1'b1;
    end else begin
        decipher_0_iibox_ce50 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce51 = 1'b1;
    end else begin
        decipher_0_iibox_ce51 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce52 = 1'b1;
    end else begin
        decipher_0_iibox_ce52 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce53 = 1'b1;
    end else begin
        decipher_0_iibox_ce53 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce54 = 1'b1;
    end else begin
        decipher_0_iibox_ce54 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce55 = 1'b1;
    end else begin
        decipher_0_iibox_ce55 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce56 = 1'b1;
    end else begin
        decipher_0_iibox_ce56 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce57 = 1'b1;
    end else begin
        decipher_0_iibox_ce57 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce58 = 1'b1;
    end else begin
        decipher_0_iibox_ce58 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce59 = 1'b1;
    end else begin
        decipher_0_iibox_ce59 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce6 = 1'b1;
    end else begin
        decipher_0_iibox_ce6 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce60 = 1'b1;
    end else begin
        decipher_0_iibox_ce60 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce61 = 1'b1;
    end else begin
        decipher_0_iibox_ce61 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce62 = 1'b1;
    end else begin
        decipher_0_iibox_ce62 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce63 = 1'b1;
    end else begin
        decipher_0_iibox_ce63 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce64 = 1'b1;
    end else begin
        decipher_0_iibox_ce64 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce65 = 1'b1;
    end else begin
        decipher_0_iibox_ce65 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce66 = 1'b1;
    end else begin
        decipher_0_iibox_ce66 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce67 = 1'b1;
    end else begin
        decipher_0_iibox_ce67 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce68 = 1'b1;
    end else begin
        decipher_0_iibox_ce68 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce69 = 1'b1;
    end else begin
        decipher_0_iibox_ce69 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce7 = 1'b1;
    end else begin
        decipher_0_iibox_ce7 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce70 = 1'b1;
    end else begin
        decipher_0_iibox_ce70 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce71 = 1'b1;
    end else begin
        decipher_0_iibox_ce71 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce72 = 1'b1;
    end else begin
        decipher_0_iibox_ce72 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce73 = 1'b1;
    end else begin
        decipher_0_iibox_ce73 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce74 = 1'b1;
    end else begin
        decipher_0_iibox_ce74 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce75 = 1'b1;
    end else begin
        decipher_0_iibox_ce75 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce76 = 1'b1;
    end else begin
        decipher_0_iibox_ce76 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce77 = 1'b1;
    end else begin
        decipher_0_iibox_ce77 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce78 = 1'b1;
    end else begin
        decipher_0_iibox_ce78 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce79 = 1'b1;
    end else begin
        decipher_0_iibox_ce79 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce8 = 1'b1;
    end else begin
        decipher_0_iibox_ce8 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce80 = 1'b1;
    end else begin
        decipher_0_iibox_ce80 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce81 = 1'b1;
    end else begin
        decipher_0_iibox_ce81 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce82 = 1'b1;
    end else begin
        decipher_0_iibox_ce82 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce83 = 1'b1;
    end else begin
        decipher_0_iibox_ce83 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce84 = 1'b1;
    end else begin
        decipher_0_iibox_ce84 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce85 = 1'b1;
    end else begin
        decipher_0_iibox_ce85 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce86 = 1'b1;
    end else begin
        decipher_0_iibox_ce86 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce87 = 1'b1;
    end else begin
        decipher_0_iibox_ce87 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce88 = 1'b1;
    end else begin
        decipher_0_iibox_ce88 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce89 = 1'b1;
    end else begin
        decipher_0_iibox_ce89 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce9 = 1'b1;
    end else begin
        decipher_0_iibox_ce9 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce90 = 1'b1;
    end else begin
        decipher_0_iibox_ce90 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce91 = 1'b1;
    end else begin
        decipher_0_iibox_ce91 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce92 = 1'b1;
    end else begin
        decipher_0_iibox_ce92 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce93 = 1'b1;
    end else begin
        decipher_0_iibox_ce93 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce94 = 1'b1;
    end else begin
        decipher_0_iibox_ce94 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce95 = 1'b1;
    end else begin
        decipher_0_iibox_ce95 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce96 = 1'b1;
    end else begin
        decipher_0_iibox_ce96 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce97 = 1'b1;
    end else begin
        decipher_0_iibox_ce97 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce98 = 1'b1;
    end else begin
        decipher_0_iibox_ce98 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce99 = 1'b1;
    end else begin
        decipher_0_iibox_ce99 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_state10_pp0_stage0_iter9 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage0_iter10 = ~(1'b1 == 1'b1);

assign ap_block_state12_pp0_stage0_iter11 = ~(1'b1 == 1'b1);

assign ap_block_state13_pp0_stage0_iter12 = ~(1'b1 == 1'b1);

assign ap_block_state14_pp0_stage0_iter13 = ~(1'b1 == 1'b1);

assign ap_block_state15_pp0_stage0_iter14 = ~(1'b1 == 1'b1);

assign ap_block_state16_pp0_stage0_iter15 = ~(1'b1 == 1'b1);

assign ap_block_state17_pp0_stage0_iter16 = ~(1'b1 == 1'b1);

assign ap_block_state18_pp0_stage0_iter17 = ~(1'b1 == 1'b1);

assign ap_block_state19_pp0_stage0_iter18 = ~(1'b1 == 1'b1);

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state20_pp0_stage0_iter19 = ~(1'b1 == 1'b1);

assign ap_block_state21_pp0_stage0_iter20 = ~(1'b1 == 1'b1);

assign ap_block_state22_pp0_stage0_iter21 = ~(1'b1 == 1'b1);

assign ap_block_state23_pp0_stage0_iter22 = ~(1'b1 == 1'b1);

assign ap_block_state24_pp0_stage0_iter23 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter8 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_enable_reg_pp0_iter0 = ap_start;

assign ap_return = (p_read13_reg_18005_pp0_iter22_reg ^ p_Result_35_fu_17909_p17);

assign decipher_0_i32box_address0 = zext_ln708_354_fu_16992_p1;

assign decipher_0_i32box_address1 = zext_ln708_353_fu_16977_p1;

assign decipher_0_i32box_address10 = zext_ln708_344_fu_16842_p1;

assign decipher_0_i32box_address100 = zext_ln708_158_fu_9810_p1;

assign decipher_0_i32box_address101 = zext_ln708_157_fu_9795_p1;

assign decipher_0_i32box_address102 = zext_ln708_156_fu_9780_p1;

assign decipher_0_i32box_address103 = zext_ln708_155_fu_9765_p1;

assign decipher_0_i32box_address104 = zext_ln708_154_fu_9750_p1;

assign decipher_0_i32box_address105 = zext_ln708_153_fu_9735_p1;

assign decipher_0_i32box_address106 = zext_ln708_152_fu_9720_p1;

assign decipher_0_i32box_address107 = zext_ln708_151_fu_9705_p1;

assign decipher_0_i32box_address108 = zext_ln708_150_fu_9690_p1;

assign decipher_0_i32box_address109 = zext_ln708_149_fu_9675_p1;

assign decipher_0_i32box_address11 = zext_ln708_343_fu_16827_p1;

assign decipher_0_i32box_address110 = zext_ln708_148_fu_9660_p1;

assign decipher_0_i32box_address111 = zext_ln708_147_fu_9645_p1;

assign decipher_0_i32box_address112 = zext_ln708_130_fu_8683_p1;

assign decipher_0_i32box_address113 = zext_ln708_129_fu_8668_p1;

assign decipher_0_i32box_address114 = zext_ln708_128_fu_8653_p1;

assign decipher_0_i32box_address115 = zext_ln708_127_fu_8638_p1;

assign decipher_0_i32box_address116 = zext_ln708_126_fu_8623_p1;

assign decipher_0_i32box_address117 = zext_ln708_125_fu_8608_p1;

assign decipher_0_i32box_address118 = zext_ln708_124_fu_8593_p1;

assign decipher_0_i32box_address119 = zext_ln708_123_fu_8578_p1;

assign decipher_0_i32box_address12 = zext_ln708_342_fu_16812_p1;

assign decipher_0_i32box_address120 = zext_ln708_122_fu_8563_p1;

assign decipher_0_i32box_address121 = zext_ln708_121_fu_8548_p1;

assign decipher_0_i32box_address122 = zext_ln708_120_fu_8533_p1;

assign decipher_0_i32box_address123 = zext_ln708_119_fu_8518_p1;

assign decipher_0_i32box_address124 = zext_ln708_118_fu_8503_p1;

assign decipher_0_i32box_address125 = zext_ln708_117_fu_8488_p1;

assign decipher_0_i32box_address126 = zext_ln708_116_fu_8473_p1;

assign decipher_0_i32box_address127 = zext_ln708_115_fu_8458_p1;

assign decipher_0_i32box_address128 = zext_ln708_98_fu_7496_p1;

assign decipher_0_i32box_address129 = zext_ln708_97_fu_7481_p1;

assign decipher_0_i32box_address13 = zext_ln708_341_fu_16797_p1;

assign decipher_0_i32box_address130 = zext_ln708_96_fu_7466_p1;

assign decipher_0_i32box_address131 = zext_ln708_95_fu_7451_p1;

assign decipher_0_i32box_address132 = zext_ln708_94_fu_7436_p1;

assign decipher_0_i32box_address133 = zext_ln708_93_fu_7421_p1;

assign decipher_0_i32box_address134 = zext_ln708_92_fu_7406_p1;

assign decipher_0_i32box_address135 = zext_ln708_91_fu_7391_p1;

assign decipher_0_i32box_address136 = zext_ln708_90_fu_7376_p1;

assign decipher_0_i32box_address137 = zext_ln708_89_fu_7361_p1;

assign decipher_0_i32box_address138 = zext_ln708_88_fu_7346_p1;

assign decipher_0_i32box_address139 = zext_ln708_87_fu_7331_p1;

assign decipher_0_i32box_address14 = zext_ln708_340_fu_16782_p1;

assign decipher_0_i32box_address140 = zext_ln708_86_fu_7316_p1;

assign decipher_0_i32box_address141 = zext_ln708_85_fu_7301_p1;

assign decipher_0_i32box_address142 = zext_ln708_84_fu_7286_p1;

assign decipher_0_i32box_address143 = zext_ln708_83_fu_7271_p1;

assign decipher_0_i32box_address144 = zext_ln708_66_fu_6309_p1;

assign decipher_0_i32box_address145 = zext_ln708_65_fu_6294_p1;

assign decipher_0_i32box_address146 = zext_ln708_64_fu_6279_p1;

assign decipher_0_i32box_address147 = zext_ln708_63_fu_6264_p1;

assign decipher_0_i32box_address148 = zext_ln708_62_fu_6249_p1;

assign decipher_0_i32box_address149 = zext_ln708_61_fu_6234_p1;

assign decipher_0_i32box_address15 = zext_ln708_339_fu_16767_p1;

assign decipher_0_i32box_address150 = zext_ln708_60_fu_6219_p1;

assign decipher_0_i32box_address151 = zext_ln708_59_fu_6204_p1;

assign decipher_0_i32box_address152 = zext_ln708_58_fu_6189_p1;

assign decipher_0_i32box_address153 = zext_ln708_57_fu_6174_p1;

assign decipher_0_i32box_address154 = zext_ln708_56_fu_6159_p1;

assign decipher_0_i32box_address155 = zext_ln708_55_fu_6144_p1;

assign decipher_0_i32box_address156 = zext_ln708_54_fu_6129_p1;

assign decipher_0_i32box_address157 = zext_ln708_53_fu_6114_p1;

assign decipher_0_i32box_address158 = zext_ln708_52_fu_6099_p1;

assign decipher_0_i32box_address159 = zext_ln708_51_fu_6084_p1;

assign decipher_0_i32box_address16 = zext_ln708_322_fu_15805_p1;

assign decipher_0_i32box_address160 = zext_ln708_34_fu_5122_p1;

assign decipher_0_i32box_address161 = zext_ln708_33_fu_5107_p1;

assign decipher_0_i32box_address162 = zext_ln708_32_fu_5092_p1;

assign decipher_0_i32box_address163 = zext_ln708_31_fu_5077_p1;

assign decipher_0_i32box_address164 = zext_ln708_30_fu_5062_p1;

assign decipher_0_i32box_address165 = zext_ln708_29_fu_5047_p1;

assign decipher_0_i32box_address166 = zext_ln708_28_fu_5032_p1;

assign decipher_0_i32box_address167 = zext_ln708_27_fu_5017_p1;

assign decipher_0_i32box_address168 = zext_ln708_26_fu_5002_p1;

assign decipher_0_i32box_address169 = zext_ln708_25_fu_4987_p1;

assign decipher_0_i32box_address17 = zext_ln708_321_fu_15790_p1;

assign decipher_0_i32box_address170 = zext_ln708_24_fu_4972_p1;

assign decipher_0_i32box_address171 = zext_ln708_23_fu_4957_p1;

assign decipher_0_i32box_address172 = zext_ln708_22_fu_4942_p1;

assign decipher_0_i32box_address173 = zext_ln708_21_fu_4927_p1;

assign decipher_0_i32box_address174 = zext_ln708_20_fu_4912_p1;

assign decipher_0_i32box_address175 = zext_ln708_19_fu_4897_p1;

assign decipher_0_i32box_address18 = zext_ln708_320_fu_15775_p1;

assign decipher_0_i32box_address19 = zext_ln708_319_fu_15760_p1;

assign decipher_0_i32box_address2 = zext_ln708_352_fu_16962_p1;

assign decipher_0_i32box_address20 = zext_ln708_318_fu_15745_p1;

assign decipher_0_i32box_address21 = zext_ln708_317_fu_15730_p1;

assign decipher_0_i32box_address22 = zext_ln708_316_fu_15715_p1;

assign decipher_0_i32box_address23 = zext_ln708_315_fu_15700_p1;

assign decipher_0_i32box_address24 = zext_ln708_314_fu_15685_p1;

assign decipher_0_i32box_address25 = zext_ln708_313_fu_15670_p1;

assign decipher_0_i32box_address26 = zext_ln708_312_fu_15655_p1;

assign decipher_0_i32box_address27 = zext_ln708_311_fu_15640_p1;

assign decipher_0_i32box_address28 = zext_ln708_310_fu_15625_p1;

assign decipher_0_i32box_address29 = zext_ln708_309_fu_15610_p1;

assign decipher_0_i32box_address3 = zext_ln708_351_fu_16947_p1;

assign decipher_0_i32box_address30 = zext_ln708_308_fu_15595_p1;

assign decipher_0_i32box_address31 = zext_ln708_307_fu_15580_p1;

assign decipher_0_i32box_address32 = zext_ln708_290_fu_14618_p1;

assign decipher_0_i32box_address33 = zext_ln708_289_fu_14603_p1;

assign decipher_0_i32box_address34 = zext_ln708_288_fu_14588_p1;

assign decipher_0_i32box_address35 = zext_ln708_287_fu_14573_p1;

assign decipher_0_i32box_address36 = zext_ln708_286_fu_14558_p1;

assign decipher_0_i32box_address37 = zext_ln708_285_fu_14543_p1;

assign decipher_0_i32box_address38 = zext_ln708_284_fu_14528_p1;

assign decipher_0_i32box_address39 = zext_ln708_283_fu_14513_p1;

assign decipher_0_i32box_address4 = zext_ln708_350_fu_16932_p1;

assign decipher_0_i32box_address40 = zext_ln708_282_fu_14498_p1;

assign decipher_0_i32box_address41 = zext_ln708_281_fu_14483_p1;

assign decipher_0_i32box_address42 = zext_ln708_280_fu_14468_p1;

assign decipher_0_i32box_address43 = zext_ln708_279_fu_14453_p1;

assign decipher_0_i32box_address44 = zext_ln708_278_fu_14438_p1;

assign decipher_0_i32box_address45 = zext_ln708_277_fu_14423_p1;

assign decipher_0_i32box_address46 = zext_ln708_276_fu_14408_p1;

assign decipher_0_i32box_address47 = zext_ln708_275_fu_14393_p1;

assign decipher_0_i32box_address48 = zext_ln708_258_fu_13431_p1;

assign decipher_0_i32box_address49 = zext_ln708_257_fu_13416_p1;

assign decipher_0_i32box_address5 = zext_ln708_349_fu_16917_p1;

assign decipher_0_i32box_address50 = zext_ln708_256_fu_13401_p1;

assign decipher_0_i32box_address51 = zext_ln708_255_fu_13386_p1;

assign decipher_0_i32box_address52 = zext_ln708_254_fu_13371_p1;

assign decipher_0_i32box_address53 = zext_ln708_253_fu_13356_p1;

assign decipher_0_i32box_address54 = zext_ln708_252_fu_13341_p1;

assign decipher_0_i32box_address55 = zext_ln708_251_fu_13326_p1;

assign decipher_0_i32box_address56 = zext_ln708_250_fu_13311_p1;

assign decipher_0_i32box_address57 = zext_ln708_249_fu_13296_p1;

assign decipher_0_i32box_address58 = zext_ln708_248_fu_13281_p1;

assign decipher_0_i32box_address59 = zext_ln708_247_fu_13266_p1;

assign decipher_0_i32box_address6 = zext_ln708_348_fu_16902_p1;

assign decipher_0_i32box_address60 = zext_ln708_246_fu_13251_p1;

assign decipher_0_i32box_address61 = zext_ln708_245_fu_13236_p1;

assign decipher_0_i32box_address62 = zext_ln708_244_fu_13221_p1;

assign decipher_0_i32box_address63 = zext_ln708_243_fu_13206_p1;

assign decipher_0_i32box_address64 = zext_ln708_226_fu_12244_p1;

assign decipher_0_i32box_address65 = zext_ln708_225_fu_12229_p1;

assign decipher_0_i32box_address66 = zext_ln708_224_fu_12214_p1;

assign decipher_0_i32box_address67 = zext_ln708_223_fu_12199_p1;

assign decipher_0_i32box_address68 = zext_ln708_222_fu_12184_p1;

assign decipher_0_i32box_address69 = zext_ln708_221_fu_12169_p1;

assign decipher_0_i32box_address7 = zext_ln708_347_fu_16887_p1;

assign decipher_0_i32box_address70 = zext_ln708_220_fu_12154_p1;

assign decipher_0_i32box_address71 = zext_ln708_219_fu_12139_p1;

assign decipher_0_i32box_address72 = zext_ln708_218_fu_12124_p1;

assign decipher_0_i32box_address73 = zext_ln708_217_fu_12109_p1;

assign decipher_0_i32box_address74 = zext_ln708_216_fu_12094_p1;

assign decipher_0_i32box_address75 = zext_ln708_215_fu_12079_p1;

assign decipher_0_i32box_address76 = zext_ln708_214_fu_12064_p1;

assign decipher_0_i32box_address77 = zext_ln708_213_fu_12049_p1;

assign decipher_0_i32box_address78 = zext_ln708_212_fu_12034_p1;

assign decipher_0_i32box_address79 = zext_ln708_211_fu_12019_p1;

assign decipher_0_i32box_address8 = zext_ln708_346_fu_16872_p1;

assign decipher_0_i32box_address80 = zext_ln708_194_fu_11057_p1;

assign decipher_0_i32box_address81 = zext_ln708_193_fu_11042_p1;

assign decipher_0_i32box_address82 = zext_ln708_192_fu_11027_p1;

assign decipher_0_i32box_address83 = zext_ln708_191_fu_11012_p1;

assign decipher_0_i32box_address84 = zext_ln708_190_fu_10997_p1;

assign decipher_0_i32box_address85 = zext_ln708_189_fu_10982_p1;

assign decipher_0_i32box_address86 = zext_ln708_188_fu_10967_p1;

assign decipher_0_i32box_address87 = zext_ln708_187_fu_10952_p1;

assign decipher_0_i32box_address88 = zext_ln708_186_fu_10937_p1;

assign decipher_0_i32box_address89 = zext_ln708_185_fu_10922_p1;

assign decipher_0_i32box_address9 = zext_ln708_345_fu_16857_p1;

assign decipher_0_i32box_address90 = zext_ln708_184_fu_10907_p1;

assign decipher_0_i32box_address91 = zext_ln708_183_fu_10892_p1;

assign decipher_0_i32box_address92 = zext_ln708_182_fu_10877_p1;

assign decipher_0_i32box_address93 = zext_ln708_181_fu_10862_p1;

assign decipher_0_i32box_address94 = zext_ln708_180_fu_10847_p1;

assign decipher_0_i32box_address95 = zext_ln708_179_fu_10832_p1;

assign decipher_0_i32box_address96 = zext_ln708_162_fu_9870_p1;

assign decipher_0_i32box_address97 = zext_ln708_161_fu_9855_p1;

assign decipher_0_i32box_address98 = zext_ln708_160_fu_9840_p1;

assign decipher_0_i32box_address99 = zext_ln708_159_fu_9825_p1;

assign decipher_0_iibox_address0 = zext_ln708_370_fu_17904_p1;

assign decipher_0_iibox_address1 = zext_ln708_369_fu_17899_p1;

assign decipher_0_iibox_address10 = zext_ln708_360_fu_17854_p1;

assign decipher_0_iibox_address100 = zext_ln708_174_fu_10762_p1;

assign decipher_0_iibox_address101 = zext_ln708_173_fu_10757_p1;

assign decipher_0_iibox_address102 = zext_ln708_172_fu_10752_p1;

assign decipher_0_iibox_address103 = zext_ln708_171_fu_10747_p1;

assign decipher_0_iibox_address104 = zext_ln708_170_fu_10742_p1;

assign decipher_0_iibox_address105 = zext_ln708_169_fu_10737_p1;

assign decipher_0_iibox_address106 = zext_ln708_168_fu_10732_p1;

assign decipher_0_iibox_address107 = zext_ln708_167_fu_10727_p1;

assign decipher_0_iibox_address108 = zext_ln708_166_fu_10722_p1;

assign decipher_0_iibox_address109 = zext_ln708_165_fu_10717_p1;

assign decipher_0_iibox_address11 = zext_ln708_359_fu_17849_p1;

assign decipher_0_iibox_address110 = zext_ln708_164_fu_10712_p1;

assign decipher_0_iibox_address111 = zext_ln708_163_fu_10707_p1;

assign decipher_0_iibox_address112 = zext_ln708_146_fu_9595_p1;

assign decipher_0_iibox_address113 = zext_ln708_145_fu_9590_p1;

assign decipher_0_iibox_address114 = zext_ln708_144_fu_9585_p1;

assign decipher_0_iibox_address115 = zext_ln708_143_fu_9580_p1;

assign decipher_0_iibox_address116 = zext_ln708_142_fu_9575_p1;

assign decipher_0_iibox_address117 = zext_ln708_141_fu_9570_p1;

assign decipher_0_iibox_address118 = zext_ln708_140_fu_9565_p1;

assign decipher_0_iibox_address119 = zext_ln708_139_fu_9560_p1;

assign decipher_0_iibox_address12 = zext_ln708_358_fu_17844_p1;

assign decipher_0_iibox_address120 = zext_ln708_138_fu_9555_p1;

assign decipher_0_iibox_address121 = zext_ln708_137_fu_9550_p1;

assign decipher_0_iibox_address122 = zext_ln708_136_fu_9545_p1;

assign decipher_0_iibox_address123 = zext_ln708_135_fu_9540_p1;

assign decipher_0_iibox_address124 = zext_ln708_134_fu_9535_p1;

assign decipher_0_iibox_address125 = zext_ln708_133_fu_9530_p1;

assign decipher_0_iibox_address126 = zext_ln708_132_fu_9525_p1;

assign decipher_0_iibox_address127 = zext_ln708_131_fu_9520_p1;

assign decipher_0_iibox_address128 = zext_ln708_114_fu_8408_p1;

assign decipher_0_iibox_address129 = zext_ln708_113_fu_8403_p1;

assign decipher_0_iibox_address13 = zext_ln708_357_fu_17839_p1;

assign decipher_0_iibox_address130 = zext_ln708_112_fu_8398_p1;

assign decipher_0_iibox_address131 = zext_ln708_111_fu_8393_p1;

assign decipher_0_iibox_address132 = zext_ln708_110_fu_8388_p1;

assign decipher_0_iibox_address133 = zext_ln708_109_fu_8383_p1;

assign decipher_0_iibox_address134 = zext_ln708_108_fu_8378_p1;

assign decipher_0_iibox_address135 = zext_ln708_107_fu_8373_p1;

assign decipher_0_iibox_address136 = zext_ln708_106_fu_8368_p1;

assign decipher_0_iibox_address137 = zext_ln708_105_fu_8363_p1;

assign decipher_0_iibox_address138 = zext_ln708_104_fu_8358_p1;

assign decipher_0_iibox_address139 = zext_ln708_103_fu_8353_p1;

assign decipher_0_iibox_address14 = zext_ln708_356_fu_17834_p1;

assign decipher_0_iibox_address140 = zext_ln708_102_fu_8348_p1;

assign decipher_0_iibox_address141 = zext_ln708_101_fu_8343_p1;

assign decipher_0_iibox_address142 = zext_ln708_100_fu_8338_p1;

assign decipher_0_iibox_address143 = zext_ln708_99_fu_8333_p1;

assign decipher_0_iibox_address144 = zext_ln708_82_fu_7221_p1;

assign decipher_0_iibox_address145 = zext_ln708_81_fu_7216_p1;

assign decipher_0_iibox_address146 = zext_ln708_80_fu_7211_p1;

assign decipher_0_iibox_address147 = zext_ln708_79_fu_7206_p1;

assign decipher_0_iibox_address148 = zext_ln708_78_fu_7201_p1;

assign decipher_0_iibox_address149 = zext_ln708_77_fu_7196_p1;

assign decipher_0_iibox_address15 = zext_ln708_355_fu_17829_p1;

assign decipher_0_iibox_address150 = zext_ln708_76_fu_7191_p1;

assign decipher_0_iibox_address151 = zext_ln708_75_fu_7186_p1;

assign decipher_0_iibox_address152 = zext_ln708_74_fu_7181_p1;

assign decipher_0_iibox_address153 = zext_ln708_73_fu_7176_p1;

assign decipher_0_iibox_address154 = zext_ln708_72_fu_7171_p1;

assign decipher_0_iibox_address155 = zext_ln708_71_fu_7166_p1;

assign decipher_0_iibox_address156 = zext_ln708_70_fu_7161_p1;

assign decipher_0_iibox_address157 = zext_ln708_69_fu_7156_p1;

assign decipher_0_iibox_address158 = zext_ln708_68_fu_7151_p1;

assign decipher_0_iibox_address159 = zext_ln708_67_fu_7146_p1;

assign decipher_0_iibox_address16 = zext_ln708_338_fu_16717_p1;

assign decipher_0_iibox_address160 = zext_ln708_50_fu_6034_p1;

assign decipher_0_iibox_address161 = zext_ln708_49_fu_6029_p1;

assign decipher_0_iibox_address162 = zext_ln708_48_fu_6024_p1;

assign decipher_0_iibox_address163 = zext_ln708_47_fu_6019_p1;

assign decipher_0_iibox_address164 = zext_ln708_46_fu_6014_p1;

assign decipher_0_iibox_address165 = zext_ln708_45_fu_6009_p1;

assign decipher_0_iibox_address166 = zext_ln708_44_fu_6004_p1;

assign decipher_0_iibox_address167 = zext_ln708_43_fu_5999_p1;

assign decipher_0_iibox_address168 = zext_ln708_42_fu_5994_p1;

assign decipher_0_iibox_address169 = zext_ln708_41_fu_5989_p1;

assign decipher_0_iibox_address17 = zext_ln708_337_fu_16712_p1;

assign decipher_0_iibox_address170 = zext_ln708_40_fu_5984_p1;

assign decipher_0_iibox_address171 = zext_ln708_39_fu_5979_p1;

assign decipher_0_iibox_address172 = zext_ln708_38_fu_5974_p1;

assign decipher_0_iibox_address173 = zext_ln708_37_fu_5969_p1;

assign decipher_0_iibox_address174 = zext_ln708_36_fu_5964_p1;

assign decipher_0_iibox_address175 = zext_ln708_35_fu_5959_p1;

assign decipher_0_iibox_address176 = zext_ln708_18_fu_4847_p1;

assign decipher_0_iibox_address177 = zext_ln708_17_fu_4832_p1;

assign decipher_0_iibox_address178 = zext_ln708_16_fu_4817_p1;

assign decipher_0_iibox_address179 = zext_ln708_15_fu_4802_p1;

assign decipher_0_iibox_address18 = zext_ln708_336_fu_16707_p1;

assign decipher_0_iibox_address180 = zext_ln708_14_fu_4787_p1;

assign decipher_0_iibox_address181 = zext_ln708_13_fu_4772_p1;

assign decipher_0_iibox_address182 = zext_ln708_12_fu_4757_p1;

assign decipher_0_iibox_address183 = zext_ln708_11_fu_4742_p1;

assign decipher_0_iibox_address184 = zext_ln708_10_fu_4727_p1;

assign decipher_0_iibox_address185 = zext_ln708_9_fu_4712_p1;

assign decipher_0_iibox_address186 = zext_ln708_8_fu_4697_p1;

assign decipher_0_iibox_address187 = zext_ln708_7_fu_4682_p1;

assign decipher_0_iibox_address188 = zext_ln708_6_fu_4667_p1;

assign decipher_0_iibox_address189 = zext_ln708_5_fu_4652_p1;

assign decipher_0_iibox_address19 = zext_ln708_335_fu_16702_p1;

assign decipher_0_iibox_address190 = zext_ln708_4_fu_4637_p1;

assign decipher_0_iibox_address191 = zext_ln708_fu_4622_p1;

assign decipher_0_iibox_address2 = zext_ln708_368_fu_17894_p1;

assign decipher_0_iibox_address20 = zext_ln708_334_fu_16697_p1;

assign decipher_0_iibox_address21 = zext_ln708_333_fu_16692_p1;

assign decipher_0_iibox_address22 = zext_ln708_332_fu_16687_p1;

assign decipher_0_iibox_address23 = zext_ln708_331_fu_16682_p1;

assign decipher_0_iibox_address24 = zext_ln708_330_fu_16677_p1;

assign decipher_0_iibox_address25 = zext_ln708_329_fu_16672_p1;

assign decipher_0_iibox_address26 = zext_ln708_328_fu_16667_p1;

assign decipher_0_iibox_address27 = zext_ln708_327_fu_16662_p1;

assign decipher_0_iibox_address28 = zext_ln708_326_fu_16657_p1;

assign decipher_0_iibox_address29 = zext_ln708_325_fu_16652_p1;

assign decipher_0_iibox_address3 = zext_ln708_367_fu_17889_p1;

assign decipher_0_iibox_address30 = zext_ln708_324_fu_16647_p1;

assign decipher_0_iibox_address31 = zext_ln708_323_fu_16642_p1;

assign decipher_0_iibox_address32 = zext_ln708_306_fu_15530_p1;

assign decipher_0_iibox_address33 = zext_ln708_305_fu_15525_p1;

assign decipher_0_iibox_address34 = zext_ln708_304_fu_15520_p1;

assign decipher_0_iibox_address35 = zext_ln708_303_fu_15515_p1;

assign decipher_0_iibox_address36 = zext_ln708_302_fu_15510_p1;

assign decipher_0_iibox_address37 = zext_ln708_301_fu_15505_p1;

assign decipher_0_iibox_address38 = zext_ln708_300_fu_15500_p1;

assign decipher_0_iibox_address39 = zext_ln708_299_fu_15495_p1;

assign decipher_0_iibox_address4 = zext_ln708_366_fu_17884_p1;

assign decipher_0_iibox_address40 = zext_ln708_298_fu_15490_p1;

assign decipher_0_iibox_address41 = zext_ln708_297_fu_15485_p1;

assign decipher_0_iibox_address42 = zext_ln708_296_fu_15480_p1;

assign decipher_0_iibox_address43 = zext_ln708_295_fu_15475_p1;

assign decipher_0_iibox_address44 = zext_ln708_294_fu_15470_p1;

assign decipher_0_iibox_address45 = zext_ln708_293_fu_15465_p1;

assign decipher_0_iibox_address46 = zext_ln708_292_fu_15460_p1;

assign decipher_0_iibox_address47 = zext_ln708_291_fu_15455_p1;

assign decipher_0_iibox_address48 = zext_ln708_274_fu_14343_p1;

assign decipher_0_iibox_address49 = zext_ln708_273_fu_14338_p1;

assign decipher_0_iibox_address5 = zext_ln708_365_fu_17879_p1;

assign decipher_0_iibox_address50 = zext_ln708_272_fu_14333_p1;

assign decipher_0_iibox_address51 = zext_ln708_271_fu_14328_p1;

assign decipher_0_iibox_address52 = zext_ln708_270_fu_14323_p1;

assign decipher_0_iibox_address53 = zext_ln708_269_fu_14318_p1;

assign decipher_0_iibox_address54 = zext_ln708_268_fu_14313_p1;

assign decipher_0_iibox_address55 = zext_ln708_267_fu_14308_p1;

assign decipher_0_iibox_address56 = zext_ln708_266_fu_14303_p1;

assign decipher_0_iibox_address57 = zext_ln708_265_fu_14298_p1;

assign decipher_0_iibox_address58 = zext_ln708_264_fu_14293_p1;

assign decipher_0_iibox_address59 = zext_ln708_263_fu_14288_p1;

assign decipher_0_iibox_address6 = zext_ln708_364_fu_17874_p1;

assign decipher_0_iibox_address60 = zext_ln708_262_fu_14283_p1;

assign decipher_0_iibox_address61 = zext_ln708_261_fu_14278_p1;

assign decipher_0_iibox_address62 = zext_ln708_260_fu_14273_p1;

assign decipher_0_iibox_address63 = zext_ln708_259_fu_14268_p1;

assign decipher_0_iibox_address64 = zext_ln708_242_fu_13156_p1;

assign decipher_0_iibox_address65 = zext_ln708_241_fu_13151_p1;

assign decipher_0_iibox_address66 = zext_ln708_240_fu_13146_p1;

assign decipher_0_iibox_address67 = zext_ln708_239_fu_13141_p1;

assign decipher_0_iibox_address68 = zext_ln708_238_fu_13136_p1;

assign decipher_0_iibox_address69 = zext_ln708_237_fu_13131_p1;

assign decipher_0_iibox_address7 = zext_ln708_363_fu_17869_p1;

assign decipher_0_iibox_address70 = zext_ln708_236_fu_13126_p1;

assign decipher_0_iibox_address71 = zext_ln708_235_fu_13121_p1;

assign decipher_0_iibox_address72 = zext_ln708_234_fu_13116_p1;

assign decipher_0_iibox_address73 = zext_ln708_233_fu_13111_p1;

assign decipher_0_iibox_address74 = zext_ln708_232_fu_13106_p1;

assign decipher_0_iibox_address75 = zext_ln708_231_fu_13101_p1;

assign decipher_0_iibox_address76 = zext_ln708_230_fu_13096_p1;

assign decipher_0_iibox_address77 = zext_ln708_229_fu_13091_p1;

assign decipher_0_iibox_address78 = zext_ln708_228_fu_13086_p1;

assign decipher_0_iibox_address79 = zext_ln708_227_fu_13081_p1;

assign decipher_0_iibox_address8 = zext_ln708_362_fu_17864_p1;

assign decipher_0_iibox_address80 = zext_ln708_210_fu_11969_p1;

assign decipher_0_iibox_address81 = zext_ln708_209_fu_11964_p1;

assign decipher_0_iibox_address82 = zext_ln708_208_fu_11959_p1;

assign decipher_0_iibox_address83 = zext_ln708_207_fu_11954_p1;

assign decipher_0_iibox_address84 = zext_ln708_206_fu_11949_p1;

assign decipher_0_iibox_address85 = zext_ln708_205_fu_11944_p1;

assign decipher_0_iibox_address86 = zext_ln708_204_fu_11939_p1;

assign decipher_0_iibox_address87 = zext_ln708_203_fu_11934_p1;

assign decipher_0_iibox_address88 = zext_ln708_202_fu_11929_p1;

assign decipher_0_iibox_address89 = zext_ln708_201_fu_11924_p1;

assign decipher_0_iibox_address9 = zext_ln708_361_fu_17859_p1;

assign decipher_0_iibox_address90 = zext_ln708_200_fu_11919_p1;

assign decipher_0_iibox_address91 = zext_ln708_199_fu_11914_p1;

assign decipher_0_iibox_address92 = zext_ln708_198_fu_11909_p1;

assign decipher_0_iibox_address93 = zext_ln708_197_fu_11904_p1;

assign decipher_0_iibox_address94 = zext_ln708_196_fu_11899_p1;

assign decipher_0_iibox_address95 = zext_ln708_195_fu_11894_p1;

assign decipher_0_iibox_address96 = zext_ln708_178_fu_10782_p1;

assign decipher_0_iibox_address97 = zext_ln708_177_fu_10777_p1;

assign decipher_0_iibox_address98 = zext_ln708_176_fu_10772_p1;

assign decipher_0_iibox_address99 = zext_ln708_175_fu_10767_p1;

assign p_Result_25_fu_6039_p17 = {{{{{{{{{{{{{{{{decipher_0_iibox_q160}, {decipher_0_iibox_q161}}, {decipher_0_iibox_q162}}, {decipher_0_iibox_q163}}, {decipher_0_iibox_q164}}, {decipher_0_iibox_q165}}, {decipher_0_iibox_q166}}, {decipher_0_iibox_q167}}, {decipher_0_iibox_q168}}, {decipher_0_iibox_q169}}, {decipher_0_iibox_q170}}, {decipher_0_iibox_q171}}, {decipher_0_iibox_q172}}, {decipher_0_iibox_q173}}, {decipher_0_iibox_q174}}, {decipher_0_iibox_q175}};

assign p_Result_26_fu_7226_p17 = {{{{{{{{{{{{{{{{decipher_0_iibox_q144}, {decipher_0_iibox_q145}}, {decipher_0_iibox_q146}}, {decipher_0_iibox_q147}}, {decipher_0_iibox_q148}}, {decipher_0_iibox_q149}}, {decipher_0_iibox_q150}}, {decipher_0_iibox_q151}}, {decipher_0_iibox_q152}}, {decipher_0_iibox_q153}}, {decipher_0_iibox_q154}}, {decipher_0_iibox_q155}}, {decipher_0_iibox_q156}}, {decipher_0_iibox_q157}}, {decipher_0_iibox_q158}}, {decipher_0_iibox_q159}};

assign p_Result_27_fu_8413_p17 = {{{{{{{{{{{{{{{{decipher_0_iibox_q128}, {decipher_0_iibox_q129}}, {decipher_0_iibox_q130}}, {decipher_0_iibox_q131}}, {decipher_0_iibox_q132}}, {decipher_0_iibox_q133}}, {decipher_0_iibox_q134}}, {decipher_0_iibox_q135}}, {decipher_0_iibox_q136}}, {decipher_0_iibox_q137}}, {decipher_0_iibox_q138}}, {decipher_0_iibox_q139}}, {decipher_0_iibox_q140}}, {decipher_0_iibox_q141}}, {decipher_0_iibox_q142}}, {decipher_0_iibox_q143}};

assign p_Result_28_fu_9600_p17 = {{{{{{{{{{{{{{{{decipher_0_iibox_q112}, {decipher_0_iibox_q113}}, {decipher_0_iibox_q114}}, {decipher_0_iibox_q115}}, {decipher_0_iibox_q116}}, {decipher_0_iibox_q117}}, {decipher_0_iibox_q118}}, {decipher_0_iibox_q119}}, {decipher_0_iibox_q120}}, {decipher_0_iibox_q121}}, {decipher_0_iibox_q122}}, {decipher_0_iibox_q123}}, {decipher_0_iibox_q124}}, {decipher_0_iibox_q125}}, {decipher_0_iibox_q126}}, {decipher_0_iibox_q127}};

assign p_Result_29_fu_10787_p17 = {{{{{{{{{{{{{{{{decipher_0_iibox_q96}, {decipher_0_iibox_q97}}, {decipher_0_iibox_q98}}, {decipher_0_iibox_q99}}, {decipher_0_iibox_q100}}, {decipher_0_iibox_q101}}, {decipher_0_iibox_q102}}, {decipher_0_iibox_q103}}, {decipher_0_iibox_q104}}, {decipher_0_iibox_q105}}, {decipher_0_iibox_q106}}, {decipher_0_iibox_q107}}, {decipher_0_iibox_q108}}, {decipher_0_iibox_q109}}, {decipher_0_iibox_q110}}, {decipher_0_iibox_q111}};

assign p_Result_30_fu_11974_p17 = {{{{{{{{{{{{{{{{decipher_0_iibox_q80}, {decipher_0_iibox_q81}}, {decipher_0_iibox_q82}}, {decipher_0_iibox_q83}}, {decipher_0_iibox_q84}}, {decipher_0_iibox_q85}}, {decipher_0_iibox_q86}}, {decipher_0_iibox_q87}}, {decipher_0_iibox_q88}}, {decipher_0_iibox_q89}}, {decipher_0_iibox_q90}}, {decipher_0_iibox_q91}}, {decipher_0_iibox_q92}}, {decipher_0_iibox_q93}}, {decipher_0_iibox_q94}}, {decipher_0_iibox_q95}};

assign p_Result_31_fu_13161_p17 = {{{{{{{{{{{{{{{{decipher_0_iibox_q64}, {decipher_0_iibox_q65}}, {decipher_0_iibox_q66}}, {decipher_0_iibox_q67}}, {decipher_0_iibox_q68}}, {decipher_0_iibox_q69}}, {decipher_0_iibox_q70}}, {decipher_0_iibox_q71}}, {decipher_0_iibox_q72}}, {decipher_0_iibox_q73}}, {decipher_0_iibox_q74}}, {decipher_0_iibox_q75}}, {decipher_0_iibox_q76}}, {decipher_0_iibox_q77}}, {decipher_0_iibox_q78}}, {decipher_0_iibox_q79}};

assign p_Result_32_fu_14348_p17 = {{{{{{{{{{{{{{{{decipher_0_iibox_q48}, {decipher_0_iibox_q49}}, {decipher_0_iibox_q50}}, {decipher_0_iibox_q51}}, {decipher_0_iibox_q52}}, {decipher_0_iibox_q53}}, {decipher_0_iibox_q54}}, {decipher_0_iibox_q55}}, {decipher_0_iibox_q56}}, {decipher_0_iibox_q57}}, {decipher_0_iibox_q58}}, {decipher_0_iibox_q59}}, {decipher_0_iibox_q60}}, {decipher_0_iibox_q61}}, {decipher_0_iibox_q62}}, {decipher_0_iibox_q63}};

assign p_Result_33_fu_15535_p17 = {{{{{{{{{{{{{{{{decipher_0_iibox_q32}, {decipher_0_iibox_q33}}, {decipher_0_iibox_q34}}, {decipher_0_iibox_q35}}, {decipher_0_iibox_q36}}, {decipher_0_iibox_q37}}, {decipher_0_iibox_q38}}, {decipher_0_iibox_q39}}, {decipher_0_iibox_q40}}, {decipher_0_iibox_q41}}, {decipher_0_iibox_q42}}, {decipher_0_iibox_q43}}, {decipher_0_iibox_q44}}, {decipher_0_iibox_q45}}, {decipher_0_iibox_q46}}, {decipher_0_iibox_q47}};

assign p_Result_34_fu_16722_p17 = {{{{{{{{{{{{{{{{decipher_0_iibox_q16}, {decipher_0_iibox_q17}}, {decipher_0_iibox_q18}}, {decipher_0_iibox_q19}}, {decipher_0_iibox_q20}}, {decipher_0_iibox_q21}}, {decipher_0_iibox_q22}}, {decipher_0_iibox_q23}}, {decipher_0_iibox_q24}}, {decipher_0_iibox_q25}}, {decipher_0_iibox_q26}}, {decipher_0_iibox_q27}}, {decipher_0_iibox_q28}}, {decipher_0_iibox_q29}}, {decipher_0_iibox_q30}}, {decipher_0_iibox_q31}};

assign p_Result_35_fu_17909_p17 = {{{{{{{{{{{{{{{{decipher_0_iibox_q0}, {decipher_0_iibox_q1}}, {decipher_0_iibox_q2}}, {decipher_0_iibox_q3}}, {decipher_0_iibox_q4}}, {decipher_0_iibox_q5}}, {decipher_0_iibox_q6}}, {decipher_0_iibox_q7}}, {decipher_0_iibox_q8}}, {decipher_0_iibox_q9}}, {decipher_0_iibox_q10}}, {decipher_0_iibox_q11}}, {decipher_0_iibox_q12}}, {decipher_0_iibox_q13}}, {decipher_0_iibox_q14}}, {decipher_0_iibox_q15}};

assign p_Result_s_fu_4852_p17 = {{{{{{{{{{{{{{{{decipher_0_iibox_q176}, {decipher_0_iibox_q177}}, {decipher_0_iibox_q178}}, {decipher_0_iibox_q179}}, {decipher_0_iibox_q180}}, {decipher_0_iibox_q181}}, {decipher_0_iibox_q182}}, {decipher_0_iibox_q183}}, {decipher_0_iibox_q184}}, {decipher_0_iibox_q185}}, {decipher_0_iibox_q186}}, {decipher_0_iibox_q187}}, {decipher_0_iibox_q188}}, {decipher_0_iibox_q189}}, {decipher_0_iibox_q190}}, {decipher_0_iibox_q191}};

assign ret_V_fu_4612_p2 = (p_read12 ^ ciphertext);

assign state_V_24_fu_4888_p2 = (p_read_2_reg_17950 ^ p_Result_s_fu_4852_p17);

assign state_V_25_fu_6075_p2 = (p_read_3_reg_17955_pp0_iter2_reg ^ p_Result_25_fu_6039_p17);

assign state_V_26_fu_7262_p2 = (p_read_4_reg_17960_pp0_iter4_reg ^ p_Result_26_fu_7226_p17);

assign state_V_27_fu_8449_p2 = (p_read_5_reg_17965_pp0_iter6_reg ^ p_Result_27_fu_8413_p17);

assign state_V_28_fu_9636_p2 = (p_read_6_reg_17970_pp0_iter8_reg ^ p_Result_28_fu_9600_p17);

assign state_V_29_fu_10823_p2 = (p_read_7_reg_17975_pp0_iter10_reg ^ p_Result_29_fu_10787_p17);

assign state_V_30_fu_13197_p2 = (p_read_9_reg_17985_pp0_iter14_reg ^ p_Result_31_fu_13161_p17);

assign state_V_31_fu_14384_p2 = (p_read_10_reg_17990_pp0_iter16_reg ^ p_Result_32_fu_14348_p17);

assign state_V_32_fu_15571_p2 = (p_read_11_reg_17995_pp0_iter18_reg ^ p_Result_33_fu_15535_p17);

assign state_V_33_fu_16758_p2 = (p_read_12_reg_18000_pp0_iter20_reg ^ p_Result_34_fu_16722_p17);

assign state_V_fu_12010_p2 = (p_read_8_reg_17980_pp0_iter12_reg ^ p_Result_30_fu_11974_p17);

assign tmp_100_fu_6396_p4 = {{decipher_0_i32box_q157[23:16]}};

assign tmp_101_fu_6406_p4 = {{decipher_0_i32box_q157[31:24]}};

assign tmp_102_fu_6119_p4 = {{state_V_25_fu_6075_p2[31:24]}};

assign tmp_103_fu_6420_p4 = {{decipher_0_i32box_q156[15:8]}};

assign tmp_104_fu_6430_p4 = {{decipher_0_i32box_q156[23:16]}};

assign tmp_105_fu_6440_p4 = {{decipher_0_i32box_q156[31:24]}};

assign tmp_106_fu_6134_p4 = {{state_V_25_fu_6075_p2[39:32]}};

assign tmp_107_fu_6454_p4 = {{decipher_0_i32box_q155[15:8]}};

assign tmp_108_fu_6464_p4 = {{decipher_0_i32box_q155[23:16]}};

assign tmp_109_fu_6474_p4 = {{decipher_0_i32box_q155[31:24]}};

assign tmp_110_fu_6149_p4 = {{state_V_25_fu_6075_p2[47:40]}};

assign tmp_111_fu_6488_p4 = {{decipher_0_i32box_q154[15:8]}};

assign tmp_112_fu_6498_p4 = {{decipher_0_i32box_q154[23:16]}};

assign tmp_113_fu_6508_p4 = {{decipher_0_i32box_q154[31:24]}};

assign tmp_114_fu_6164_p4 = {{state_V_25_fu_6075_p2[55:48]}};

assign tmp_115_fu_6522_p4 = {{decipher_0_i32box_q153[15:8]}};

assign tmp_116_fu_6532_p4 = {{decipher_0_i32box_q153[23:16]}};

assign tmp_117_fu_6542_p4 = {{decipher_0_i32box_q153[31:24]}};

assign tmp_118_fu_6179_p4 = {{state_V_25_fu_6075_p2[63:56]}};

assign tmp_119_fu_6556_p4 = {{decipher_0_i32box_q152[15:8]}};

assign tmp_120_fu_6566_p4 = {{decipher_0_i32box_q152[23:16]}};

assign tmp_121_fu_6576_p4 = {{decipher_0_i32box_q152[31:24]}};

assign tmp_122_fu_6194_p4 = {{state_V_25_fu_6075_p2[71:64]}};

assign tmp_123_fu_6590_p4 = {{decipher_0_i32box_q151[15:8]}};

assign tmp_124_fu_6600_p4 = {{decipher_0_i32box_q151[23:16]}};

assign tmp_125_fu_6610_p4 = {{decipher_0_i32box_q151[31:24]}};

assign tmp_126_fu_6209_p4 = {{state_V_25_fu_6075_p2[79:72]}};

assign tmp_127_fu_6624_p4 = {{decipher_0_i32box_q150[15:8]}};

assign tmp_128_fu_6634_p4 = {{decipher_0_i32box_q150[23:16]}};

assign tmp_129_fu_6644_p4 = {{decipher_0_i32box_q150[31:24]}};

assign tmp_130_fu_6224_p4 = {{state_V_25_fu_6075_p2[87:80]}};

assign tmp_131_fu_6658_p4 = {{decipher_0_i32box_q149[15:8]}};

assign tmp_132_fu_6668_p4 = {{decipher_0_i32box_q149[23:16]}};

assign tmp_133_fu_6678_p4 = {{decipher_0_i32box_q149[31:24]}};

assign tmp_134_fu_6239_p4 = {{state_V_25_fu_6075_p2[95:88]}};

assign tmp_135_fu_6692_p4 = {{decipher_0_i32box_q148[15:8]}};

assign tmp_136_fu_6702_p4 = {{decipher_0_i32box_q148[23:16]}};

assign tmp_137_fu_6712_p4 = {{decipher_0_i32box_q148[31:24]}};

assign tmp_138_fu_6254_p4 = {{state_V_25_fu_6075_p2[103:96]}};

assign tmp_139_fu_6726_p4 = {{decipher_0_i32box_q147[15:8]}};

assign tmp_140_fu_6736_p4 = {{decipher_0_i32box_q147[23:16]}};

assign tmp_141_fu_6746_p4 = {{decipher_0_i32box_q147[31:24]}};

assign tmp_142_fu_6269_p4 = {{state_V_25_fu_6075_p2[111:104]}};

assign tmp_143_fu_6760_p4 = {{decipher_0_i32box_q146[15:8]}};

assign tmp_144_fu_6770_p4 = {{decipher_0_i32box_q146[23:16]}};

assign tmp_145_fu_6780_p4 = {{decipher_0_i32box_q146[31:24]}};

assign tmp_146_fu_6284_p4 = {{state_V_25_fu_6075_p2[119:112]}};

assign tmp_147_fu_6794_p4 = {{decipher_0_i32box_q145[15:8]}};

assign tmp_148_fu_6804_p4 = {{decipher_0_i32box_q145[23:16]}};

assign tmp_149_fu_6814_p4 = {{decipher_0_i32box_q145[31:24]}};

assign tmp_14_fu_4642_p4 = {{ret_V_fu_4612_p2[87:80]}};

assign tmp_150_fu_6299_p4 = {{state_V_25_fu_6075_p2[127:120]}};

assign tmp_151_fu_6828_p4 = {{decipher_0_i32box_q144[15:8]}};

assign tmp_152_fu_6838_p4 = {{decipher_0_i32box_q144[23:16]}};

assign tmp_153_fu_6848_p4 = {{decipher_0_i32box_q144[31:24]}};

assign tmp_154_fu_7505_p4 = {{decipher_0_i32box_q143[15:8]}};

assign tmp_155_fu_7515_p4 = {{decipher_0_i32box_q143[23:16]}};

assign tmp_156_fu_7525_p4 = {{decipher_0_i32box_q143[31:24]}};

assign tmp_157_fu_7276_p4 = {{state_V_26_fu_7262_p2[15:8]}};

assign tmp_158_fu_7539_p4 = {{decipher_0_i32box_q142[15:8]}};

assign tmp_159_fu_7549_p4 = {{decipher_0_i32box_q142[23:16]}};

assign tmp_15_fu_4657_p4 = {{ret_V_fu_4612_p2[63:56]}};

assign tmp_160_fu_7559_p4 = {{decipher_0_i32box_q142[31:24]}};

assign tmp_161_fu_7291_p4 = {{state_V_26_fu_7262_p2[23:16]}};

assign tmp_162_fu_7573_p4 = {{decipher_0_i32box_q141[15:8]}};

assign tmp_163_fu_7583_p4 = {{decipher_0_i32box_q141[23:16]}};

assign tmp_164_fu_7593_p4 = {{decipher_0_i32box_q141[31:24]}};

assign tmp_165_fu_7306_p4 = {{state_V_26_fu_7262_p2[31:24]}};

assign tmp_166_fu_7607_p4 = {{decipher_0_i32box_q140[15:8]}};

assign tmp_167_fu_7617_p4 = {{decipher_0_i32box_q140[23:16]}};

assign tmp_168_fu_7627_p4 = {{decipher_0_i32box_q140[31:24]}};

assign tmp_169_fu_7321_p4 = {{state_V_26_fu_7262_p2[39:32]}};

assign tmp_16_fu_4672_p4 = {{ret_V_fu_4612_p2[39:32]}};

assign tmp_170_fu_7641_p4 = {{decipher_0_i32box_q139[15:8]}};

assign tmp_171_fu_7651_p4 = {{decipher_0_i32box_q139[23:16]}};

assign tmp_172_fu_7661_p4 = {{decipher_0_i32box_q139[31:24]}};

assign tmp_173_fu_7336_p4 = {{state_V_26_fu_7262_p2[47:40]}};

assign tmp_174_fu_7675_p4 = {{decipher_0_i32box_q138[15:8]}};

assign tmp_175_fu_7685_p4 = {{decipher_0_i32box_q138[23:16]}};

assign tmp_176_fu_7695_p4 = {{decipher_0_i32box_q138[31:24]}};

assign tmp_177_fu_7351_p4 = {{state_V_26_fu_7262_p2[55:48]}};

assign tmp_178_fu_7709_p4 = {{decipher_0_i32box_q137[15:8]}};

assign tmp_179_fu_7719_p4 = {{decipher_0_i32box_q137[23:16]}};

assign tmp_17_fu_4687_p4 = {{ret_V_fu_4612_p2[15:8]}};

assign tmp_180_fu_7729_p4 = {{decipher_0_i32box_q137[31:24]}};

assign tmp_181_fu_7366_p4 = {{state_V_26_fu_7262_p2[63:56]}};

assign tmp_182_fu_7743_p4 = {{decipher_0_i32box_q136[15:8]}};

assign tmp_183_fu_7753_p4 = {{decipher_0_i32box_q136[23:16]}};

assign tmp_184_fu_7763_p4 = {{decipher_0_i32box_q136[31:24]}};

assign tmp_185_fu_7381_p4 = {{state_V_26_fu_7262_p2[71:64]}};

assign tmp_186_fu_7777_p4 = {{decipher_0_i32box_q135[15:8]}};

assign tmp_187_fu_7787_p4 = {{decipher_0_i32box_q135[23:16]}};

assign tmp_188_fu_7797_p4 = {{decipher_0_i32box_q135[31:24]}};

assign tmp_189_fu_7396_p4 = {{state_V_26_fu_7262_p2[79:72]}};

assign tmp_18_fu_4702_p4 = {{ret_V_fu_4612_p2[119:112]}};

assign tmp_190_fu_7811_p4 = {{decipher_0_i32box_q134[15:8]}};

assign tmp_191_fu_7821_p4 = {{decipher_0_i32box_q134[23:16]}};

assign tmp_192_fu_7831_p4 = {{decipher_0_i32box_q134[31:24]}};

assign tmp_193_fu_7411_p4 = {{state_V_26_fu_7262_p2[87:80]}};

assign tmp_194_fu_7845_p4 = {{decipher_0_i32box_q133[15:8]}};

assign tmp_195_fu_7855_p4 = {{decipher_0_i32box_q133[23:16]}};

assign tmp_196_fu_7865_p4 = {{decipher_0_i32box_q133[31:24]}};

assign tmp_197_fu_7426_p4 = {{state_V_26_fu_7262_p2[95:88]}};

assign tmp_198_fu_7879_p4 = {{decipher_0_i32box_q132[15:8]}};

assign tmp_199_fu_7889_p4 = {{decipher_0_i32box_q132[23:16]}};

assign tmp_19_fu_4717_p4 = {{ret_V_fu_4612_p2[95:88]}};

assign tmp_1_V_10_fu_17787_p2 = (xor_ln1545_526_fu_17781_p2 ^ xor_ln1545_525_fu_17775_p2);

assign tmp_1_V_1_fu_7104_p2 = (xor_ln1545_94_fu_7098_p2 ^ xor_ln1545_93_fu_7092_p2);

assign tmp_1_V_2_fu_8291_p2 = (xor_ln1545_142_fu_8285_p2 ^ xor_ln1545_141_fu_8279_p2);

assign tmp_1_V_3_fu_9478_p2 = (xor_ln1545_190_fu_9472_p2 ^ xor_ln1545_189_fu_9466_p2);

assign tmp_1_V_4_fu_10665_p2 = (xor_ln1545_238_fu_10659_p2 ^ xor_ln1545_237_fu_10653_p2);

assign tmp_1_V_5_fu_11852_p2 = (xor_ln1545_286_fu_11846_p2 ^ xor_ln1545_285_fu_11840_p2);

assign tmp_1_V_6_fu_13039_p2 = (xor_ln1545_334_fu_13033_p2 ^ xor_ln1545_333_fu_13027_p2);

assign tmp_1_V_7_fu_14226_p2 = (xor_ln1545_382_fu_14220_p2 ^ xor_ln1545_381_fu_14214_p2);

assign tmp_1_V_8_fu_15413_p2 = (xor_ln1545_430_fu_15407_p2 ^ xor_ln1545_429_fu_15401_p2);

assign tmp_1_V_9_fu_16600_p2 = (xor_ln1545_478_fu_16594_p2 ^ xor_ln1545_477_fu_16588_p2);

assign tmp_1_V_fu_5917_p2 = (xor_ln1545_46_fu_5911_p2 ^ xor_ln1545_45_fu_5905_p2);

assign tmp_200_fu_7899_p4 = {{decipher_0_i32box_q132[31:24]}};

assign tmp_201_fu_7441_p4 = {{state_V_26_fu_7262_p2[103:96]}};

assign tmp_202_fu_7913_p4 = {{decipher_0_i32box_q131[15:8]}};

assign tmp_203_fu_7923_p4 = {{decipher_0_i32box_q131[23:16]}};

assign tmp_204_fu_7933_p4 = {{decipher_0_i32box_q131[31:24]}};

assign tmp_205_fu_7456_p4 = {{state_V_26_fu_7262_p2[111:104]}};

assign tmp_206_fu_7947_p4 = {{decipher_0_i32box_q130[15:8]}};

assign tmp_207_fu_7957_p4 = {{decipher_0_i32box_q130[23:16]}};

assign tmp_208_fu_7967_p4 = {{decipher_0_i32box_q130[31:24]}};

assign tmp_209_fu_7471_p4 = {{state_V_26_fu_7262_p2[119:112]}};

assign tmp_20_fu_4732_p4 = {{ret_V_fu_4612_p2[71:64]}};

assign tmp_210_fu_7981_p4 = {{decipher_0_i32box_q129[15:8]}};

assign tmp_211_fu_7991_p4 = {{decipher_0_i32box_q129[23:16]}};

assign tmp_212_fu_8001_p4 = {{decipher_0_i32box_q129[31:24]}};

assign tmp_213_fu_7486_p4 = {{state_V_26_fu_7262_p2[127:120]}};

assign tmp_214_fu_8015_p4 = {{decipher_0_i32box_q128[15:8]}};

assign tmp_215_fu_8025_p4 = {{decipher_0_i32box_q128[23:16]}};

assign tmp_216_fu_8035_p4 = {{decipher_0_i32box_q128[31:24]}};

assign tmp_217_fu_8692_p4 = {{decipher_0_i32box_q127[15:8]}};

assign tmp_218_fu_8702_p4 = {{decipher_0_i32box_q127[23:16]}};

assign tmp_219_fu_8712_p4 = {{decipher_0_i32box_q127[31:24]}};

assign tmp_21_fu_4747_p4 = {{ret_V_fu_4612_p2[47:40]}};

assign tmp_220_fu_8463_p4 = {{state_V_27_fu_8449_p2[15:8]}};

assign tmp_221_fu_8726_p4 = {{decipher_0_i32box_q126[15:8]}};

assign tmp_222_fu_8736_p4 = {{decipher_0_i32box_q126[23:16]}};

assign tmp_223_fu_8746_p4 = {{decipher_0_i32box_q126[31:24]}};

assign tmp_224_fu_8478_p4 = {{state_V_27_fu_8449_p2[23:16]}};

assign tmp_225_fu_8760_p4 = {{decipher_0_i32box_q125[15:8]}};

assign tmp_226_fu_8770_p4 = {{decipher_0_i32box_q125[23:16]}};

assign tmp_227_fu_8780_p4 = {{decipher_0_i32box_q125[31:24]}};

assign tmp_228_fu_8493_p4 = {{state_V_27_fu_8449_p2[31:24]}};

assign tmp_229_fu_8794_p4 = {{decipher_0_i32box_q124[15:8]}};

assign tmp_22_fu_4762_p4 = {{ret_V_fu_4612_p2[23:16]}};

assign tmp_230_fu_8804_p4 = {{decipher_0_i32box_q124[23:16]}};

assign tmp_231_fu_8814_p4 = {{decipher_0_i32box_q124[31:24]}};

assign tmp_232_fu_8508_p4 = {{state_V_27_fu_8449_p2[39:32]}};

assign tmp_233_fu_8828_p4 = {{decipher_0_i32box_q123[15:8]}};

assign tmp_234_fu_8838_p4 = {{decipher_0_i32box_q123[23:16]}};

assign tmp_235_fu_8848_p4 = {{decipher_0_i32box_q123[31:24]}};

assign tmp_236_fu_8523_p4 = {{state_V_27_fu_8449_p2[47:40]}};

assign tmp_237_fu_8862_p4 = {{decipher_0_i32box_q122[15:8]}};

assign tmp_238_fu_8872_p4 = {{decipher_0_i32box_q122[23:16]}};

assign tmp_239_fu_8882_p4 = {{decipher_0_i32box_q122[31:24]}};

assign tmp_23_fu_4777_p4 = {{ret_V_fu_4612_p2[127:120]}};

assign tmp_240_fu_8538_p4 = {{state_V_27_fu_8449_p2[55:48]}};

assign tmp_241_fu_8896_p4 = {{decipher_0_i32box_q121[15:8]}};

assign tmp_242_fu_8906_p4 = {{decipher_0_i32box_q121[23:16]}};

assign tmp_243_fu_8916_p4 = {{decipher_0_i32box_q121[31:24]}};

assign tmp_244_fu_8553_p4 = {{state_V_27_fu_8449_p2[63:56]}};

assign tmp_245_fu_8930_p4 = {{decipher_0_i32box_q120[15:8]}};

assign tmp_246_fu_8940_p4 = {{decipher_0_i32box_q120[23:16]}};

assign tmp_247_fu_8950_p4 = {{decipher_0_i32box_q120[31:24]}};

assign tmp_248_fu_8568_p4 = {{state_V_27_fu_8449_p2[71:64]}};

assign tmp_249_fu_8964_p4 = {{decipher_0_i32box_q119[15:8]}};

assign tmp_24_fu_4792_p4 = {{ret_V_fu_4612_p2[103:96]}};

assign tmp_250_fu_8974_p4 = {{decipher_0_i32box_q119[23:16]}};

assign tmp_251_fu_8984_p4 = {{decipher_0_i32box_q119[31:24]}};

assign tmp_252_fu_8583_p4 = {{state_V_27_fu_8449_p2[79:72]}};

assign tmp_253_fu_8998_p4 = {{decipher_0_i32box_q118[15:8]}};

assign tmp_254_fu_9008_p4 = {{decipher_0_i32box_q118[23:16]}};

assign tmp_255_fu_9018_p4 = {{decipher_0_i32box_q118[31:24]}};

assign tmp_256_fu_8598_p4 = {{state_V_27_fu_8449_p2[87:80]}};

assign tmp_257_fu_9032_p4 = {{decipher_0_i32box_q117[15:8]}};

assign tmp_258_fu_9042_p4 = {{decipher_0_i32box_q117[23:16]}};

assign tmp_259_fu_9052_p4 = {{decipher_0_i32box_q117[31:24]}};

assign tmp_25_fu_4807_p4 = {{ret_V_fu_4612_p2[79:72]}};

assign tmp_260_fu_8613_p4 = {{state_V_27_fu_8449_p2[95:88]}};

assign tmp_261_fu_9066_p4 = {{decipher_0_i32box_q116[15:8]}};

assign tmp_262_fu_9076_p4 = {{decipher_0_i32box_q116[23:16]}};

assign tmp_263_fu_9086_p4 = {{decipher_0_i32box_q116[31:24]}};

assign tmp_264_fu_8628_p4 = {{state_V_27_fu_8449_p2[103:96]}};

assign tmp_265_fu_9100_p4 = {{decipher_0_i32box_q115[15:8]}};

assign tmp_266_fu_9110_p4 = {{decipher_0_i32box_q115[23:16]}};

assign tmp_267_fu_9120_p4 = {{decipher_0_i32box_q115[31:24]}};

assign tmp_268_fu_8643_p4 = {{state_V_27_fu_8449_p2[111:104]}};

assign tmp_269_fu_9134_p4 = {{decipher_0_i32box_q114[15:8]}};

assign tmp_26_fu_4822_p4 = {{ret_V_fu_4612_p2[55:48]}};

assign tmp_270_fu_9144_p4 = {{decipher_0_i32box_q114[23:16]}};

assign tmp_271_fu_9154_p4 = {{decipher_0_i32box_q114[31:24]}};

assign tmp_272_fu_8658_p4 = {{state_V_27_fu_8449_p2[119:112]}};

assign tmp_273_fu_9168_p4 = {{decipher_0_i32box_q113[15:8]}};

assign tmp_274_fu_9178_p4 = {{decipher_0_i32box_q113[23:16]}};

assign tmp_275_fu_9188_p4 = {{decipher_0_i32box_q113[31:24]}};

assign tmp_276_fu_8673_p4 = {{state_V_27_fu_8449_p2[127:120]}};

assign tmp_277_fu_9202_p4 = {{decipher_0_i32box_q112[15:8]}};

assign tmp_278_fu_9212_p4 = {{decipher_0_i32box_q112[23:16]}};

assign tmp_279_fu_9222_p4 = {{decipher_0_i32box_q112[31:24]}};

assign tmp_27_fu_4837_p4 = {{ret_V_fu_4612_p2[31:24]}};

assign tmp_280_fu_9879_p4 = {{decipher_0_i32box_q111[15:8]}};

assign tmp_281_fu_9889_p4 = {{decipher_0_i32box_q111[23:16]}};

assign tmp_282_fu_9899_p4 = {{decipher_0_i32box_q111[31:24]}};

assign tmp_283_fu_9650_p4 = {{state_V_28_fu_9636_p2[15:8]}};

assign tmp_284_fu_9913_p4 = {{decipher_0_i32box_q110[15:8]}};

assign tmp_285_fu_9923_p4 = {{decipher_0_i32box_q110[23:16]}};

assign tmp_286_fu_9933_p4 = {{decipher_0_i32box_q110[31:24]}};

assign tmp_287_fu_9665_p4 = {{state_V_28_fu_9636_p2[23:16]}};

assign tmp_288_fu_9947_p4 = {{decipher_0_i32box_q109[15:8]}};

assign tmp_289_fu_9957_p4 = {{decipher_0_i32box_q109[23:16]}};

assign tmp_28_fu_5131_p4 = {{decipher_0_i32box_q175[15:8]}};

assign tmp_290_fu_9967_p4 = {{decipher_0_i32box_q109[31:24]}};

assign tmp_291_fu_9680_p4 = {{state_V_28_fu_9636_p2[31:24]}};

assign tmp_292_fu_9981_p4 = {{decipher_0_i32box_q108[15:8]}};

assign tmp_293_fu_9991_p4 = {{decipher_0_i32box_q108[23:16]}};

assign tmp_294_fu_10001_p4 = {{decipher_0_i32box_q108[31:24]}};

assign tmp_295_fu_9695_p4 = {{state_V_28_fu_9636_p2[39:32]}};

assign tmp_296_fu_10015_p4 = {{decipher_0_i32box_q107[15:8]}};

assign tmp_297_fu_10025_p4 = {{decipher_0_i32box_q107[23:16]}};

assign tmp_298_fu_10035_p4 = {{decipher_0_i32box_q107[31:24]}};

assign tmp_299_fu_9710_p4 = {{state_V_28_fu_9636_p2[47:40]}};

assign tmp_29_fu_5141_p4 = {{decipher_0_i32box_q175[23:16]}};

assign tmp_2_1_V_10_fu_17733_p2 = (xor_ln1545_517_fu_17727_p2 ^ xor_ln1545_516_fu_17721_p2);

assign tmp_2_1_V_1_fu_7050_p2 = (xor_ln1545_85_fu_7044_p2 ^ xor_ln1545_84_fu_7038_p2);

assign tmp_2_1_V_2_fu_8237_p2 = (xor_ln1545_133_fu_8231_p2 ^ xor_ln1545_132_fu_8225_p2);

assign tmp_2_1_V_3_fu_9424_p2 = (xor_ln1545_181_fu_9418_p2 ^ xor_ln1545_180_fu_9412_p2);

assign tmp_2_1_V_4_fu_10611_p2 = (xor_ln1545_229_fu_10605_p2 ^ xor_ln1545_228_fu_10599_p2);

assign tmp_2_1_V_5_fu_11798_p2 = (xor_ln1545_277_fu_11792_p2 ^ xor_ln1545_276_fu_11786_p2);

assign tmp_2_1_V_6_fu_12985_p2 = (xor_ln1545_325_fu_12979_p2 ^ xor_ln1545_324_fu_12973_p2);

assign tmp_2_1_V_7_fu_14172_p2 = (xor_ln1545_373_fu_14166_p2 ^ xor_ln1545_372_fu_14160_p2);

assign tmp_2_1_V_8_fu_15359_p2 = (xor_ln1545_421_fu_15353_p2 ^ xor_ln1545_420_fu_15347_p2);

assign tmp_2_1_V_9_fu_16546_p2 = (xor_ln1545_469_fu_16540_p2 ^ xor_ln1545_468_fu_16534_p2);

assign tmp_2_1_V_fu_5863_p2 = (xor_ln1545_37_fu_5857_p2 ^ xor_ln1545_36_fu_5851_p2);

assign tmp_2_2_V_10_fu_17805_p2 = (xor_ln1545_529_fu_17799_p2 ^ xor_ln1545_528_fu_17793_p2);

assign tmp_2_2_V_1_fu_7122_p2 = (xor_ln1545_97_fu_7116_p2 ^ xor_ln1545_96_fu_7110_p2);

assign tmp_2_2_V_2_fu_8309_p2 = (xor_ln1545_145_fu_8303_p2 ^ xor_ln1545_144_fu_8297_p2);

assign tmp_2_2_V_3_fu_9496_p2 = (xor_ln1545_193_fu_9490_p2 ^ xor_ln1545_192_fu_9484_p2);

assign tmp_2_2_V_4_fu_10683_p2 = (xor_ln1545_241_fu_10677_p2 ^ xor_ln1545_240_fu_10671_p2);

assign tmp_2_2_V_5_fu_11870_p2 = (xor_ln1545_289_fu_11864_p2 ^ xor_ln1545_288_fu_11858_p2);

assign tmp_2_2_V_6_fu_13057_p2 = (xor_ln1545_337_fu_13051_p2 ^ xor_ln1545_336_fu_13045_p2);

assign tmp_2_2_V_7_fu_14244_p2 = (xor_ln1545_385_fu_14238_p2 ^ xor_ln1545_384_fu_14232_p2);

assign tmp_2_2_V_8_fu_15431_p2 = (xor_ln1545_433_fu_15425_p2 ^ xor_ln1545_432_fu_15419_p2);

assign tmp_2_2_V_9_fu_16618_p2 = (xor_ln1545_481_fu_16612_p2 ^ xor_ln1545_480_fu_16606_p2);

assign tmp_2_2_V_fu_5935_p2 = (xor_ln1545_49_fu_5929_p2 ^ xor_ln1545_48_fu_5923_p2);

assign tmp_300_fu_10049_p4 = {{decipher_0_i32box_q106[15:8]}};

assign tmp_301_fu_10059_p4 = {{decipher_0_i32box_q106[23:16]}};

assign tmp_302_fu_10069_p4 = {{decipher_0_i32box_q106[31:24]}};

assign tmp_303_fu_9725_p4 = {{state_V_28_fu_9636_p2[55:48]}};

assign tmp_304_fu_10083_p4 = {{decipher_0_i32box_q105[15:8]}};

assign tmp_305_fu_10093_p4 = {{decipher_0_i32box_q105[23:16]}};

assign tmp_306_fu_10103_p4 = {{decipher_0_i32box_q105[31:24]}};

assign tmp_307_fu_9740_p4 = {{state_V_28_fu_9636_p2[63:56]}};

assign tmp_308_fu_10117_p4 = {{decipher_0_i32box_q104[15:8]}};

assign tmp_309_fu_10127_p4 = {{decipher_0_i32box_q104[23:16]}};

assign tmp_30_fu_5151_p4 = {{decipher_0_i32box_q175[31:24]}};

assign tmp_310_fu_10137_p4 = {{decipher_0_i32box_q104[31:24]}};

assign tmp_311_fu_9755_p4 = {{state_V_28_fu_9636_p2[71:64]}};

assign tmp_312_fu_10151_p4 = {{decipher_0_i32box_q103[15:8]}};

assign tmp_313_fu_10161_p4 = {{decipher_0_i32box_q103[23:16]}};

assign tmp_314_fu_10171_p4 = {{decipher_0_i32box_q103[31:24]}};

assign tmp_315_fu_9770_p4 = {{state_V_28_fu_9636_p2[79:72]}};

assign tmp_316_fu_10185_p4 = {{decipher_0_i32box_q102[15:8]}};

assign tmp_317_fu_10195_p4 = {{decipher_0_i32box_q102[23:16]}};

assign tmp_318_fu_10205_p4 = {{decipher_0_i32box_q102[31:24]}};

assign tmp_319_fu_9785_p4 = {{state_V_28_fu_9636_p2[87:80]}};

assign tmp_31_fu_4902_p4 = {{state_V_24_fu_4888_p2[15:8]}};

assign tmp_320_fu_10219_p4 = {{decipher_0_i32box_q101[15:8]}};

assign tmp_321_fu_10229_p4 = {{decipher_0_i32box_q101[23:16]}};

assign tmp_322_fu_10239_p4 = {{decipher_0_i32box_q101[31:24]}};

assign tmp_323_fu_9800_p4 = {{state_V_28_fu_9636_p2[95:88]}};

assign tmp_324_fu_10253_p4 = {{decipher_0_i32box_q100[15:8]}};

assign tmp_325_fu_10263_p4 = {{decipher_0_i32box_q100[23:16]}};

assign tmp_326_fu_10273_p4 = {{decipher_0_i32box_q100[31:24]}};

assign tmp_327_fu_9815_p4 = {{state_V_28_fu_9636_p2[103:96]}};

assign tmp_328_fu_10287_p4 = {{decipher_0_i32box_q99[15:8]}};

assign tmp_329_fu_10297_p4 = {{decipher_0_i32box_q99[23:16]}};

assign tmp_32_fu_5165_p4 = {{decipher_0_i32box_q174[15:8]}};

assign tmp_330_fu_10307_p4 = {{decipher_0_i32box_q99[31:24]}};

assign tmp_331_fu_9830_p4 = {{state_V_28_fu_9636_p2[111:104]}};

assign tmp_332_fu_10321_p4 = {{decipher_0_i32box_q98[15:8]}};

assign tmp_333_fu_10331_p4 = {{decipher_0_i32box_q98[23:16]}};

assign tmp_334_fu_10341_p4 = {{decipher_0_i32box_q98[31:24]}};

assign tmp_335_fu_9845_p4 = {{state_V_28_fu_9636_p2[119:112]}};

assign tmp_336_fu_10355_p4 = {{decipher_0_i32box_q97[15:8]}};

assign tmp_337_fu_10365_p4 = {{decipher_0_i32box_q97[23:16]}};

assign tmp_338_fu_10375_p4 = {{decipher_0_i32box_q97[31:24]}};

assign tmp_339_fu_9860_p4 = {{state_V_28_fu_9636_p2[127:120]}};

assign tmp_33_fu_5175_p4 = {{decipher_0_i32box_q174[23:16]}};

assign tmp_340_fu_10389_p4 = {{decipher_0_i32box_q96[15:8]}};

assign tmp_341_fu_10399_p4 = {{decipher_0_i32box_q96[23:16]}};

assign tmp_342_fu_10409_p4 = {{decipher_0_i32box_q96[31:24]}};

assign tmp_343_fu_11066_p4 = {{decipher_0_i32box_q95[15:8]}};

assign tmp_344_fu_11076_p4 = {{decipher_0_i32box_q95[23:16]}};

assign tmp_345_fu_11086_p4 = {{decipher_0_i32box_q95[31:24]}};

assign tmp_346_fu_10837_p4 = {{state_V_29_fu_10823_p2[15:8]}};

assign tmp_347_fu_11100_p4 = {{decipher_0_i32box_q94[15:8]}};

assign tmp_348_fu_11110_p4 = {{decipher_0_i32box_q94[23:16]}};

assign tmp_349_fu_11120_p4 = {{decipher_0_i32box_q94[31:24]}};

assign tmp_34_fu_5185_p4 = {{decipher_0_i32box_q174[31:24]}};

assign tmp_350_fu_10852_p4 = {{state_V_29_fu_10823_p2[23:16]}};

assign tmp_351_fu_11134_p4 = {{decipher_0_i32box_q93[15:8]}};

assign tmp_352_fu_11144_p4 = {{decipher_0_i32box_q93[23:16]}};

assign tmp_353_fu_11154_p4 = {{decipher_0_i32box_q93[31:24]}};

assign tmp_354_fu_10867_p4 = {{state_V_29_fu_10823_p2[31:24]}};

assign tmp_355_fu_11168_p4 = {{decipher_0_i32box_q92[15:8]}};

assign tmp_356_fu_11178_p4 = {{decipher_0_i32box_q92[23:16]}};

assign tmp_357_fu_11188_p4 = {{decipher_0_i32box_q92[31:24]}};

assign tmp_358_fu_10882_p4 = {{state_V_29_fu_10823_p2[39:32]}};

assign tmp_359_fu_11202_p4 = {{decipher_0_i32box_q91[15:8]}};

assign tmp_35_fu_4917_p4 = {{state_V_24_fu_4888_p2[23:16]}};

assign tmp_360_fu_11212_p4 = {{decipher_0_i32box_q91[23:16]}};

assign tmp_361_fu_11222_p4 = {{decipher_0_i32box_q91[31:24]}};

assign tmp_362_fu_10897_p4 = {{state_V_29_fu_10823_p2[47:40]}};

assign tmp_363_fu_11236_p4 = {{decipher_0_i32box_q90[15:8]}};

assign tmp_364_fu_11246_p4 = {{decipher_0_i32box_q90[23:16]}};

assign tmp_365_fu_11256_p4 = {{decipher_0_i32box_q90[31:24]}};

assign tmp_366_fu_10912_p4 = {{state_V_29_fu_10823_p2[55:48]}};

assign tmp_367_fu_11270_p4 = {{decipher_0_i32box_q89[15:8]}};

assign tmp_368_fu_11280_p4 = {{decipher_0_i32box_q89[23:16]}};

assign tmp_369_fu_11290_p4 = {{decipher_0_i32box_q89[31:24]}};

assign tmp_36_fu_5199_p4 = {{decipher_0_i32box_q173[15:8]}};

assign tmp_370_fu_10927_p4 = {{state_V_29_fu_10823_p2[63:56]}};

assign tmp_371_fu_11304_p4 = {{decipher_0_i32box_q88[15:8]}};

assign tmp_372_fu_11314_p4 = {{decipher_0_i32box_q88[23:16]}};

assign tmp_373_fu_11324_p4 = {{decipher_0_i32box_q88[31:24]}};

assign tmp_374_fu_10942_p4 = {{state_V_29_fu_10823_p2[71:64]}};

assign tmp_375_fu_11338_p4 = {{decipher_0_i32box_q87[15:8]}};

assign tmp_376_fu_11348_p4 = {{decipher_0_i32box_q87[23:16]}};

assign tmp_377_fu_11358_p4 = {{decipher_0_i32box_q87[31:24]}};

assign tmp_378_fu_10957_p4 = {{state_V_29_fu_10823_p2[79:72]}};

assign tmp_379_fu_11372_p4 = {{decipher_0_i32box_q86[15:8]}};

assign tmp_37_fu_5209_p4 = {{decipher_0_i32box_q173[23:16]}};

assign tmp_380_fu_11382_p4 = {{decipher_0_i32box_q86[23:16]}};

assign tmp_381_fu_11392_p4 = {{decipher_0_i32box_q86[31:24]}};

assign tmp_382_fu_10972_p4 = {{state_V_29_fu_10823_p2[87:80]}};

assign tmp_383_fu_11406_p4 = {{decipher_0_i32box_q85[15:8]}};

assign tmp_384_fu_11416_p4 = {{decipher_0_i32box_q85[23:16]}};

assign tmp_385_fu_11426_p4 = {{decipher_0_i32box_q85[31:24]}};

assign tmp_386_fu_10987_p4 = {{state_V_29_fu_10823_p2[95:88]}};

assign tmp_387_fu_11440_p4 = {{decipher_0_i32box_q84[15:8]}};

assign tmp_388_fu_11450_p4 = {{decipher_0_i32box_q84[23:16]}};

assign tmp_389_fu_11460_p4 = {{decipher_0_i32box_q84[31:24]}};

assign tmp_38_fu_5219_p4 = {{decipher_0_i32box_q173[31:24]}};

assign tmp_390_fu_11002_p4 = {{state_V_29_fu_10823_p2[103:96]}};

assign tmp_391_fu_11474_p4 = {{decipher_0_i32box_q83[15:8]}};

assign tmp_392_fu_11484_p4 = {{decipher_0_i32box_q83[23:16]}};

assign tmp_393_fu_11494_p4 = {{decipher_0_i32box_q83[31:24]}};

assign tmp_394_fu_11017_p4 = {{state_V_29_fu_10823_p2[111:104]}};

assign tmp_395_fu_11508_p4 = {{decipher_0_i32box_q82[15:8]}};

assign tmp_396_fu_11518_p4 = {{decipher_0_i32box_q82[23:16]}};

assign tmp_397_fu_11528_p4 = {{decipher_0_i32box_q82[31:24]}};

assign tmp_398_fu_11032_p4 = {{state_V_29_fu_10823_p2[119:112]}};

assign tmp_399_fu_11542_p4 = {{decipher_0_i32box_q81[15:8]}};

assign tmp_39_fu_4932_p4 = {{state_V_24_fu_4888_p2[31:24]}};

assign tmp_3_V_10_fu_17607_p2 = (xor_ln1545_496_fu_17601_p2 ^ xor_ln1545_495_fu_17595_p2);

assign tmp_3_V_1_fu_6924_p2 = (xor_ln1545_64_fu_6918_p2 ^ xor_ln1545_63_fu_6912_p2);

assign tmp_3_V_2_fu_8111_p2 = (xor_ln1545_112_fu_8105_p2 ^ xor_ln1545_111_fu_8099_p2);

assign tmp_3_V_3_fu_9298_p2 = (xor_ln1545_160_fu_9292_p2 ^ xor_ln1545_159_fu_9286_p2);

assign tmp_3_V_4_fu_10485_p2 = (xor_ln1545_208_fu_10479_p2 ^ xor_ln1545_207_fu_10473_p2);

assign tmp_3_V_5_fu_11672_p2 = (xor_ln1545_256_fu_11666_p2 ^ xor_ln1545_255_fu_11660_p2);

assign tmp_3_V_6_fu_12859_p2 = (xor_ln1545_304_fu_12853_p2 ^ xor_ln1545_303_fu_12847_p2);

assign tmp_3_V_7_fu_14046_p2 = (xor_ln1545_352_fu_14040_p2 ^ xor_ln1545_351_fu_14034_p2);

assign tmp_3_V_8_fu_15233_p2 = (xor_ln1545_400_fu_15227_p2 ^ xor_ln1545_399_fu_15221_p2);

assign tmp_3_V_9_fu_16420_p2 = (xor_ln1545_448_fu_16414_p2 ^ xor_ln1545_447_fu_16408_p2);

assign tmp_3_V_fu_5737_p2 = (xor_ln1545_16_fu_5731_p2 ^ xor_ln1545_15_fu_5725_p2);

assign tmp_400_fu_11552_p4 = {{decipher_0_i32box_q81[23:16]}};

assign tmp_401_fu_11562_p4 = {{decipher_0_i32box_q81[31:24]}};

assign tmp_402_fu_11047_p4 = {{state_V_29_fu_10823_p2[127:120]}};

assign tmp_403_fu_11576_p4 = {{decipher_0_i32box_q80[15:8]}};

assign tmp_404_fu_11586_p4 = {{decipher_0_i32box_q80[23:16]}};

assign tmp_405_fu_11596_p4 = {{decipher_0_i32box_q80[31:24]}};

assign tmp_406_fu_12253_p4 = {{decipher_0_i32box_q79[15:8]}};

assign tmp_407_fu_12263_p4 = {{decipher_0_i32box_q79[23:16]}};

assign tmp_408_fu_12273_p4 = {{decipher_0_i32box_q79[31:24]}};

assign tmp_409_fu_12024_p4 = {{state_V_fu_12010_p2[15:8]}};

assign tmp_40_fu_5233_p4 = {{decipher_0_i32box_q172[15:8]}};

assign tmp_410_fu_12287_p4 = {{decipher_0_i32box_q78[15:8]}};

assign tmp_411_fu_12297_p4 = {{decipher_0_i32box_q78[23:16]}};

assign tmp_412_fu_12307_p4 = {{decipher_0_i32box_q78[31:24]}};

assign tmp_413_fu_12039_p4 = {{state_V_fu_12010_p2[23:16]}};

assign tmp_414_fu_12321_p4 = {{decipher_0_i32box_q77[15:8]}};

assign tmp_415_fu_12331_p4 = {{decipher_0_i32box_q77[23:16]}};

assign tmp_416_fu_12341_p4 = {{decipher_0_i32box_q77[31:24]}};

assign tmp_417_fu_12054_p4 = {{state_V_fu_12010_p2[31:24]}};

assign tmp_418_fu_12355_p4 = {{decipher_0_i32box_q76[15:8]}};

assign tmp_419_fu_12365_p4 = {{decipher_0_i32box_q76[23:16]}};

assign tmp_41_fu_5243_p4 = {{decipher_0_i32box_q172[23:16]}};

assign tmp_420_fu_12375_p4 = {{decipher_0_i32box_q76[31:24]}};

assign tmp_421_fu_12069_p4 = {{state_V_fu_12010_p2[39:32]}};

assign tmp_422_fu_12389_p4 = {{decipher_0_i32box_q75[15:8]}};

assign tmp_423_fu_12399_p4 = {{decipher_0_i32box_q75[23:16]}};

assign tmp_424_fu_12409_p4 = {{decipher_0_i32box_q75[31:24]}};

assign tmp_425_fu_12084_p4 = {{state_V_fu_12010_p2[47:40]}};

assign tmp_426_fu_12423_p4 = {{decipher_0_i32box_q74[15:8]}};

assign tmp_427_fu_12433_p4 = {{decipher_0_i32box_q74[23:16]}};

assign tmp_428_fu_12443_p4 = {{decipher_0_i32box_q74[31:24]}};

assign tmp_429_fu_12099_p4 = {{state_V_fu_12010_p2[55:48]}};

assign tmp_42_fu_5253_p4 = {{decipher_0_i32box_q172[31:24]}};

assign tmp_430_fu_12457_p4 = {{decipher_0_i32box_q73[15:8]}};

assign tmp_431_fu_12467_p4 = {{decipher_0_i32box_q73[23:16]}};

assign tmp_432_fu_12477_p4 = {{decipher_0_i32box_q73[31:24]}};

assign tmp_433_fu_12114_p4 = {{state_V_fu_12010_p2[63:56]}};

assign tmp_434_fu_12491_p4 = {{decipher_0_i32box_q72[15:8]}};

assign tmp_435_fu_12501_p4 = {{decipher_0_i32box_q72[23:16]}};

assign tmp_436_fu_12511_p4 = {{decipher_0_i32box_q72[31:24]}};

assign tmp_437_fu_12129_p4 = {{state_V_fu_12010_p2[71:64]}};

assign tmp_438_fu_12525_p4 = {{decipher_0_i32box_q71[15:8]}};

assign tmp_439_fu_12535_p4 = {{decipher_0_i32box_q71[23:16]}};

assign tmp_43_fu_4947_p4 = {{state_V_24_fu_4888_p2[39:32]}};

assign tmp_440_fu_12545_p4 = {{decipher_0_i32box_q71[31:24]}};

assign tmp_441_fu_12144_p4 = {{state_V_fu_12010_p2[79:72]}};

assign tmp_442_fu_12559_p4 = {{decipher_0_i32box_q70[15:8]}};

assign tmp_443_fu_12569_p4 = {{decipher_0_i32box_q70[23:16]}};

assign tmp_444_fu_12579_p4 = {{decipher_0_i32box_q70[31:24]}};

assign tmp_445_fu_12159_p4 = {{state_V_fu_12010_p2[87:80]}};

assign tmp_446_fu_12593_p4 = {{decipher_0_i32box_q69[15:8]}};

assign tmp_447_fu_12603_p4 = {{decipher_0_i32box_q69[23:16]}};

assign tmp_448_fu_12613_p4 = {{decipher_0_i32box_q69[31:24]}};

assign tmp_449_fu_12174_p4 = {{state_V_fu_12010_p2[95:88]}};

assign tmp_44_fu_5267_p4 = {{decipher_0_i32box_q171[15:8]}};

assign tmp_450_fu_12627_p4 = {{decipher_0_i32box_q68[15:8]}};

assign tmp_451_fu_12637_p4 = {{decipher_0_i32box_q68[23:16]}};

assign tmp_452_fu_12647_p4 = {{decipher_0_i32box_q68[31:24]}};

assign tmp_453_fu_12189_p4 = {{state_V_fu_12010_p2[103:96]}};

assign tmp_454_fu_12661_p4 = {{decipher_0_i32box_q67[15:8]}};

assign tmp_455_fu_12671_p4 = {{decipher_0_i32box_q67[23:16]}};

assign tmp_456_fu_12681_p4 = {{decipher_0_i32box_q67[31:24]}};

assign tmp_457_fu_12204_p4 = {{state_V_fu_12010_p2[111:104]}};

assign tmp_458_fu_12695_p4 = {{decipher_0_i32box_q66[15:8]}};

assign tmp_459_fu_12705_p4 = {{decipher_0_i32box_q66[23:16]}};

assign tmp_45_fu_5277_p4 = {{decipher_0_i32box_q171[23:16]}};

assign tmp_460_fu_12715_p4 = {{decipher_0_i32box_q66[31:24]}};

assign tmp_461_fu_12219_p4 = {{state_V_fu_12010_p2[119:112]}};

assign tmp_462_fu_12729_p4 = {{decipher_0_i32box_q65[15:8]}};

assign tmp_463_fu_12739_p4 = {{decipher_0_i32box_q65[23:16]}};

assign tmp_464_fu_12749_p4 = {{decipher_0_i32box_q65[31:24]}};

assign tmp_465_fu_12234_p4 = {{state_V_fu_12010_p2[127:120]}};

assign tmp_466_fu_12763_p4 = {{decipher_0_i32box_q64[15:8]}};

assign tmp_467_fu_12773_p4 = {{decipher_0_i32box_q64[23:16]}};

assign tmp_468_fu_12783_p4 = {{decipher_0_i32box_q64[31:24]}};

assign tmp_469_fu_13440_p4 = {{decipher_0_i32box_q63[15:8]}};

assign tmp_46_fu_5287_p4 = {{decipher_0_i32box_q171[31:24]}};

assign tmp_470_fu_13450_p4 = {{decipher_0_i32box_q63[23:16]}};

assign tmp_471_fu_13460_p4 = {{decipher_0_i32box_q63[31:24]}};

assign tmp_472_fu_13211_p4 = {{state_V_30_fu_13197_p2[15:8]}};

assign tmp_473_fu_13474_p4 = {{decipher_0_i32box_q62[15:8]}};

assign tmp_474_fu_13484_p4 = {{decipher_0_i32box_q62[23:16]}};

assign tmp_475_fu_13494_p4 = {{decipher_0_i32box_q62[31:24]}};

assign tmp_476_fu_13226_p4 = {{state_V_30_fu_13197_p2[23:16]}};

assign tmp_477_fu_13508_p4 = {{decipher_0_i32box_q61[15:8]}};

assign tmp_478_fu_13518_p4 = {{decipher_0_i32box_q61[23:16]}};

assign tmp_479_fu_13528_p4 = {{decipher_0_i32box_q61[31:24]}};

assign tmp_47_fu_4962_p4 = {{state_V_24_fu_4888_p2[47:40]}};

assign tmp_480_fu_13241_p4 = {{state_V_30_fu_13197_p2[31:24]}};

assign tmp_481_fu_13542_p4 = {{decipher_0_i32box_q60[15:8]}};

assign tmp_482_fu_13552_p4 = {{decipher_0_i32box_q60[23:16]}};

assign tmp_483_fu_13562_p4 = {{decipher_0_i32box_q60[31:24]}};

assign tmp_484_fu_13256_p4 = {{state_V_30_fu_13197_p2[39:32]}};

assign tmp_485_fu_13576_p4 = {{decipher_0_i32box_q59[15:8]}};

assign tmp_486_fu_13586_p4 = {{decipher_0_i32box_q59[23:16]}};

assign tmp_487_fu_13596_p4 = {{decipher_0_i32box_q59[31:24]}};

assign tmp_488_fu_13271_p4 = {{state_V_30_fu_13197_p2[47:40]}};

assign tmp_489_fu_13610_p4 = {{decipher_0_i32box_q58[15:8]}};

assign tmp_48_fu_5301_p4 = {{decipher_0_i32box_q170[15:8]}};

assign tmp_490_fu_13620_p4 = {{decipher_0_i32box_q58[23:16]}};

assign tmp_491_fu_13630_p4 = {{decipher_0_i32box_q58[31:24]}};

assign tmp_492_fu_13286_p4 = {{state_V_30_fu_13197_p2[55:48]}};

assign tmp_493_fu_13644_p4 = {{decipher_0_i32box_q57[15:8]}};

assign tmp_494_fu_13654_p4 = {{decipher_0_i32box_q57[23:16]}};

assign tmp_495_fu_13664_p4 = {{decipher_0_i32box_q57[31:24]}};

assign tmp_496_fu_13301_p4 = {{state_V_30_fu_13197_p2[63:56]}};

assign tmp_497_fu_13678_p4 = {{decipher_0_i32box_q56[15:8]}};

assign tmp_498_fu_13688_p4 = {{decipher_0_i32box_q56[23:16]}};

assign tmp_499_fu_13698_p4 = {{decipher_0_i32box_q56[31:24]}};

assign tmp_49_fu_5311_p4 = {{decipher_0_i32box_q170[23:16]}};

assign tmp_500_fu_13316_p4 = {{state_V_30_fu_13197_p2[71:64]}};

assign tmp_501_fu_13712_p4 = {{decipher_0_i32box_q55[15:8]}};

assign tmp_502_fu_13722_p4 = {{decipher_0_i32box_q55[23:16]}};

assign tmp_503_fu_13732_p4 = {{decipher_0_i32box_q55[31:24]}};

assign tmp_504_fu_13331_p4 = {{state_V_30_fu_13197_p2[79:72]}};

assign tmp_505_fu_13746_p4 = {{decipher_0_i32box_q54[15:8]}};

assign tmp_506_fu_13756_p4 = {{decipher_0_i32box_q54[23:16]}};

assign tmp_507_fu_13766_p4 = {{decipher_0_i32box_q54[31:24]}};

assign tmp_508_fu_13346_p4 = {{state_V_30_fu_13197_p2[87:80]}};

assign tmp_509_fu_13780_p4 = {{decipher_0_i32box_q53[15:8]}};

assign tmp_50_fu_5321_p4 = {{decipher_0_i32box_q170[31:24]}};

assign tmp_510_fu_13790_p4 = {{decipher_0_i32box_q53[23:16]}};

assign tmp_511_fu_13800_p4 = {{decipher_0_i32box_q53[31:24]}};

assign tmp_512_fu_13361_p4 = {{state_V_30_fu_13197_p2[95:88]}};

assign tmp_513_fu_13814_p4 = {{decipher_0_i32box_q52[15:8]}};

assign tmp_514_fu_13824_p4 = {{decipher_0_i32box_q52[23:16]}};

assign tmp_515_fu_13834_p4 = {{decipher_0_i32box_q52[31:24]}};

assign tmp_516_fu_13376_p4 = {{state_V_30_fu_13197_p2[103:96]}};

assign tmp_517_fu_13848_p4 = {{decipher_0_i32box_q51[15:8]}};

assign tmp_518_fu_13858_p4 = {{decipher_0_i32box_q51[23:16]}};

assign tmp_519_fu_13868_p4 = {{decipher_0_i32box_q51[31:24]}};

assign tmp_51_fu_4977_p4 = {{state_V_24_fu_4888_p2[55:48]}};

assign tmp_520_fu_13391_p4 = {{state_V_30_fu_13197_p2[111:104]}};

assign tmp_521_fu_13882_p4 = {{decipher_0_i32box_q50[15:8]}};

assign tmp_522_fu_13892_p4 = {{decipher_0_i32box_q50[23:16]}};

assign tmp_523_fu_13902_p4 = {{decipher_0_i32box_q50[31:24]}};

assign tmp_524_fu_13406_p4 = {{state_V_30_fu_13197_p2[119:112]}};

assign tmp_525_fu_13916_p4 = {{decipher_0_i32box_q49[15:8]}};

assign tmp_526_fu_13926_p4 = {{decipher_0_i32box_q49[23:16]}};

assign tmp_527_fu_13936_p4 = {{decipher_0_i32box_q49[31:24]}};

assign tmp_528_fu_13421_p4 = {{state_V_30_fu_13197_p2[127:120]}};

assign tmp_529_fu_13950_p4 = {{decipher_0_i32box_q48[15:8]}};

assign tmp_52_fu_5335_p4 = {{decipher_0_i32box_q169[15:8]}};

assign tmp_530_fu_13960_p4 = {{decipher_0_i32box_q48[23:16]}};

assign tmp_531_fu_13970_p4 = {{decipher_0_i32box_q48[31:24]}};

assign tmp_532_fu_14627_p4 = {{decipher_0_i32box_q47[15:8]}};

assign tmp_533_fu_14637_p4 = {{decipher_0_i32box_q47[23:16]}};

assign tmp_534_fu_14647_p4 = {{decipher_0_i32box_q47[31:24]}};

assign tmp_535_fu_14398_p4 = {{state_V_31_fu_14384_p2[15:8]}};

assign tmp_536_fu_14661_p4 = {{decipher_0_i32box_q46[15:8]}};

assign tmp_537_fu_14671_p4 = {{decipher_0_i32box_q46[23:16]}};

assign tmp_538_fu_14681_p4 = {{decipher_0_i32box_q46[31:24]}};

assign tmp_539_fu_14413_p4 = {{state_V_31_fu_14384_p2[23:16]}};

assign tmp_53_fu_5345_p4 = {{decipher_0_i32box_q169[23:16]}};

assign tmp_540_fu_14695_p4 = {{decipher_0_i32box_q45[15:8]}};

assign tmp_541_fu_14705_p4 = {{decipher_0_i32box_q45[23:16]}};

assign tmp_542_fu_14715_p4 = {{decipher_0_i32box_q45[31:24]}};

assign tmp_543_fu_14428_p4 = {{state_V_31_fu_14384_p2[31:24]}};

assign tmp_544_fu_14729_p4 = {{decipher_0_i32box_q44[15:8]}};

assign tmp_545_fu_14739_p4 = {{decipher_0_i32box_q44[23:16]}};

assign tmp_546_fu_14749_p4 = {{decipher_0_i32box_q44[31:24]}};

assign tmp_547_fu_14443_p4 = {{state_V_31_fu_14384_p2[39:32]}};

assign tmp_548_fu_14763_p4 = {{decipher_0_i32box_q43[15:8]}};

assign tmp_549_fu_14773_p4 = {{decipher_0_i32box_q43[23:16]}};

assign tmp_54_fu_5355_p4 = {{decipher_0_i32box_q169[31:24]}};

assign tmp_550_fu_14783_p4 = {{decipher_0_i32box_q43[31:24]}};

assign tmp_551_fu_14458_p4 = {{state_V_31_fu_14384_p2[47:40]}};

assign tmp_552_fu_14797_p4 = {{decipher_0_i32box_q42[15:8]}};

assign tmp_553_fu_14807_p4 = {{decipher_0_i32box_q42[23:16]}};

assign tmp_554_fu_14817_p4 = {{decipher_0_i32box_q42[31:24]}};

assign tmp_555_fu_14473_p4 = {{state_V_31_fu_14384_p2[55:48]}};

assign tmp_556_fu_14831_p4 = {{decipher_0_i32box_q41[15:8]}};

assign tmp_557_fu_14841_p4 = {{decipher_0_i32box_q41[23:16]}};

assign tmp_558_fu_14851_p4 = {{decipher_0_i32box_q41[31:24]}};

assign tmp_559_fu_14488_p4 = {{state_V_31_fu_14384_p2[63:56]}};

assign tmp_55_fu_4992_p4 = {{state_V_24_fu_4888_p2[63:56]}};

assign tmp_560_fu_14865_p4 = {{decipher_0_i32box_q40[15:8]}};

assign tmp_561_fu_14875_p4 = {{decipher_0_i32box_q40[23:16]}};

assign tmp_562_fu_14885_p4 = {{decipher_0_i32box_q40[31:24]}};

assign tmp_563_fu_14503_p4 = {{state_V_31_fu_14384_p2[71:64]}};

assign tmp_564_fu_14899_p4 = {{decipher_0_i32box_q39[15:8]}};

assign tmp_565_fu_14909_p4 = {{decipher_0_i32box_q39[23:16]}};

assign tmp_566_fu_14919_p4 = {{decipher_0_i32box_q39[31:24]}};

assign tmp_567_fu_14518_p4 = {{state_V_31_fu_14384_p2[79:72]}};

assign tmp_568_fu_14933_p4 = {{decipher_0_i32box_q38[15:8]}};

assign tmp_569_fu_14943_p4 = {{decipher_0_i32box_q38[23:16]}};

assign tmp_56_fu_5369_p4 = {{decipher_0_i32box_q168[15:8]}};

assign tmp_570_fu_14953_p4 = {{decipher_0_i32box_q38[31:24]}};

assign tmp_571_fu_14533_p4 = {{state_V_31_fu_14384_p2[87:80]}};

assign tmp_572_fu_14967_p4 = {{decipher_0_i32box_q37[15:8]}};

assign tmp_573_fu_14977_p4 = {{decipher_0_i32box_q37[23:16]}};

assign tmp_574_fu_14987_p4 = {{decipher_0_i32box_q37[31:24]}};

assign tmp_575_fu_14548_p4 = {{state_V_31_fu_14384_p2[95:88]}};

assign tmp_576_fu_15001_p4 = {{decipher_0_i32box_q36[15:8]}};

assign tmp_577_fu_15011_p4 = {{decipher_0_i32box_q36[23:16]}};

assign tmp_578_fu_15021_p4 = {{decipher_0_i32box_q36[31:24]}};

assign tmp_579_fu_14563_p4 = {{state_V_31_fu_14384_p2[103:96]}};

assign tmp_57_fu_5379_p4 = {{decipher_0_i32box_q168[23:16]}};

assign tmp_580_fu_15035_p4 = {{decipher_0_i32box_q35[15:8]}};

assign tmp_581_fu_15045_p4 = {{decipher_0_i32box_q35[23:16]}};

assign tmp_582_fu_15055_p4 = {{decipher_0_i32box_q35[31:24]}};

assign tmp_583_fu_14578_p4 = {{state_V_31_fu_14384_p2[111:104]}};

assign tmp_584_fu_15069_p4 = {{decipher_0_i32box_q34[15:8]}};

assign tmp_585_fu_15079_p4 = {{decipher_0_i32box_q34[23:16]}};

assign tmp_586_fu_15089_p4 = {{decipher_0_i32box_q34[31:24]}};

assign tmp_587_fu_14593_p4 = {{state_V_31_fu_14384_p2[119:112]}};

assign tmp_588_fu_15103_p4 = {{decipher_0_i32box_q33[15:8]}};

assign tmp_589_fu_15113_p4 = {{decipher_0_i32box_q33[23:16]}};

assign tmp_58_fu_5389_p4 = {{decipher_0_i32box_q168[31:24]}};

assign tmp_590_fu_15123_p4 = {{decipher_0_i32box_q33[31:24]}};

assign tmp_591_fu_14608_p4 = {{state_V_31_fu_14384_p2[127:120]}};

assign tmp_592_fu_15137_p4 = {{decipher_0_i32box_q32[15:8]}};

assign tmp_593_fu_15147_p4 = {{decipher_0_i32box_q32[23:16]}};

assign tmp_594_fu_15157_p4 = {{decipher_0_i32box_q32[31:24]}};

assign tmp_595_fu_15814_p4 = {{decipher_0_i32box_q31[15:8]}};

assign tmp_596_fu_15824_p4 = {{decipher_0_i32box_q31[23:16]}};

assign tmp_597_fu_15834_p4 = {{decipher_0_i32box_q31[31:24]}};

assign tmp_598_fu_15585_p4 = {{state_V_32_fu_15571_p2[15:8]}};

assign tmp_599_fu_15848_p4 = {{decipher_0_i32box_q30[15:8]}};

assign tmp_59_fu_5007_p4 = {{state_V_24_fu_4888_p2[71:64]}};

assign tmp_600_fu_15858_p4 = {{decipher_0_i32box_q30[23:16]}};

assign tmp_601_fu_15868_p4 = {{decipher_0_i32box_q30[31:24]}};

assign tmp_602_fu_15600_p4 = {{state_V_32_fu_15571_p2[23:16]}};

assign tmp_603_fu_15882_p4 = {{decipher_0_i32box_q29[15:8]}};

assign tmp_604_fu_15892_p4 = {{decipher_0_i32box_q29[23:16]}};

assign tmp_605_fu_15902_p4 = {{decipher_0_i32box_q29[31:24]}};

assign tmp_606_fu_15615_p4 = {{state_V_32_fu_15571_p2[31:24]}};

assign tmp_607_fu_15916_p4 = {{decipher_0_i32box_q28[15:8]}};

assign tmp_608_fu_15926_p4 = {{decipher_0_i32box_q28[23:16]}};

assign tmp_609_fu_15936_p4 = {{decipher_0_i32box_q28[31:24]}};

assign tmp_60_fu_5403_p4 = {{decipher_0_i32box_q167[15:8]}};

assign tmp_610_fu_15630_p4 = {{state_V_32_fu_15571_p2[39:32]}};

assign tmp_611_fu_15950_p4 = {{decipher_0_i32box_q27[15:8]}};

assign tmp_612_fu_15960_p4 = {{decipher_0_i32box_q27[23:16]}};

assign tmp_613_fu_15970_p4 = {{decipher_0_i32box_q27[31:24]}};

assign tmp_614_fu_15645_p4 = {{state_V_32_fu_15571_p2[47:40]}};

assign tmp_615_fu_15984_p4 = {{decipher_0_i32box_q26[15:8]}};

assign tmp_616_fu_15994_p4 = {{decipher_0_i32box_q26[23:16]}};

assign tmp_617_fu_16004_p4 = {{decipher_0_i32box_q26[31:24]}};

assign tmp_618_fu_15660_p4 = {{state_V_32_fu_15571_p2[55:48]}};

assign tmp_619_fu_16018_p4 = {{decipher_0_i32box_q25[15:8]}};

assign tmp_61_fu_5413_p4 = {{decipher_0_i32box_q167[23:16]}};

assign tmp_620_fu_16028_p4 = {{decipher_0_i32box_q25[23:16]}};

assign tmp_621_fu_16038_p4 = {{decipher_0_i32box_q25[31:24]}};

assign tmp_622_fu_15675_p4 = {{state_V_32_fu_15571_p2[63:56]}};

assign tmp_623_fu_16052_p4 = {{decipher_0_i32box_q24[15:8]}};

assign tmp_624_fu_16062_p4 = {{decipher_0_i32box_q24[23:16]}};

assign tmp_625_fu_16072_p4 = {{decipher_0_i32box_q24[31:24]}};

assign tmp_626_fu_15690_p4 = {{state_V_32_fu_15571_p2[71:64]}};

assign tmp_627_fu_16086_p4 = {{decipher_0_i32box_q23[15:8]}};

assign tmp_628_fu_16096_p4 = {{decipher_0_i32box_q23[23:16]}};

assign tmp_629_fu_16106_p4 = {{decipher_0_i32box_q23[31:24]}};

assign tmp_62_fu_5423_p4 = {{decipher_0_i32box_q167[31:24]}};

assign tmp_630_fu_15705_p4 = {{state_V_32_fu_15571_p2[79:72]}};

assign tmp_631_fu_16120_p4 = {{decipher_0_i32box_q22[15:8]}};

assign tmp_632_fu_16130_p4 = {{decipher_0_i32box_q22[23:16]}};

assign tmp_633_fu_16140_p4 = {{decipher_0_i32box_q22[31:24]}};

assign tmp_634_fu_15720_p4 = {{state_V_32_fu_15571_p2[87:80]}};

assign tmp_635_fu_16154_p4 = {{decipher_0_i32box_q21[15:8]}};

assign tmp_636_fu_16164_p4 = {{decipher_0_i32box_q21[23:16]}};

assign tmp_637_fu_16174_p4 = {{decipher_0_i32box_q21[31:24]}};

assign tmp_638_fu_15735_p4 = {{state_V_32_fu_15571_p2[95:88]}};

assign tmp_639_fu_16188_p4 = {{decipher_0_i32box_q20[15:8]}};

assign tmp_63_fu_5022_p4 = {{state_V_24_fu_4888_p2[79:72]}};

assign tmp_640_fu_16198_p4 = {{decipher_0_i32box_q20[23:16]}};

assign tmp_641_fu_16208_p4 = {{decipher_0_i32box_q20[31:24]}};

assign tmp_642_fu_15750_p4 = {{state_V_32_fu_15571_p2[103:96]}};

assign tmp_643_fu_16222_p4 = {{decipher_0_i32box_q19[15:8]}};

assign tmp_644_fu_16232_p4 = {{decipher_0_i32box_q19[23:16]}};

assign tmp_645_fu_16242_p4 = {{decipher_0_i32box_q19[31:24]}};

assign tmp_646_fu_15765_p4 = {{state_V_32_fu_15571_p2[111:104]}};

assign tmp_647_fu_16256_p4 = {{decipher_0_i32box_q18[15:8]}};

assign tmp_648_fu_16266_p4 = {{decipher_0_i32box_q18[23:16]}};

assign tmp_649_fu_16276_p4 = {{decipher_0_i32box_q18[31:24]}};

assign tmp_64_fu_5437_p4 = {{decipher_0_i32box_q166[15:8]}};

assign tmp_650_fu_15780_p4 = {{state_V_32_fu_15571_p2[119:112]}};

assign tmp_651_fu_16290_p4 = {{decipher_0_i32box_q17[15:8]}};

assign tmp_652_fu_16300_p4 = {{decipher_0_i32box_q17[23:16]}};

assign tmp_653_fu_16310_p4 = {{decipher_0_i32box_q17[31:24]}};

assign tmp_654_fu_15795_p4 = {{state_V_32_fu_15571_p2[127:120]}};

assign tmp_655_fu_16324_p4 = {{decipher_0_i32box_q16[15:8]}};

assign tmp_656_fu_16334_p4 = {{decipher_0_i32box_q16[23:16]}};

assign tmp_657_fu_16344_p4 = {{decipher_0_i32box_q16[31:24]}};

assign tmp_658_fu_17001_p4 = {{decipher_0_i32box_q15[15:8]}};

assign tmp_659_fu_17011_p4 = {{decipher_0_i32box_q15[23:16]}};

assign tmp_65_fu_5447_p4 = {{decipher_0_i32box_q166[23:16]}};

assign tmp_660_fu_17021_p4 = {{decipher_0_i32box_q15[31:24]}};

assign tmp_661_fu_16772_p4 = {{state_V_33_fu_16758_p2[15:8]}};

assign tmp_662_fu_17035_p4 = {{decipher_0_i32box_q14[15:8]}};

assign tmp_663_fu_17045_p4 = {{decipher_0_i32box_q14[23:16]}};

assign tmp_664_fu_17055_p4 = {{decipher_0_i32box_q14[31:24]}};

assign tmp_665_fu_16787_p4 = {{state_V_33_fu_16758_p2[23:16]}};

assign tmp_666_fu_17069_p4 = {{decipher_0_i32box_q13[15:8]}};

assign tmp_667_fu_17079_p4 = {{decipher_0_i32box_q13[23:16]}};

assign tmp_668_fu_17089_p4 = {{decipher_0_i32box_q13[31:24]}};

assign tmp_669_fu_16802_p4 = {{state_V_33_fu_16758_p2[31:24]}};

assign tmp_66_fu_5457_p4 = {{decipher_0_i32box_q166[31:24]}};

assign tmp_670_fu_17103_p4 = {{decipher_0_i32box_q12[15:8]}};

assign tmp_671_fu_17113_p4 = {{decipher_0_i32box_q12[23:16]}};

assign tmp_672_fu_17123_p4 = {{decipher_0_i32box_q12[31:24]}};

assign tmp_673_fu_16817_p4 = {{state_V_33_fu_16758_p2[39:32]}};

assign tmp_674_fu_17137_p4 = {{decipher_0_i32box_q11[15:8]}};

assign tmp_675_fu_17147_p4 = {{decipher_0_i32box_q11[23:16]}};

assign tmp_676_fu_17157_p4 = {{decipher_0_i32box_q11[31:24]}};

assign tmp_677_fu_16832_p4 = {{state_V_33_fu_16758_p2[47:40]}};

assign tmp_678_fu_17171_p4 = {{decipher_0_i32box_q10[15:8]}};

assign tmp_679_fu_17181_p4 = {{decipher_0_i32box_q10[23:16]}};

assign tmp_67_fu_5037_p4 = {{state_V_24_fu_4888_p2[87:80]}};

assign tmp_680_fu_17191_p4 = {{decipher_0_i32box_q10[31:24]}};

assign tmp_681_fu_16847_p4 = {{state_V_33_fu_16758_p2[55:48]}};

assign tmp_682_fu_17205_p4 = {{decipher_0_i32box_q9[15:8]}};

assign tmp_683_fu_17215_p4 = {{decipher_0_i32box_q9[23:16]}};

assign tmp_684_fu_17225_p4 = {{decipher_0_i32box_q9[31:24]}};

assign tmp_685_fu_16862_p4 = {{state_V_33_fu_16758_p2[63:56]}};

assign tmp_686_fu_17239_p4 = {{decipher_0_i32box_q8[15:8]}};

assign tmp_687_fu_17249_p4 = {{decipher_0_i32box_q8[23:16]}};

assign tmp_688_fu_17259_p4 = {{decipher_0_i32box_q8[31:24]}};

assign tmp_689_fu_16877_p4 = {{state_V_33_fu_16758_p2[71:64]}};

assign tmp_68_fu_5471_p4 = {{decipher_0_i32box_q165[15:8]}};

assign tmp_690_fu_17273_p4 = {{decipher_0_i32box_q7[15:8]}};

assign tmp_691_fu_17283_p4 = {{decipher_0_i32box_q7[23:16]}};

assign tmp_692_fu_17293_p4 = {{decipher_0_i32box_q7[31:24]}};

assign tmp_693_fu_16892_p4 = {{state_V_33_fu_16758_p2[79:72]}};

assign tmp_694_fu_17307_p4 = {{decipher_0_i32box_q6[15:8]}};

assign tmp_695_fu_17317_p4 = {{decipher_0_i32box_q6[23:16]}};

assign tmp_696_fu_17327_p4 = {{decipher_0_i32box_q6[31:24]}};

assign tmp_697_fu_16907_p4 = {{state_V_33_fu_16758_p2[87:80]}};

assign tmp_698_fu_17341_p4 = {{decipher_0_i32box_q5[15:8]}};

assign tmp_699_fu_17351_p4 = {{decipher_0_i32box_q5[23:16]}};

assign tmp_69_fu_5481_p4 = {{decipher_0_i32box_q165[23:16]}};

assign tmp_700_fu_17361_p4 = {{decipher_0_i32box_q5[31:24]}};

assign tmp_701_fu_16922_p4 = {{state_V_33_fu_16758_p2[95:88]}};

assign tmp_702_fu_17375_p4 = {{decipher_0_i32box_q4[15:8]}};

assign tmp_703_fu_17385_p4 = {{decipher_0_i32box_q4[23:16]}};

assign tmp_704_fu_17395_p4 = {{decipher_0_i32box_q4[31:24]}};

assign tmp_705_fu_16937_p4 = {{state_V_33_fu_16758_p2[103:96]}};

assign tmp_706_fu_17409_p4 = {{decipher_0_i32box_q3[15:8]}};

assign tmp_707_fu_17419_p4 = {{decipher_0_i32box_q3[23:16]}};

assign tmp_708_fu_17429_p4 = {{decipher_0_i32box_q3[31:24]}};

assign tmp_709_fu_16952_p4 = {{state_V_33_fu_16758_p2[111:104]}};

assign tmp_70_fu_5491_p4 = {{decipher_0_i32box_q165[31:24]}};

assign tmp_710_fu_17443_p4 = {{decipher_0_i32box_q2[15:8]}};

assign tmp_711_fu_17453_p4 = {{decipher_0_i32box_q2[23:16]}};

assign tmp_712_fu_17463_p4 = {{decipher_0_i32box_q2[31:24]}};

assign tmp_713_fu_16967_p4 = {{state_V_33_fu_16758_p2[119:112]}};

assign tmp_714_fu_17477_p4 = {{decipher_0_i32box_q1[15:8]}};

assign tmp_715_fu_17487_p4 = {{decipher_0_i32box_q1[23:16]}};

assign tmp_716_fu_17497_p4 = {{decipher_0_i32box_q1[31:24]}};

assign tmp_717_fu_16982_p4 = {{state_V_33_fu_16758_p2[127:120]}};

assign tmp_718_fu_17511_p4 = {{decipher_0_i32box_q0[15:8]}};

assign tmp_719_fu_17521_p4 = {{decipher_0_i32box_q0[23:16]}};

assign tmp_71_fu_5052_p4 = {{state_V_24_fu_4888_p2[95:88]}};

assign tmp_720_fu_17531_p4 = {{decipher_0_i32box_q0[31:24]}};

assign tmp_72_fu_5505_p4 = {{decipher_0_i32box_q164[15:8]}};

assign tmp_73_fu_5515_p4 = {{decipher_0_i32box_q164[23:16]}};

assign tmp_74_fu_5525_p4 = {{decipher_0_i32box_q164[31:24]}};

assign tmp_75_fu_5067_p4 = {{state_V_24_fu_4888_p2[103:96]}};

assign tmp_76_fu_5539_p4 = {{decipher_0_i32box_q163[15:8]}};

assign tmp_77_fu_5549_p4 = {{decipher_0_i32box_q163[23:16]}};

assign tmp_78_fu_5559_p4 = {{decipher_0_i32box_q163[31:24]}};

assign tmp_79_fu_5082_p4 = {{state_V_24_fu_4888_p2[111:104]}};

assign tmp_80_fu_5573_p4 = {{decipher_0_i32box_q162[15:8]}};

assign tmp_81_fu_5583_p4 = {{decipher_0_i32box_q162[23:16]}};

assign tmp_82_fu_5593_p4 = {{decipher_0_i32box_q162[31:24]}};

assign tmp_83_fu_5097_p4 = {{state_V_24_fu_4888_p2[119:112]}};

assign tmp_84_fu_5607_p4 = {{decipher_0_i32box_q161[15:8]}};

assign tmp_85_fu_5617_p4 = {{decipher_0_i32box_q161[23:16]}};

assign tmp_86_fu_5627_p4 = {{decipher_0_i32box_q161[31:24]}};

assign tmp_87_fu_5112_p4 = {{state_V_24_fu_4888_p2[127:120]}};

assign tmp_88_fu_5641_p4 = {{decipher_0_i32box_q160[15:8]}};

assign tmp_89_fu_5651_p4 = {{decipher_0_i32box_q160[23:16]}};

assign tmp_90_fu_5661_p4 = {{decipher_0_i32box_q160[31:24]}};

assign tmp_91_fu_6318_p4 = {{decipher_0_i32box_q159[15:8]}};

assign tmp_92_fu_6328_p4 = {{decipher_0_i32box_q159[23:16]}};

assign tmp_93_fu_6338_p4 = {{decipher_0_i32box_q159[31:24]}};

assign tmp_94_fu_6089_p4 = {{state_V_25_fu_6075_p2[15:8]}};

assign tmp_95_fu_6352_p4 = {{decipher_0_i32box_q158[15:8]}};

assign tmp_96_fu_6362_p4 = {{decipher_0_i32box_q158[23:16]}};

assign tmp_97_fu_6372_p4 = {{decipher_0_i32box_q158[31:24]}};

assign tmp_98_fu_6104_p4 = {{state_V_25_fu_6075_p2[23:16]}};

assign tmp_99_fu_6386_p4 = {{decipher_0_i32box_q157[15:8]}};

assign tmp_s_fu_4627_p4 = {{ret_V_fu_4612_p2[111:104]}};

assign trunc_ln674_100_fu_12351_p1 = decipher_0_i32box_q76[7:0];

assign trunc_ln674_101_fu_12385_p1 = decipher_0_i32box_q75[7:0];

assign trunc_ln674_102_fu_12419_p1 = decipher_0_i32box_q74[7:0];

assign trunc_ln674_103_fu_12453_p1 = decipher_0_i32box_q73[7:0];

assign trunc_ln674_104_fu_12487_p1 = decipher_0_i32box_q72[7:0];

assign trunc_ln674_105_fu_12521_p1 = decipher_0_i32box_q71[7:0];

assign trunc_ln674_106_fu_12555_p1 = decipher_0_i32box_q70[7:0];

assign trunc_ln674_107_fu_12589_p1 = decipher_0_i32box_q69[7:0];

assign trunc_ln674_108_fu_12623_p1 = decipher_0_i32box_q68[7:0];

assign trunc_ln674_109_fu_12657_p1 = decipher_0_i32box_q67[7:0];

assign trunc_ln674_10_fu_5433_p1 = decipher_0_i32box_q166[7:0];

assign trunc_ln674_110_fu_12691_p1 = decipher_0_i32box_q66[7:0];

assign trunc_ln674_111_fu_12725_p1 = decipher_0_i32box_q65[7:0];

assign trunc_ln674_112_fu_12759_p1 = decipher_0_i32box_q64[7:0];

assign trunc_ln674_113_fu_13436_p1 = decipher_0_i32box_q63[7:0];

assign trunc_ln674_114_fu_13470_p1 = decipher_0_i32box_q62[7:0];

assign trunc_ln674_115_fu_13504_p1 = decipher_0_i32box_q61[7:0];

assign trunc_ln674_116_fu_13538_p1 = decipher_0_i32box_q60[7:0];

assign trunc_ln674_117_fu_13572_p1 = decipher_0_i32box_q59[7:0];

assign trunc_ln674_118_fu_13606_p1 = decipher_0_i32box_q58[7:0];

assign trunc_ln674_119_fu_13640_p1 = decipher_0_i32box_q57[7:0];

assign trunc_ln674_11_fu_5467_p1 = decipher_0_i32box_q165[7:0];

assign trunc_ln674_120_fu_13674_p1 = decipher_0_i32box_q56[7:0];

assign trunc_ln674_121_fu_13708_p1 = decipher_0_i32box_q55[7:0];

assign trunc_ln674_122_fu_13742_p1 = decipher_0_i32box_q54[7:0];

assign trunc_ln674_123_fu_13776_p1 = decipher_0_i32box_q53[7:0];

assign trunc_ln674_124_fu_13810_p1 = decipher_0_i32box_q52[7:0];

assign trunc_ln674_125_fu_13844_p1 = decipher_0_i32box_q51[7:0];

assign trunc_ln674_126_fu_13878_p1 = decipher_0_i32box_q50[7:0];

assign trunc_ln674_127_fu_13912_p1 = decipher_0_i32box_q49[7:0];

assign trunc_ln674_128_fu_13946_p1 = decipher_0_i32box_q48[7:0];

assign trunc_ln674_129_fu_14623_p1 = decipher_0_i32box_q47[7:0];

assign trunc_ln674_12_fu_5501_p1 = decipher_0_i32box_q164[7:0];

assign trunc_ln674_130_fu_14657_p1 = decipher_0_i32box_q46[7:0];

assign trunc_ln674_131_fu_14691_p1 = decipher_0_i32box_q45[7:0];

assign trunc_ln674_132_fu_14725_p1 = decipher_0_i32box_q44[7:0];

assign trunc_ln674_133_fu_14759_p1 = decipher_0_i32box_q43[7:0];

assign trunc_ln674_134_fu_14793_p1 = decipher_0_i32box_q42[7:0];

assign trunc_ln674_135_fu_14827_p1 = decipher_0_i32box_q41[7:0];

assign trunc_ln674_136_fu_14861_p1 = decipher_0_i32box_q40[7:0];

assign trunc_ln674_137_fu_14895_p1 = decipher_0_i32box_q39[7:0];

assign trunc_ln674_138_fu_14929_p1 = decipher_0_i32box_q38[7:0];

assign trunc_ln674_139_fu_14963_p1 = decipher_0_i32box_q37[7:0];

assign trunc_ln674_13_fu_5535_p1 = decipher_0_i32box_q163[7:0];

assign trunc_ln674_140_fu_14997_p1 = decipher_0_i32box_q36[7:0];

assign trunc_ln674_141_fu_15031_p1 = decipher_0_i32box_q35[7:0];

assign trunc_ln674_142_fu_15065_p1 = decipher_0_i32box_q34[7:0];

assign trunc_ln674_143_fu_15099_p1 = decipher_0_i32box_q33[7:0];

assign trunc_ln674_144_fu_15133_p1 = decipher_0_i32box_q32[7:0];

assign trunc_ln674_145_fu_15810_p1 = decipher_0_i32box_q31[7:0];

assign trunc_ln674_146_fu_15844_p1 = decipher_0_i32box_q30[7:0];

assign trunc_ln674_147_fu_15878_p1 = decipher_0_i32box_q29[7:0];

assign trunc_ln674_148_fu_15912_p1 = decipher_0_i32box_q28[7:0];

assign trunc_ln674_149_fu_15946_p1 = decipher_0_i32box_q27[7:0];

assign trunc_ln674_14_fu_5569_p1 = decipher_0_i32box_q162[7:0];

assign trunc_ln674_150_fu_15980_p1 = decipher_0_i32box_q26[7:0];

assign trunc_ln674_151_fu_16014_p1 = decipher_0_i32box_q25[7:0];

assign trunc_ln674_152_fu_16048_p1 = decipher_0_i32box_q24[7:0];

assign trunc_ln674_153_fu_16082_p1 = decipher_0_i32box_q23[7:0];

assign trunc_ln674_154_fu_16116_p1 = decipher_0_i32box_q22[7:0];

assign trunc_ln674_155_fu_16150_p1 = decipher_0_i32box_q21[7:0];

assign trunc_ln674_156_fu_16184_p1 = decipher_0_i32box_q20[7:0];

assign trunc_ln674_157_fu_16218_p1 = decipher_0_i32box_q19[7:0];

assign trunc_ln674_158_fu_16252_p1 = decipher_0_i32box_q18[7:0];

assign trunc_ln674_159_fu_16286_p1 = decipher_0_i32box_q17[7:0];

assign trunc_ln674_15_fu_5603_p1 = decipher_0_i32box_q161[7:0];

assign trunc_ln674_160_fu_16320_p1 = decipher_0_i32box_q16[7:0];

assign trunc_ln674_161_fu_16997_p1 = decipher_0_i32box_q15[7:0];

assign trunc_ln674_162_fu_17031_p1 = decipher_0_i32box_q14[7:0];

assign trunc_ln674_163_fu_17065_p1 = decipher_0_i32box_q13[7:0];

assign trunc_ln674_164_fu_17099_p1 = decipher_0_i32box_q12[7:0];

assign trunc_ln674_165_fu_17133_p1 = decipher_0_i32box_q11[7:0];

assign trunc_ln674_166_fu_17167_p1 = decipher_0_i32box_q10[7:0];

assign trunc_ln674_167_fu_17201_p1 = decipher_0_i32box_q9[7:0];

assign trunc_ln674_168_fu_17235_p1 = decipher_0_i32box_q8[7:0];

assign trunc_ln674_169_fu_17269_p1 = decipher_0_i32box_q7[7:0];

assign trunc_ln674_16_fu_5637_p1 = decipher_0_i32box_q160[7:0];

assign trunc_ln674_170_fu_17303_p1 = decipher_0_i32box_q6[7:0];

assign trunc_ln674_171_fu_17337_p1 = decipher_0_i32box_q5[7:0];

assign trunc_ln674_172_fu_17371_p1 = decipher_0_i32box_q4[7:0];

assign trunc_ln674_173_fu_17405_p1 = decipher_0_i32box_q3[7:0];

assign trunc_ln674_174_fu_17439_p1 = decipher_0_i32box_q2[7:0];

assign trunc_ln674_175_fu_17473_p1 = decipher_0_i32box_q1[7:0];

assign trunc_ln674_176_fu_17507_p1 = decipher_0_i32box_q0[7:0];

assign trunc_ln674_17_fu_6314_p1 = decipher_0_i32box_q159[7:0];

assign trunc_ln674_18_fu_6348_p1 = decipher_0_i32box_q158[7:0];

assign trunc_ln674_19_fu_6382_p1 = decipher_0_i32box_q157[7:0];

assign trunc_ln674_20_fu_6416_p1 = decipher_0_i32box_q156[7:0];

assign trunc_ln674_21_fu_6450_p1 = decipher_0_i32box_q155[7:0];

assign trunc_ln674_22_fu_6484_p1 = decipher_0_i32box_q154[7:0];

assign trunc_ln674_23_fu_6518_p1 = decipher_0_i32box_q153[7:0];

assign trunc_ln674_24_fu_6552_p1 = decipher_0_i32box_q152[7:0];

assign trunc_ln674_25_fu_6586_p1 = decipher_0_i32box_q151[7:0];

assign trunc_ln674_26_fu_6620_p1 = decipher_0_i32box_q150[7:0];

assign trunc_ln674_27_fu_6654_p1 = decipher_0_i32box_q149[7:0];

assign trunc_ln674_28_fu_6688_p1 = decipher_0_i32box_q148[7:0];

assign trunc_ln674_29_fu_6722_p1 = decipher_0_i32box_q147[7:0];

assign trunc_ln674_2_fu_5161_p1 = decipher_0_i32box_q174[7:0];

assign trunc_ln674_30_fu_6756_p1 = decipher_0_i32box_q146[7:0];

assign trunc_ln674_31_fu_6790_p1 = decipher_0_i32box_q145[7:0];

assign trunc_ln674_32_fu_6824_p1 = decipher_0_i32box_q144[7:0];

assign trunc_ln674_33_fu_7501_p1 = decipher_0_i32box_q143[7:0];

assign trunc_ln674_34_fu_7535_p1 = decipher_0_i32box_q142[7:0];

assign trunc_ln674_35_fu_7569_p1 = decipher_0_i32box_q141[7:0];

assign trunc_ln674_36_fu_7603_p1 = decipher_0_i32box_q140[7:0];

assign trunc_ln674_37_fu_7637_p1 = decipher_0_i32box_q139[7:0];

assign trunc_ln674_38_fu_7671_p1 = decipher_0_i32box_q138[7:0];

assign trunc_ln674_39_fu_7705_p1 = decipher_0_i32box_q137[7:0];

assign trunc_ln674_3_fu_5195_p1 = decipher_0_i32box_q173[7:0];

assign trunc_ln674_40_fu_7739_p1 = decipher_0_i32box_q136[7:0];

assign trunc_ln674_41_fu_7773_p1 = decipher_0_i32box_q135[7:0];

assign trunc_ln674_42_fu_7807_p1 = decipher_0_i32box_q134[7:0];

assign trunc_ln674_43_fu_7841_p1 = decipher_0_i32box_q133[7:0];

assign trunc_ln674_44_fu_7875_p1 = decipher_0_i32box_q132[7:0];

assign trunc_ln674_45_fu_7909_p1 = decipher_0_i32box_q131[7:0];

assign trunc_ln674_46_fu_7943_p1 = decipher_0_i32box_q130[7:0];

assign trunc_ln674_47_fu_7977_p1 = decipher_0_i32box_q129[7:0];

assign trunc_ln674_48_fu_8011_p1 = decipher_0_i32box_q128[7:0];

assign trunc_ln674_49_fu_8688_p1 = decipher_0_i32box_q127[7:0];

assign trunc_ln674_4_fu_5229_p1 = decipher_0_i32box_q172[7:0];

assign trunc_ln674_50_fu_8722_p1 = decipher_0_i32box_q126[7:0];

assign trunc_ln674_51_fu_8756_p1 = decipher_0_i32box_q125[7:0];

assign trunc_ln674_52_fu_8790_p1 = decipher_0_i32box_q124[7:0];

assign trunc_ln674_53_fu_8824_p1 = decipher_0_i32box_q123[7:0];

assign trunc_ln674_54_fu_8858_p1 = decipher_0_i32box_q122[7:0];

assign trunc_ln674_55_fu_8892_p1 = decipher_0_i32box_q121[7:0];

assign trunc_ln674_56_fu_8926_p1 = decipher_0_i32box_q120[7:0];

assign trunc_ln674_57_fu_8960_p1 = decipher_0_i32box_q119[7:0];

assign trunc_ln674_58_fu_8994_p1 = decipher_0_i32box_q118[7:0];

assign trunc_ln674_59_fu_9028_p1 = decipher_0_i32box_q117[7:0];

assign trunc_ln674_5_fu_5263_p1 = decipher_0_i32box_q171[7:0];

assign trunc_ln674_60_fu_9062_p1 = decipher_0_i32box_q116[7:0];

assign trunc_ln674_61_fu_9096_p1 = decipher_0_i32box_q115[7:0];

assign trunc_ln674_62_fu_9130_p1 = decipher_0_i32box_q114[7:0];

assign trunc_ln674_63_fu_9164_p1 = decipher_0_i32box_q113[7:0];

assign trunc_ln674_64_fu_9198_p1 = decipher_0_i32box_q112[7:0];

assign trunc_ln674_65_fu_9875_p1 = decipher_0_i32box_q111[7:0];

assign trunc_ln674_66_fu_9909_p1 = decipher_0_i32box_q110[7:0];

assign trunc_ln674_67_fu_9943_p1 = decipher_0_i32box_q109[7:0];

assign trunc_ln674_68_fu_9977_p1 = decipher_0_i32box_q108[7:0];

assign trunc_ln674_69_fu_10011_p1 = decipher_0_i32box_q107[7:0];

assign trunc_ln674_6_fu_5297_p1 = decipher_0_i32box_q170[7:0];

assign trunc_ln674_70_fu_10045_p1 = decipher_0_i32box_q106[7:0];

assign trunc_ln674_71_fu_10079_p1 = decipher_0_i32box_q105[7:0];

assign trunc_ln674_72_fu_10113_p1 = decipher_0_i32box_q104[7:0];

assign trunc_ln674_73_fu_10147_p1 = decipher_0_i32box_q103[7:0];

assign trunc_ln674_74_fu_10181_p1 = decipher_0_i32box_q102[7:0];

assign trunc_ln674_75_fu_10215_p1 = decipher_0_i32box_q101[7:0];

assign trunc_ln674_76_fu_10249_p1 = decipher_0_i32box_q100[7:0];

assign trunc_ln674_77_fu_10283_p1 = decipher_0_i32box_q99[7:0];

assign trunc_ln674_78_fu_10317_p1 = decipher_0_i32box_q98[7:0];

assign trunc_ln674_79_fu_10351_p1 = decipher_0_i32box_q97[7:0];

assign trunc_ln674_7_fu_5331_p1 = decipher_0_i32box_q169[7:0];

assign trunc_ln674_80_fu_10385_p1 = decipher_0_i32box_q96[7:0];

assign trunc_ln674_81_fu_11062_p1 = decipher_0_i32box_q95[7:0];

assign trunc_ln674_82_fu_11096_p1 = decipher_0_i32box_q94[7:0];

assign trunc_ln674_83_fu_11130_p1 = decipher_0_i32box_q93[7:0];

assign trunc_ln674_84_fu_11164_p1 = decipher_0_i32box_q92[7:0];

assign trunc_ln674_85_fu_11198_p1 = decipher_0_i32box_q91[7:0];

assign trunc_ln674_86_fu_11232_p1 = decipher_0_i32box_q90[7:0];

assign trunc_ln674_87_fu_11266_p1 = decipher_0_i32box_q89[7:0];

assign trunc_ln674_88_fu_11300_p1 = decipher_0_i32box_q88[7:0];

assign trunc_ln674_89_fu_11334_p1 = decipher_0_i32box_q87[7:0];

assign trunc_ln674_8_fu_5365_p1 = decipher_0_i32box_q168[7:0];

assign trunc_ln674_90_fu_11368_p1 = decipher_0_i32box_q86[7:0];

assign trunc_ln674_91_fu_11402_p1 = decipher_0_i32box_q85[7:0];

assign trunc_ln674_92_fu_11436_p1 = decipher_0_i32box_q84[7:0];

assign trunc_ln674_93_fu_11470_p1 = decipher_0_i32box_q83[7:0];

assign trunc_ln674_94_fu_11504_p1 = decipher_0_i32box_q82[7:0];

assign trunc_ln674_95_fu_11538_p1 = decipher_0_i32box_q81[7:0];

assign trunc_ln674_96_fu_11572_p1 = decipher_0_i32box_q80[7:0];

assign trunc_ln674_97_fu_12249_p1 = decipher_0_i32box_q79[7:0];

assign trunc_ln674_98_fu_12283_p1 = decipher_0_i32box_q78[7:0];

assign trunc_ln674_99_fu_12317_p1 = decipher_0_i32box_q77[7:0];

assign trunc_ln674_9_fu_5399_p1 = decipher_0_i32box_q167[7:0];

assign trunc_ln674_fu_5127_p1 = decipher_0_i32box_q175[7:0];

assign trunc_ln708_10_fu_15576_p1 = state_V_32_fu_15571_p2[7:0];

assign trunc_ln708_11_fu_16763_p1 = state_V_33_fu_16758_p2[7:0];

assign trunc_ln708_1_fu_4893_p1 = state_V_24_fu_4888_p2[7:0];

assign trunc_ln708_2_fu_6080_p1 = state_V_25_fu_6075_p2[7:0];

assign trunc_ln708_3_fu_7267_p1 = state_V_26_fu_7262_p2[7:0];

assign trunc_ln708_4_fu_8454_p1 = state_V_27_fu_8449_p2[7:0];

assign trunc_ln708_5_fu_9641_p1 = state_V_28_fu_9636_p2[7:0];

assign trunc_ln708_6_fu_10828_p1 = state_V_29_fu_10823_p2[7:0];

assign trunc_ln708_7_fu_12015_p1 = state_V_fu_12010_p2[7:0];

assign trunc_ln708_8_fu_13202_p1 = state_V_30_fu_13197_p2[7:0];

assign trunc_ln708_9_fu_14389_p1 = state_V_31_fu_14384_p2[7:0];

assign trunc_ln708_fu_4618_p1 = ret_V_fu_4612_p2[7:0];

assign xor_ln1545_100_fu_7140_p2 = (xor_ln1545_99_fu_7128_p2 ^ xor_ln1545_101_fu_7134_p2);

assign xor_ln1545_101_fu_7134_p2 = (trunc_ln674_31_fu_6790_p1 ^ tmp_153_fu_6848_p4);

assign xor_ln1545_102_fu_8045_p2 = (tmp_158_fu_7539_p4 ^ tmp_156_fu_7525_p4);

assign xor_ln1545_103_fu_8057_p2 = (xor_ln1545_104_fu_8051_p2 ^ xor_ln1545_102_fu_8045_p2);

assign xor_ln1545_104_fu_8051_p2 = (trunc_ln674_36_fu_7603_p1 ^ tmp_163_fu_7583_p4);

assign xor_ln1545_105_fu_8063_p2 = (trunc_ln674_33_fu_7501_p1 ^ tmp_160_fu_7559_p4);

assign xor_ln1545_106_fu_8075_p2 = (xor_ln1545_107_fu_8069_p2 ^ xor_ln1545_105_fu_8063_p2);

assign xor_ln1545_107_fu_8069_p2 = (tmp_167_fu_7617_p4 ^ tmp_162_fu_7573_p4);

assign xor_ln1545_108_fu_8081_p2 = (trunc_ln674_34_fu_7535_p1 ^ tmp_155_fu_7515_p4);

assign xor_ln1545_109_fu_8093_p2 = (xor_ln1545_110_fu_8087_p2 ^ xor_ln1545_108_fu_8081_p2);

assign xor_ln1545_10_fu_5701_p2 = (xor_ln1545_9_fu_5689_p2 ^ xor_ln1545_11_fu_5695_p2);

assign xor_ln1545_110_fu_8087_p2 = (tmp_166_fu_7607_p4 ^ tmp_164_fu_7593_p4);

assign xor_ln1545_111_fu_8099_p2 = (tmp_159_fu_7549_p4 ^ tmp_154_fu_7505_p4);

assign xor_ln1545_112_fu_8105_p2 = (trunc_ln674_35_fu_7569_p1 ^ tmp_168_fu_7627_p4);

assign xor_ln1545_114_fu_8117_p2 = (tmp_174_fu_7675_p4 ^ tmp_172_fu_7661_p4);

assign xor_ln1545_115_fu_8129_p2 = (xor_ln1545_116_fu_8123_p2 ^ xor_ln1545_114_fu_8117_p2);

assign xor_ln1545_116_fu_8123_p2 = (trunc_ln674_40_fu_7739_p1 ^ tmp_179_fu_7719_p4);

assign xor_ln1545_117_fu_8135_p2 = (trunc_ln674_37_fu_7637_p1 ^ tmp_176_fu_7695_p4);

assign xor_ln1545_118_fu_8147_p2 = (xor_ln1545_119_fu_8141_p2 ^ xor_ln1545_117_fu_8135_p2);

assign xor_ln1545_119_fu_8141_p2 = (tmp_183_fu_7753_p4 ^ tmp_178_fu_7709_p4);

assign xor_ln1545_11_fu_5695_p2 = (tmp_41_fu_5243_p4 ^ tmp_36_fu_5199_p4);

assign xor_ln1545_120_fu_8153_p2 = (trunc_ln674_38_fu_7671_p1 ^ tmp_171_fu_7651_p4);

assign xor_ln1545_121_fu_8165_p2 = (xor_ln1545_122_fu_8159_p2 ^ xor_ln1545_120_fu_8153_p2);

assign xor_ln1545_122_fu_8159_p2 = (tmp_182_fu_7743_p4 ^ tmp_180_fu_7729_p4);

assign xor_ln1545_123_fu_8171_p2 = (tmp_175_fu_7685_p4 ^ tmp_170_fu_7641_p4);

assign xor_ln1545_124_fu_8183_p2 = (xor_ln1545_125_fu_8177_p2 ^ xor_ln1545_123_fu_8171_p2);

assign xor_ln1545_125_fu_8177_p2 = (trunc_ln674_39_fu_7705_p1 ^ tmp_184_fu_7763_p4);

assign xor_ln1545_126_fu_8189_p2 = (tmp_190_fu_7811_p4 ^ tmp_188_fu_7797_p4);

assign xor_ln1545_127_fu_8201_p2 = (xor_ln1545_128_fu_8195_p2 ^ xor_ln1545_126_fu_8189_p2);

assign xor_ln1545_128_fu_8195_p2 = (trunc_ln674_44_fu_7875_p1 ^ tmp_195_fu_7855_p4);

assign xor_ln1545_129_fu_8207_p2 = (trunc_ln674_41_fu_7773_p1 ^ tmp_192_fu_7831_p4);

assign xor_ln1545_12_fu_5707_p2 = (trunc_ln674_2_fu_5161_p1 ^ tmp_29_fu_5141_p4);

assign xor_ln1545_130_fu_8219_p2 = (xor_ln1545_131_fu_8213_p2 ^ xor_ln1545_129_fu_8207_p2);

assign xor_ln1545_131_fu_8213_p2 = (tmp_199_fu_7889_p4 ^ tmp_194_fu_7845_p4);

assign xor_ln1545_132_fu_8225_p2 = (trunc_ln674_42_fu_7807_p1 ^ tmp_187_fu_7787_p4);

assign xor_ln1545_133_fu_8231_p2 = (tmp_198_fu_7879_p4 ^ tmp_196_fu_7865_p4);

assign xor_ln1545_135_fu_8243_p2 = (tmp_191_fu_7821_p4 ^ tmp_186_fu_7777_p4);

assign xor_ln1545_136_fu_8255_p2 = (xor_ln1545_137_fu_8249_p2 ^ xor_ln1545_135_fu_8243_p2);

assign xor_ln1545_137_fu_8249_p2 = (trunc_ln674_43_fu_7841_p1 ^ tmp_200_fu_7899_p4);

assign xor_ln1545_138_fu_8261_p2 = (tmp_206_fu_7947_p4 ^ tmp_204_fu_7933_p4);

assign xor_ln1545_139_fu_8273_p2 = (xor_ln1545_140_fu_8267_p2 ^ xor_ln1545_138_fu_8261_p2);

assign xor_ln1545_13_fu_5719_p2 = (xor_ln1545_14_fu_5713_p2 ^ xor_ln1545_12_fu_5707_p2);

assign xor_ln1545_140_fu_8267_p2 = (trunc_ln674_48_fu_8011_p1 ^ tmp_211_fu_7991_p4);

assign xor_ln1545_141_fu_8279_p2 = (trunc_ln674_45_fu_7909_p1 ^ tmp_208_fu_7967_p4);

assign xor_ln1545_142_fu_8285_p2 = (tmp_215_fu_8025_p4 ^ tmp_210_fu_7981_p4);

assign xor_ln1545_144_fu_8297_p2 = (trunc_ln674_46_fu_7943_p1 ^ tmp_203_fu_7923_p4);

assign xor_ln1545_145_fu_8303_p2 = (tmp_214_fu_8015_p4 ^ tmp_212_fu_8001_p4);

assign xor_ln1545_147_fu_8315_p2 = (tmp_207_fu_7957_p4 ^ tmp_202_fu_7913_p4);

assign xor_ln1545_148_fu_8327_p2 = (xor_ln1545_149_fu_8321_p2 ^ xor_ln1545_147_fu_8315_p2);

assign xor_ln1545_149_fu_8321_p2 = (trunc_ln674_47_fu_7977_p1 ^ tmp_216_fu_8035_p4);

assign xor_ln1545_14_fu_5713_p2 = (tmp_40_fu_5233_p4 ^ tmp_38_fu_5219_p4);

assign xor_ln1545_150_fu_9232_p2 = (tmp_221_fu_8726_p4 ^ tmp_219_fu_8712_p4);

assign xor_ln1545_151_fu_9244_p2 = (xor_ln1545_152_fu_9238_p2 ^ xor_ln1545_150_fu_9232_p2);

assign xor_ln1545_152_fu_9238_p2 = (trunc_ln674_52_fu_8790_p1 ^ tmp_226_fu_8770_p4);

assign xor_ln1545_153_fu_9250_p2 = (trunc_ln674_49_fu_8688_p1 ^ tmp_223_fu_8746_p4);

assign xor_ln1545_154_fu_9262_p2 = (xor_ln1545_155_fu_9256_p2 ^ xor_ln1545_153_fu_9250_p2);

assign xor_ln1545_155_fu_9256_p2 = (tmp_230_fu_8804_p4 ^ tmp_225_fu_8760_p4);

assign xor_ln1545_156_fu_9268_p2 = (trunc_ln674_50_fu_8722_p1 ^ tmp_218_fu_8702_p4);

assign xor_ln1545_157_fu_9280_p2 = (xor_ln1545_158_fu_9274_p2 ^ xor_ln1545_156_fu_9268_p2);

assign xor_ln1545_158_fu_9274_p2 = (tmp_229_fu_8794_p4 ^ tmp_227_fu_8780_p4);

assign xor_ln1545_159_fu_9286_p2 = (tmp_222_fu_8736_p4 ^ tmp_217_fu_8692_p4);

assign xor_ln1545_15_fu_5725_p2 = (tmp_33_fu_5175_p4 ^ tmp_28_fu_5131_p4);

assign xor_ln1545_160_fu_9292_p2 = (trunc_ln674_51_fu_8756_p1 ^ tmp_231_fu_8814_p4);

assign xor_ln1545_162_fu_9304_p2 = (tmp_237_fu_8862_p4 ^ tmp_235_fu_8848_p4);

assign xor_ln1545_163_fu_9316_p2 = (xor_ln1545_164_fu_9310_p2 ^ xor_ln1545_162_fu_9304_p2);

assign xor_ln1545_164_fu_9310_p2 = (trunc_ln674_56_fu_8926_p1 ^ tmp_242_fu_8906_p4);

assign xor_ln1545_165_fu_9322_p2 = (trunc_ln674_53_fu_8824_p1 ^ tmp_239_fu_8882_p4);

assign xor_ln1545_166_fu_9334_p2 = (xor_ln1545_167_fu_9328_p2 ^ xor_ln1545_165_fu_9322_p2);

assign xor_ln1545_167_fu_9328_p2 = (tmp_246_fu_8940_p4 ^ tmp_241_fu_8896_p4);

assign xor_ln1545_168_fu_9340_p2 = (trunc_ln674_54_fu_8858_p1 ^ tmp_234_fu_8838_p4);

assign xor_ln1545_169_fu_9352_p2 = (xor_ln1545_170_fu_9346_p2 ^ xor_ln1545_168_fu_9340_p2);

assign xor_ln1545_16_fu_5731_p2 = (trunc_ln674_3_fu_5195_p1 ^ tmp_42_fu_5253_p4);

assign xor_ln1545_170_fu_9346_p2 = (tmp_245_fu_8930_p4 ^ tmp_243_fu_8916_p4);

assign xor_ln1545_171_fu_9358_p2 = (tmp_238_fu_8872_p4 ^ tmp_233_fu_8828_p4);

assign xor_ln1545_172_fu_9370_p2 = (xor_ln1545_173_fu_9364_p2 ^ xor_ln1545_171_fu_9358_p2);

assign xor_ln1545_173_fu_9364_p2 = (trunc_ln674_55_fu_8892_p1 ^ tmp_247_fu_8950_p4);

assign xor_ln1545_174_fu_9376_p2 = (tmp_253_fu_8998_p4 ^ tmp_251_fu_8984_p4);

assign xor_ln1545_175_fu_9388_p2 = (xor_ln1545_176_fu_9382_p2 ^ xor_ln1545_174_fu_9376_p2);

assign xor_ln1545_176_fu_9382_p2 = (trunc_ln674_60_fu_9062_p1 ^ tmp_258_fu_9042_p4);

assign xor_ln1545_177_fu_9394_p2 = (trunc_ln674_57_fu_8960_p1 ^ tmp_255_fu_9018_p4);

assign xor_ln1545_178_fu_9406_p2 = (xor_ln1545_179_fu_9400_p2 ^ xor_ln1545_177_fu_9394_p2);

assign xor_ln1545_179_fu_9400_p2 = (tmp_262_fu_9076_p4 ^ tmp_257_fu_9032_p4);

assign xor_ln1545_180_fu_9412_p2 = (trunc_ln674_58_fu_8994_p1 ^ tmp_250_fu_8974_p4);

assign xor_ln1545_181_fu_9418_p2 = (tmp_261_fu_9066_p4 ^ tmp_259_fu_9052_p4);

assign xor_ln1545_183_fu_9430_p2 = (tmp_254_fu_9008_p4 ^ tmp_249_fu_8964_p4);

assign xor_ln1545_184_fu_9442_p2 = (xor_ln1545_185_fu_9436_p2 ^ xor_ln1545_183_fu_9430_p2);

assign xor_ln1545_185_fu_9436_p2 = (trunc_ln674_59_fu_9028_p1 ^ tmp_263_fu_9086_p4);

assign xor_ln1545_186_fu_9448_p2 = (tmp_269_fu_9134_p4 ^ tmp_267_fu_9120_p4);

assign xor_ln1545_187_fu_9460_p2 = (xor_ln1545_188_fu_9454_p2 ^ xor_ln1545_186_fu_9448_p2);

assign xor_ln1545_188_fu_9454_p2 = (trunc_ln674_64_fu_9198_p1 ^ tmp_274_fu_9178_p4);

assign xor_ln1545_189_fu_9466_p2 = (trunc_ln674_61_fu_9096_p1 ^ tmp_271_fu_9154_p4);

assign xor_ln1545_18_fu_5743_p2 = (tmp_48_fu_5301_p4 ^ tmp_46_fu_5287_p4);

assign xor_ln1545_190_fu_9472_p2 = (tmp_278_fu_9212_p4 ^ tmp_273_fu_9168_p4);

assign xor_ln1545_192_fu_9484_p2 = (trunc_ln674_62_fu_9130_p1 ^ tmp_266_fu_9110_p4);

assign xor_ln1545_193_fu_9490_p2 = (tmp_277_fu_9202_p4 ^ tmp_275_fu_9188_p4);

assign xor_ln1545_195_fu_9502_p2 = (tmp_270_fu_9144_p4 ^ tmp_265_fu_9100_p4);

assign xor_ln1545_196_fu_9514_p2 = (xor_ln1545_197_fu_9508_p2 ^ xor_ln1545_195_fu_9502_p2);

assign xor_ln1545_197_fu_9508_p2 = (trunc_ln674_63_fu_9164_p1 ^ tmp_279_fu_9222_p4);

assign xor_ln1545_198_fu_10419_p2 = (tmp_284_fu_9913_p4 ^ tmp_282_fu_9899_p4);

assign xor_ln1545_199_fu_10431_p2 = (xor_ln1545_200_fu_10425_p2 ^ xor_ln1545_198_fu_10419_p2);

assign xor_ln1545_19_fu_5755_p2 = (xor_ln1545_20_fu_5749_p2 ^ xor_ln1545_18_fu_5743_p2);

assign xor_ln1545_200_fu_10425_p2 = (trunc_ln674_68_fu_9977_p1 ^ tmp_289_fu_9957_p4);

assign xor_ln1545_201_fu_10437_p2 = (trunc_ln674_65_fu_9875_p1 ^ tmp_286_fu_9933_p4);

assign xor_ln1545_202_fu_10449_p2 = (xor_ln1545_203_fu_10443_p2 ^ xor_ln1545_201_fu_10437_p2);

assign xor_ln1545_203_fu_10443_p2 = (tmp_293_fu_9991_p4 ^ tmp_288_fu_9947_p4);

assign xor_ln1545_204_fu_10455_p2 = (trunc_ln674_66_fu_9909_p1 ^ tmp_281_fu_9889_p4);

assign xor_ln1545_205_fu_10467_p2 = (xor_ln1545_206_fu_10461_p2 ^ xor_ln1545_204_fu_10455_p2);

assign xor_ln1545_206_fu_10461_p2 = (tmp_292_fu_9981_p4 ^ tmp_290_fu_9967_p4);

assign xor_ln1545_207_fu_10473_p2 = (tmp_285_fu_9923_p4 ^ tmp_280_fu_9879_p4);

assign xor_ln1545_208_fu_10479_p2 = (trunc_ln674_67_fu_9943_p1 ^ tmp_294_fu_10001_p4);

assign xor_ln1545_20_fu_5749_p2 = (trunc_ln674_8_fu_5365_p1 ^ tmp_53_fu_5345_p4);

assign xor_ln1545_210_fu_10491_p2 = (tmp_300_fu_10049_p4 ^ tmp_298_fu_10035_p4);

assign xor_ln1545_211_fu_10503_p2 = (xor_ln1545_212_fu_10497_p2 ^ xor_ln1545_210_fu_10491_p2);

assign xor_ln1545_212_fu_10497_p2 = (trunc_ln674_72_fu_10113_p1 ^ tmp_305_fu_10093_p4);

assign xor_ln1545_213_fu_10509_p2 = (trunc_ln674_69_fu_10011_p1 ^ tmp_302_fu_10069_p4);

assign xor_ln1545_214_fu_10521_p2 = (xor_ln1545_215_fu_10515_p2 ^ xor_ln1545_213_fu_10509_p2);

assign xor_ln1545_215_fu_10515_p2 = (tmp_309_fu_10127_p4 ^ tmp_304_fu_10083_p4);

assign xor_ln1545_216_fu_10527_p2 = (trunc_ln674_70_fu_10045_p1 ^ tmp_297_fu_10025_p4);

assign xor_ln1545_217_fu_10539_p2 = (xor_ln1545_218_fu_10533_p2 ^ xor_ln1545_216_fu_10527_p2);

assign xor_ln1545_218_fu_10533_p2 = (tmp_308_fu_10117_p4 ^ tmp_306_fu_10103_p4);

assign xor_ln1545_219_fu_10545_p2 = (tmp_301_fu_10059_p4 ^ tmp_296_fu_10015_p4);

assign xor_ln1545_21_fu_5761_p2 = (trunc_ln674_5_fu_5263_p1 ^ tmp_50_fu_5321_p4);

assign xor_ln1545_220_fu_10557_p2 = (xor_ln1545_221_fu_10551_p2 ^ xor_ln1545_219_fu_10545_p2);

assign xor_ln1545_221_fu_10551_p2 = (trunc_ln674_71_fu_10079_p1 ^ tmp_310_fu_10137_p4);

assign xor_ln1545_222_fu_10563_p2 = (tmp_316_fu_10185_p4 ^ tmp_314_fu_10171_p4);

assign xor_ln1545_223_fu_10575_p2 = (xor_ln1545_224_fu_10569_p2 ^ xor_ln1545_222_fu_10563_p2);

assign xor_ln1545_224_fu_10569_p2 = (trunc_ln674_76_fu_10249_p1 ^ tmp_321_fu_10229_p4);

assign xor_ln1545_225_fu_10581_p2 = (trunc_ln674_73_fu_10147_p1 ^ tmp_318_fu_10205_p4);

assign xor_ln1545_226_fu_10593_p2 = (xor_ln1545_227_fu_10587_p2 ^ xor_ln1545_225_fu_10581_p2);

assign xor_ln1545_227_fu_10587_p2 = (tmp_325_fu_10263_p4 ^ tmp_320_fu_10219_p4);

assign xor_ln1545_228_fu_10599_p2 = (trunc_ln674_74_fu_10181_p1 ^ tmp_313_fu_10161_p4);

assign xor_ln1545_229_fu_10605_p2 = (tmp_324_fu_10253_p4 ^ tmp_322_fu_10239_p4);

assign xor_ln1545_22_fu_5773_p2 = (xor_ln1545_23_fu_5767_p2 ^ xor_ln1545_21_fu_5761_p2);

assign xor_ln1545_231_fu_10617_p2 = (tmp_317_fu_10195_p4 ^ tmp_312_fu_10151_p4);

assign xor_ln1545_232_fu_10629_p2 = (xor_ln1545_233_fu_10623_p2 ^ xor_ln1545_231_fu_10617_p2);

assign xor_ln1545_233_fu_10623_p2 = (trunc_ln674_75_fu_10215_p1 ^ tmp_326_fu_10273_p4);

assign xor_ln1545_234_fu_10635_p2 = (tmp_332_fu_10321_p4 ^ tmp_330_fu_10307_p4);

assign xor_ln1545_235_fu_10647_p2 = (xor_ln1545_236_fu_10641_p2 ^ xor_ln1545_234_fu_10635_p2);

assign xor_ln1545_236_fu_10641_p2 = (trunc_ln674_80_fu_10385_p1 ^ tmp_337_fu_10365_p4);

assign xor_ln1545_237_fu_10653_p2 = (trunc_ln674_77_fu_10283_p1 ^ tmp_334_fu_10341_p4);

assign xor_ln1545_238_fu_10659_p2 = (tmp_341_fu_10399_p4 ^ tmp_336_fu_10355_p4);

assign xor_ln1545_23_fu_5767_p2 = (tmp_57_fu_5379_p4 ^ tmp_52_fu_5335_p4);

assign xor_ln1545_240_fu_10671_p2 = (trunc_ln674_78_fu_10317_p1 ^ tmp_329_fu_10297_p4);

assign xor_ln1545_241_fu_10677_p2 = (tmp_340_fu_10389_p4 ^ tmp_338_fu_10375_p4);

assign xor_ln1545_243_fu_10689_p2 = (tmp_333_fu_10331_p4 ^ tmp_328_fu_10287_p4);

assign xor_ln1545_244_fu_10701_p2 = (xor_ln1545_245_fu_10695_p2 ^ xor_ln1545_243_fu_10689_p2);

assign xor_ln1545_245_fu_10695_p2 = (trunc_ln674_79_fu_10351_p1 ^ tmp_342_fu_10409_p4);

assign xor_ln1545_246_fu_11606_p2 = (tmp_347_fu_11100_p4 ^ tmp_345_fu_11086_p4);

assign xor_ln1545_247_fu_11618_p2 = (xor_ln1545_248_fu_11612_p2 ^ xor_ln1545_246_fu_11606_p2);

assign xor_ln1545_248_fu_11612_p2 = (trunc_ln674_84_fu_11164_p1 ^ tmp_352_fu_11144_p4);

assign xor_ln1545_249_fu_11624_p2 = (trunc_ln674_81_fu_11062_p1 ^ tmp_349_fu_11120_p4);

assign xor_ln1545_24_fu_5779_p2 = (trunc_ln674_6_fu_5297_p1 ^ tmp_45_fu_5277_p4);

assign xor_ln1545_250_fu_11636_p2 = (xor_ln1545_251_fu_11630_p2 ^ xor_ln1545_249_fu_11624_p2);

assign xor_ln1545_251_fu_11630_p2 = (tmp_356_fu_11178_p4 ^ tmp_351_fu_11134_p4);

assign xor_ln1545_252_fu_11642_p2 = (trunc_ln674_82_fu_11096_p1 ^ tmp_344_fu_11076_p4);

assign xor_ln1545_253_fu_11654_p2 = (xor_ln1545_254_fu_11648_p2 ^ xor_ln1545_252_fu_11642_p2);

assign xor_ln1545_254_fu_11648_p2 = (tmp_355_fu_11168_p4 ^ tmp_353_fu_11154_p4);

assign xor_ln1545_255_fu_11660_p2 = (tmp_348_fu_11110_p4 ^ tmp_343_fu_11066_p4);

assign xor_ln1545_256_fu_11666_p2 = (trunc_ln674_83_fu_11130_p1 ^ tmp_357_fu_11188_p4);

assign xor_ln1545_258_fu_11678_p2 = (tmp_363_fu_11236_p4 ^ tmp_361_fu_11222_p4);

assign xor_ln1545_259_fu_11690_p2 = (xor_ln1545_260_fu_11684_p2 ^ xor_ln1545_258_fu_11678_p2);

assign xor_ln1545_25_fu_5791_p2 = (xor_ln1545_26_fu_5785_p2 ^ xor_ln1545_24_fu_5779_p2);

assign xor_ln1545_260_fu_11684_p2 = (trunc_ln674_88_fu_11300_p1 ^ tmp_368_fu_11280_p4);

assign xor_ln1545_261_fu_11696_p2 = (trunc_ln674_85_fu_11198_p1 ^ tmp_365_fu_11256_p4);

assign xor_ln1545_262_fu_11708_p2 = (xor_ln1545_263_fu_11702_p2 ^ xor_ln1545_261_fu_11696_p2);

assign xor_ln1545_263_fu_11702_p2 = (tmp_372_fu_11314_p4 ^ tmp_367_fu_11270_p4);

assign xor_ln1545_264_fu_11714_p2 = (trunc_ln674_86_fu_11232_p1 ^ tmp_360_fu_11212_p4);

assign xor_ln1545_265_fu_11726_p2 = (xor_ln1545_266_fu_11720_p2 ^ xor_ln1545_264_fu_11714_p2);

assign xor_ln1545_266_fu_11720_p2 = (tmp_371_fu_11304_p4 ^ tmp_369_fu_11290_p4);

assign xor_ln1545_267_fu_11732_p2 = (tmp_364_fu_11246_p4 ^ tmp_359_fu_11202_p4);

assign xor_ln1545_268_fu_11744_p2 = (xor_ln1545_269_fu_11738_p2 ^ xor_ln1545_267_fu_11732_p2);

assign xor_ln1545_269_fu_11738_p2 = (trunc_ln674_87_fu_11266_p1 ^ tmp_373_fu_11324_p4);

assign xor_ln1545_26_fu_5785_p2 = (tmp_56_fu_5369_p4 ^ tmp_54_fu_5355_p4);

assign xor_ln1545_270_fu_11750_p2 = (tmp_379_fu_11372_p4 ^ tmp_377_fu_11358_p4);

assign xor_ln1545_271_fu_11762_p2 = (xor_ln1545_272_fu_11756_p2 ^ xor_ln1545_270_fu_11750_p2);

assign xor_ln1545_272_fu_11756_p2 = (trunc_ln674_92_fu_11436_p1 ^ tmp_384_fu_11416_p4);

assign xor_ln1545_273_fu_11768_p2 = (trunc_ln674_89_fu_11334_p1 ^ tmp_381_fu_11392_p4);

assign xor_ln1545_274_fu_11780_p2 = (xor_ln1545_275_fu_11774_p2 ^ xor_ln1545_273_fu_11768_p2);

assign xor_ln1545_275_fu_11774_p2 = (tmp_388_fu_11450_p4 ^ tmp_383_fu_11406_p4);

assign xor_ln1545_276_fu_11786_p2 = (trunc_ln674_90_fu_11368_p1 ^ tmp_376_fu_11348_p4);

assign xor_ln1545_277_fu_11792_p2 = (tmp_387_fu_11440_p4 ^ tmp_385_fu_11426_p4);

assign xor_ln1545_279_fu_11804_p2 = (tmp_380_fu_11382_p4 ^ tmp_375_fu_11338_p4);

assign xor_ln1545_27_fu_5797_p2 = (tmp_49_fu_5311_p4 ^ tmp_44_fu_5267_p4);

assign xor_ln1545_280_fu_11816_p2 = (xor_ln1545_281_fu_11810_p2 ^ xor_ln1545_279_fu_11804_p2);

assign xor_ln1545_281_fu_11810_p2 = (trunc_ln674_91_fu_11402_p1 ^ tmp_389_fu_11460_p4);

assign xor_ln1545_282_fu_11822_p2 = (tmp_395_fu_11508_p4 ^ tmp_393_fu_11494_p4);

assign xor_ln1545_283_fu_11834_p2 = (xor_ln1545_284_fu_11828_p2 ^ xor_ln1545_282_fu_11822_p2);

assign xor_ln1545_284_fu_11828_p2 = (trunc_ln674_96_fu_11572_p1 ^ tmp_400_fu_11552_p4);

assign xor_ln1545_285_fu_11840_p2 = (trunc_ln674_93_fu_11470_p1 ^ tmp_397_fu_11528_p4);

assign xor_ln1545_286_fu_11846_p2 = (tmp_404_fu_11586_p4 ^ tmp_399_fu_11542_p4);

assign xor_ln1545_288_fu_11858_p2 = (trunc_ln674_94_fu_11504_p1 ^ tmp_392_fu_11484_p4);

assign xor_ln1545_289_fu_11864_p2 = (tmp_403_fu_11576_p4 ^ tmp_401_fu_11562_p4);

assign xor_ln1545_28_fu_5809_p2 = (xor_ln1545_29_fu_5803_p2 ^ xor_ln1545_27_fu_5797_p2);

assign xor_ln1545_291_fu_11876_p2 = (tmp_396_fu_11518_p4 ^ tmp_391_fu_11474_p4);

assign xor_ln1545_292_fu_11888_p2 = (xor_ln1545_293_fu_11882_p2 ^ xor_ln1545_291_fu_11876_p2);

assign xor_ln1545_293_fu_11882_p2 = (trunc_ln674_95_fu_11538_p1 ^ tmp_405_fu_11596_p4);

assign xor_ln1545_294_fu_12793_p2 = (tmp_410_fu_12287_p4 ^ tmp_408_fu_12273_p4);

assign xor_ln1545_295_fu_12805_p2 = (xor_ln1545_296_fu_12799_p2 ^ xor_ln1545_294_fu_12793_p2);

assign xor_ln1545_296_fu_12799_p2 = (trunc_ln674_100_fu_12351_p1 ^ tmp_415_fu_12331_p4);

assign xor_ln1545_297_fu_12811_p2 = (trunc_ln674_97_fu_12249_p1 ^ tmp_412_fu_12307_p4);

assign xor_ln1545_298_fu_12823_p2 = (xor_ln1545_299_fu_12817_p2 ^ xor_ln1545_297_fu_12811_p2);

assign xor_ln1545_299_fu_12817_p2 = (tmp_419_fu_12365_p4 ^ tmp_414_fu_12321_p4);

assign xor_ln1545_29_fu_5803_p2 = (trunc_ln674_7_fu_5331_p1 ^ tmp_58_fu_5389_p4);

assign xor_ln1545_300_fu_12829_p2 = (trunc_ln674_98_fu_12283_p1 ^ tmp_407_fu_12263_p4);

assign xor_ln1545_301_fu_12841_p2 = (xor_ln1545_302_fu_12835_p2 ^ xor_ln1545_300_fu_12829_p2);

assign xor_ln1545_302_fu_12835_p2 = (tmp_418_fu_12355_p4 ^ tmp_416_fu_12341_p4);

assign xor_ln1545_303_fu_12847_p2 = (tmp_411_fu_12297_p4 ^ tmp_406_fu_12253_p4);

assign xor_ln1545_304_fu_12853_p2 = (trunc_ln674_99_fu_12317_p1 ^ tmp_420_fu_12375_p4);

assign xor_ln1545_306_fu_12865_p2 = (tmp_426_fu_12423_p4 ^ tmp_424_fu_12409_p4);

assign xor_ln1545_307_fu_12877_p2 = (xor_ln1545_308_fu_12871_p2 ^ xor_ln1545_306_fu_12865_p2);

assign xor_ln1545_308_fu_12871_p2 = (trunc_ln674_104_fu_12487_p1 ^ tmp_431_fu_12467_p4);

assign xor_ln1545_309_fu_12883_p2 = (trunc_ln674_101_fu_12385_p1 ^ tmp_428_fu_12443_p4);

assign xor_ln1545_30_fu_5815_p2 = (tmp_64_fu_5437_p4 ^ tmp_62_fu_5423_p4);

assign xor_ln1545_310_fu_12895_p2 = (xor_ln1545_311_fu_12889_p2 ^ xor_ln1545_309_fu_12883_p2);

assign xor_ln1545_311_fu_12889_p2 = (tmp_435_fu_12501_p4 ^ tmp_430_fu_12457_p4);

assign xor_ln1545_312_fu_12901_p2 = (trunc_ln674_102_fu_12419_p1 ^ tmp_423_fu_12399_p4);

assign xor_ln1545_313_fu_12913_p2 = (xor_ln1545_314_fu_12907_p2 ^ xor_ln1545_312_fu_12901_p2);

assign xor_ln1545_314_fu_12907_p2 = (tmp_434_fu_12491_p4 ^ tmp_432_fu_12477_p4);

assign xor_ln1545_315_fu_12919_p2 = (tmp_427_fu_12433_p4 ^ tmp_422_fu_12389_p4);

assign xor_ln1545_316_fu_12931_p2 = (xor_ln1545_317_fu_12925_p2 ^ xor_ln1545_315_fu_12919_p2);

assign xor_ln1545_317_fu_12925_p2 = (trunc_ln674_103_fu_12453_p1 ^ tmp_436_fu_12511_p4);

assign xor_ln1545_318_fu_12937_p2 = (tmp_442_fu_12559_p4 ^ tmp_440_fu_12545_p4);

assign xor_ln1545_319_fu_12949_p2 = (xor_ln1545_320_fu_12943_p2 ^ xor_ln1545_318_fu_12937_p2);

assign xor_ln1545_31_fu_5827_p2 = (xor_ln1545_32_fu_5821_p2 ^ xor_ln1545_30_fu_5815_p2);

assign xor_ln1545_320_fu_12943_p2 = (trunc_ln674_108_fu_12623_p1 ^ tmp_447_fu_12603_p4);

assign xor_ln1545_321_fu_12955_p2 = (trunc_ln674_105_fu_12521_p1 ^ tmp_444_fu_12579_p4);

assign xor_ln1545_322_fu_12967_p2 = (xor_ln1545_323_fu_12961_p2 ^ xor_ln1545_321_fu_12955_p2);

assign xor_ln1545_323_fu_12961_p2 = (tmp_451_fu_12637_p4 ^ tmp_446_fu_12593_p4);

assign xor_ln1545_324_fu_12973_p2 = (trunc_ln674_106_fu_12555_p1 ^ tmp_439_fu_12535_p4);

assign xor_ln1545_325_fu_12979_p2 = (tmp_450_fu_12627_p4 ^ tmp_448_fu_12613_p4);

assign xor_ln1545_327_fu_12991_p2 = (tmp_443_fu_12569_p4 ^ tmp_438_fu_12525_p4);

assign xor_ln1545_328_fu_13003_p2 = (xor_ln1545_329_fu_12997_p2 ^ xor_ln1545_327_fu_12991_p2);

assign xor_ln1545_329_fu_12997_p2 = (trunc_ln674_107_fu_12589_p1 ^ tmp_452_fu_12647_p4);

assign xor_ln1545_32_fu_5821_p2 = (trunc_ln674_12_fu_5501_p1 ^ tmp_69_fu_5481_p4);

assign xor_ln1545_330_fu_13009_p2 = (tmp_458_fu_12695_p4 ^ tmp_456_fu_12681_p4);

assign xor_ln1545_331_fu_13021_p2 = (xor_ln1545_332_fu_13015_p2 ^ xor_ln1545_330_fu_13009_p2);

assign xor_ln1545_332_fu_13015_p2 = (trunc_ln674_112_fu_12759_p1 ^ tmp_463_fu_12739_p4);

assign xor_ln1545_333_fu_13027_p2 = (trunc_ln674_109_fu_12657_p1 ^ tmp_460_fu_12715_p4);

assign xor_ln1545_334_fu_13033_p2 = (tmp_467_fu_12773_p4 ^ tmp_462_fu_12729_p4);

assign xor_ln1545_336_fu_13045_p2 = (trunc_ln674_110_fu_12691_p1 ^ tmp_455_fu_12671_p4);

assign xor_ln1545_337_fu_13051_p2 = (tmp_466_fu_12763_p4 ^ tmp_464_fu_12749_p4);

assign xor_ln1545_339_fu_13063_p2 = (tmp_459_fu_12705_p4 ^ tmp_454_fu_12661_p4);

assign xor_ln1545_33_fu_5833_p2 = (trunc_ln674_9_fu_5399_p1 ^ tmp_66_fu_5457_p4);

assign xor_ln1545_340_fu_13075_p2 = (xor_ln1545_341_fu_13069_p2 ^ xor_ln1545_339_fu_13063_p2);

assign xor_ln1545_341_fu_13069_p2 = (trunc_ln674_111_fu_12725_p1 ^ tmp_468_fu_12783_p4);

assign xor_ln1545_342_fu_13980_p2 = (tmp_473_fu_13474_p4 ^ tmp_471_fu_13460_p4);

assign xor_ln1545_343_fu_13992_p2 = (xor_ln1545_344_fu_13986_p2 ^ xor_ln1545_342_fu_13980_p2);

assign xor_ln1545_344_fu_13986_p2 = (trunc_ln674_116_fu_13538_p1 ^ tmp_478_fu_13518_p4);

assign xor_ln1545_345_fu_13998_p2 = (trunc_ln674_113_fu_13436_p1 ^ tmp_475_fu_13494_p4);

assign xor_ln1545_346_fu_14010_p2 = (xor_ln1545_347_fu_14004_p2 ^ xor_ln1545_345_fu_13998_p2);

assign xor_ln1545_347_fu_14004_p2 = (tmp_482_fu_13552_p4 ^ tmp_477_fu_13508_p4);

assign xor_ln1545_348_fu_14016_p2 = (trunc_ln674_114_fu_13470_p1 ^ tmp_470_fu_13450_p4);

assign xor_ln1545_349_fu_14028_p2 = (xor_ln1545_350_fu_14022_p2 ^ xor_ln1545_348_fu_14016_p2);

assign xor_ln1545_34_fu_5845_p2 = (xor_ln1545_35_fu_5839_p2 ^ xor_ln1545_33_fu_5833_p2);

assign xor_ln1545_350_fu_14022_p2 = (tmp_481_fu_13542_p4 ^ tmp_479_fu_13528_p4);

assign xor_ln1545_351_fu_14034_p2 = (tmp_474_fu_13484_p4 ^ tmp_469_fu_13440_p4);

assign xor_ln1545_352_fu_14040_p2 = (trunc_ln674_115_fu_13504_p1 ^ tmp_483_fu_13562_p4);

assign xor_ln1545_354_fu_14052_p2 = (tmp_489_fu_13610_p4 ^ tmp_487_fu_13596_p4);

assign xor_ln1545_355_fu_14064_p2 = (xor_ln1545_356_fu_14058_p2 ^ xor_ln1545_354_fu_14052_p2);

assign xor_ln1545_356_fu_14058_p2 = (trunc_ln674_120_fu_13674_p1 ^ tmp_494_fu_13654_p4);

assign xor_ln1545_357_fu_14070_p2 = (trunc_ln674_117_fu_13572_p1 ^ tmp_491_fu_13630_p4);

assign xor_ln1545_358_fu_14082_p2 = (xor_ln1545_359_fu_14076_p2 ^ xor_ln1545_357_fu_14070_p2);

assign xor_ln1545_359_fu_14076_p2 = (tmp_498_fu_13688_p4 ^ tmp_493_fu_13644_p4);

assign xor_ln1545_35_fu_5839_p2 = (tmp_73_fu_5515_p4 ^ tmp_68_fu_5471_p4);

assign xor_ln1545_360_fu_14088_p2 = (trunc_ln674_118_fu_13606_p1 ^ tmp_486_fu_13586_p4);

assign xor_ln1545_361_fu_14100_p2 = (xor_ln1545_362_fu_14094_p2 ^ xor_ln1545_360_fu_14088_p2);

assign xor_ln1545_362_fu_14094_p2 = (tmp_497_fu_13678_p4 ^ tmp_495_fu_13664_p4);

assign xor_ln1545_363_fu_14106_p2 = (tmp_490_fu_13620_p4 ^ tmp_485_fu_13576_p4);

assign xor_ln1545_364_fu_14118_p2 = (xor_ln1545_365_fu_14112_p2 ^ xor_ln1545_363_fu_14106_p2);

assign xor_ln1545_365_fu_14112_p2 = (trunc_ln674_119_fu_13640_p1 ^ tmp_499_fu_13698_p4);

assign xor_ln1545_366_fu_14124_p2 = (tmp_505_fu_13746_p4 ^ tmp_503_fu_13732_p4);

assign xor_ln1545_367_fu_14136_p2 = (xor_ln1545_368_fu_14130_p2 ^ xor_ln1545_366_fu_14124_p2);

assign xor_ln1545_368_fu_14130_p2 = (trunc_ln674_124_fu_13810_p1 ^ tmp_510_fu_13790_p4);

assign xor_ln1545_369_fu_14142_p2 = (trunc_ln674_121_fu_13708_p1 ^ tmp_507_fu_13766_p4);

assign xor_ln1545_36_fu_5851_p2 = (trunc_ln674_10_fu_5433_p1 ^ tmp_61_fu_5413_p4);

assign xor_ln1545_370_fu_14154_p2 = (xor_ln1545_371_fu_14148_p2 ^ xor_ln1545_369_fu_14142_p2);

assign xor_ln1545_371_fu_14148_p2 = (tmp_514_fu_13824_p4 ^ tmp_509_fu_13780_p4);

assign xor_ln1545_372_fu_14160_p2 = (trunc_ln674_122_fu_13742_p1 ^ tmp_502_fu_13722_p4);

assign xor_ln1545_373_fu_14166_p2 = (tmp_513_fu_13814_p4 ^ tmp_511_fu_13800_p4);

assign xor_ln1545_375_fu_14178_p2 = (tmp_506_fu_13756_p4 ^ tmp_501_fu_13712_p4);

assign xor_ln1545_376_fu_14190_p2 = (xor_ln1545_377_fu_14184_p2 ^ xor_ln1545_375_fu_14178_p2);

assign xor_ln1545_377_fu_14184_p2 = (trunc_ln674_123_fu_13776_p1 ^ tmp_515_fu_13834_p4);

assign xor_ln1545_378_fu_14196_p2 = (tmp_521_fu_13882_p4 ^ tmp_519_fu_13868_p4);

assign xor_ln1545_379_fu_14208_p2 = (xor_ln1545_380_fu_14202_p2 ^ xor_ln1545_378_fu_14196_p2);

assign xor_ln1545_37_fu_5857_p2 = (tmp_72_fu_5505_p4 ^ tmp_70_fu_5491_p4);

assign xor_ln1545_380_fu_14202_p2 = (trunc_ln674_128_fu_13946_p1 ^ tmp_526_fu_13926_p4);

assign xor_ln1545_381_fu_14214_p2 = (trunc_ln674_125_fu_13844_p1 ^ tmp_523_fu_13902_p4);

assign xor_ln1545_382_fu_14220_p2 = (tmp_530_fu_13960_p4 ^ tmp_525_fu_13916_p4);

assign xor_ln1545_384_fu_14232_p2 = (trunc_ln674_126_fu_13878_p1 ^ tmp_518_fu_13858_p4);

assign xor_ln1545_385_fu_14238_p2 = (tmp_529_fu_13950_p4 ^ tmp_527_fu_13936_p4);

assign xor_ln1545_387_fu_14250_p2 = (tmp_522_fu_13892_p4 ^ tmp_517_fu_13848_p4);

assign xor_ln1545_388_fu_14262_p2 = (xor_ln1545_389_fu_14256_p2 ^ xor_ln1545_387_fu_14250_p2);

assign xor_ln1545_389_fu_14256_p2 = (trunc_ln674_127_fu_13912_p1 ^ tmp_531_fu_13970_p4);

assign xor_ln1545_390_fu_15167_p2 = (tmp_536_fu_14661_p4 ^ tmp_534_fu_14647_p4);

assign xor_ln1545_391_fu_15179_p2 = (xor_ln1545_392_fu_15173_p2 ^ xor_ln1545_390_fu_15167_p2);

assign xor_ln1545_392_fu_15173_p2 = (trunc_ln674_132_fu_14725_p1 ^ tmp_541_fu_14705_p4);

assign xor_ln1545_393_fu_15185_p2 = (trunc_ln674_129_fu_14623_p1 ^ tmp_538_fu_14681_p4);

assign xor_ln1545_394_fu_15197_p2 = (xor_ln1545_395_fu_15191_p2 ^ xor_ln1545_393_fu_15185_p2);

assign xor_ln1545_395_fu_15191_p2 = (tmp_545_fu_14739_p4 ^ tmp_540_fu_14695_p4);

assign xor_ln1545_396_fu_15203_p2 = (trunc_ln674_130_fu_14657_p1 ^ tmp_533_fu_14637_p4);

assign xor_ln1545_397_fu_15215_p2 = (xor_ln1545_398_fu_15209_p2 ^ xor_ln1545_396_fu_15203_p2);

assign xor_ln1545_398_fu_15209_p2 = (tmp_544_fu_14729_p4 ^ tmp_542_fu_14715_p4);

assign xor_ln1545_399_fu_15221_p2 = (tmp_537_fu_14671_p4 ^ tmp_532_fu_14627_p4);

assign xor_ln1545_39_fu_5869_p2 = (tmp_65_fu_5447_p4 ^ tmp_60_fu_5403_p4);

assign xor_ln1545_400_fu_15227_p2 = (trunc_ln674_131_fu_14691_p1 ^ tmp_546_fu_14749_p4);

assign xor_ln1545_402_fu_15239_p2 = (tmp_552_fu_14797_p4 ^ tmp_550_fu_14783_p4);

assign xor_ln1545_403_fu_15251_p2 = (xor_ln1545_404_fu_15245_p2 ^ xor_ln1545_402_fu_15239_p2);

assign xor_ln1545_404_fu_15245_p2 = (trunc_ln674_136_fu_14861_p1 ^ tmp_557_fu_14841_p4);

assign xor_ln1545_405_fu_15257_p2 = (trunc_ln674_133_fu_14759_p1 ^ tmp_554_fu_14817_p4);

assign xor_ln1545_406_fu_15269_p2 = (xor_ln1545_407_fu_15263_p2 ^ xor_ln1545_405_fu_15257_p2);

assign xor_ln1545_407_fu_15263_p2 = (tmp_561_fu_14875_p4 ^ tmp_556_fu_14831_p4);

assign xor_ln1545_408_fu_15275_p2 = (trunc_ln674_134_fu_14793_p1 ^ tmp_549_fu_14773_p4);

assign xor_ln1545_409_fu_15287_p2 = (xor_ln1545_410_fu_15281_p2 ^ xor_ln1545_408_fu_15275_p2);

assign xor_ln1545_40_fu_5881_p2 = (xor_ln1545_41_fu_5875_p2 ^ xor_ln1545_39_fu_5869_p2);

assign xor_ln1545_410_fu_15281_p2 = (tmp_560_fu_14865_p4 ^ tmp_558_fu_14851_p4);

assign xor_ln1545_411_fu_15293_p2 = (tmp_553_fu_14807_p4 ^ tmp_548_fu_14763_p4);

assign xor_ln1545_412_fu_15305_p2 = (xor_ln1545_413_fu_15299_p2 ^ xor_ln1545_411_fu_15293_p2);

assign xor_ln1545_413_fu_15299_p2 = (trunc_ln674_135_fu_14827_p1 ^ tmp_562_fu_14885_p4);

assign xor_ln1545_414_fu_15311_p2 = (tmp_568_fu_14933_p4 ^ tmp_566_fu_14919_p4);

assign xor_ln1545_415_fu_15323_p2 = (xor_ln1545_416_fu_15317_p2 ^ xor_ln1545_414_fu_15311_p2);

assign xor_ln1545_416_fu_15317_p2 = (trunc_ln674_140_fu_14997_p1 ^ tmp_573_fu_14977_p4);

assign xor_ln1545_417_fu_15329_p2 = (trunc_ln674_137_fu_14895_p1 ^ tmp_570_fu_14953_p4);

assign xor_ln1545_418_fu_15341_p2 = (xor_ln1545_419_fu_15335_p2 ^ xor_ln1545_417_fu_15329_p2);

assign xor_ln1545_419_fu_15335_p2 = (tmp_577_fu_15011_p4 ^ tmp_572_fu_14967_p4);

assign xor_ln1545_41_fu_5875_p2 = (trunc_ln674_11_fu_5467_p1 ^ tmp_74_fu_5525_p4);

assign xor_ln1545_420_fu_15347_p2 = (trunc_ln674_138_fu_14929_p1 ^ tmp_565_fu_14909_p4);

assign xor_ln1545_421_fu_15353_p2 = (tmp_576_fu_15001_p4 ^ tmp_574_fu_14987_p4);

assign xor_ln1545_423_fu_15365_p2 = (tmp_569_fu_14943_p4 ^ tmp_564_fu_14899_p4);

assign xor_ln1545_424_fu_15377_p2 = (xor_ln1545_425_fu_15371_p2 ^ xor_ln1545_423_fu_15365_p2);

assign xor_ln1545_425_fu_15371_p2 = (trunc_ln674_139_fu_14963_p1 ^ tmp_578_fu_15021_p4);

assign xor_ln1545_426_fu_15383_p2 = (tmp_584_fu_15069_p4 ^ tmp_582_fu_15055_p4);

assign xor_ln1545_427_fu_15395_p2 = (xor_ln1545_428_fu_15389_p2 ^ xor_ln1545_426_fu_15383_p2);

assign xor_ln1545_428_fu_15389_p2 = (trunc_ln674_144_fu_15133_p1 ^ tmp_589_fu_15113_p4);

assign xor_ln1545_429_fu_15401_p2 = (trunc_ln674_141_fu_15031_p1 ^ tmp_586_fu_15089_p4);

assign xor_ln1545_42_fu_5887_p2 = (tmp_80_fu_5573_p4 ^ tmp_78_fu_5559_p4);

assign xor_ln1545_430_fu_15407_p2 = (tmp_593_fu_15147_p4 ^ tmp_588_fu_15103_p4);

assign xor_ln1545_432_fu_15419_p2 = (trunc_ln674_142_fu_15065_p1 ^ tmp_581_fu_15045_p4);

assign xor_ln1545_433_fu_15425_p2 = (tmp_592_fu_15137_p4 ^ tmp_590_fu_15123_p4);

assign xor_ln1545_435_fu_15437_p2 = (tmp_585_fu_15079_p4 ^ tmp_580_fu_15035_p4);

assign xor_ln1545_436_fu_15449_p2 = (xor_ln1545_437_fu_15443_p2 ^ xor_ln1545_435_fu_15437_p2);

assign xor_ln1545_437_fu_15443_p2 = (trunc_ln674_143_fu_15099_p1 ^ tmp_594_fu_15157_p4);

assign xor_ln1545_438_fu_16354_p2 = (tmp_599_fu_15848_p4 ^ tmp_597_fu_15834_p4);

assign xor_ln1545_439_fu_16366_p2 = (xor_ln1545_440_fu_16360_p2 ^ xor_ln1545_438_fu_16354_p2);

assign xor_ln1545_43_fu_5899_p2 = (xor_ln1545_44_fu_5893_p2 ^ xor_ln1545_42_fu_5887_p2);

assign xor_ln1545_440_fu_16360_p2 = (trunc_ln674_148_fu_15912_p1 ^ tmp_604_fu_15892_p4);

assign xor_ln1545_441_fu_16372_p2 = (trunc_ln674_145_fu_15810_p1 ^ tmp_601_fu_15868_p4);

assign xor_ln1545_442_fu_16384_p2 = (xor_ln1545_443_fu_16378_p2 ^ xor_ln1545_441_fu_16372_p2);

assign xor_ln1545_443_fu_16378_p2 = (tmp_608_fu_15926_p4 ^ tmp_603_fu_15882_p4);

assign xor_ln1545_444_fu_16390_p2 = (trunc_ln674_146_fu_15844_p1 ^ tmp_596_fu_15824_p4);

assign xor_ln1545_445_fu_16402_p2 = (xor_ln1545_446_fu_16396_p2 ^ xor_ln1545_444_fu_16390_p2);

assign xor_ln1545_446_fu_16396_p2 = (tmp_607_fu_15916_p4 ^ tmp_605_fu_15902_p4);

assign xor_ln1545_447_fu_16408_p2 = (tmp_600_fu_15858_p4 ^ tmp_595_fu_15814_p4);

assign xor_ln1545_448_fu_16414_p2 = (trunc_ln674_147_fu_15878_p1 ^ tmp_609_fu_15936_p4);

assign xor_ln1545_44_fu_5893_p2 = (trunc_ln674_16_fu_5637_p1 ^ tmp_85_fu_5617_p4);

assign xor_ln1545_450_fu_16426_p2 = (tmp_615_fu_15984_p4 ^ tmp_613_fu_15970_p4);

assign xor_ln1545_451_fu_16438_p2 = (xor_ln1545_452_fu_16432_p2 ^ xor_ln1545_450_fu_16426_p2);

assign xor_ln1545_452_fu_16432_p2 = (trunc_ln674_152_fu_16048_p1 ^ tmp_620_fu_16028_p4);

assign xor_ln1545_453_fu_16444_p2 = (trunc_ln674_149_fu_15946_p1 ^ tmp_617_fu_16004_p4);

assign xor_ln1545_454_fu_16456_p2 = (xor_ln1545_455_fu_16450_p2 ^ xor_ln1545_453_fu_16444_p2);

assign xor_ln1545_455_fu_16450_p2 = (tmp_624_fu_16062_p4 ^ tmp_619_fu_16018_p4);

assign xor_ln1545_456_fu_16462_p2 = (trunc_ln674_150_fu_15980_p1 ^ tmp_612_fu_15960_p4);

assign xor_ln1545_457_fu_16474_p2 = (xor_ln1545_458_fu_16468_p2 ^ xor_ln1545_456_fu_16462_p2);

assign xor_ln1545_458_fu_16468_p2 = (tmp_623_fu_16052_p4 ^ tmp_621_fu_16038_p4);

assign xor_ln1545_459_fu_16480_p2 = (tmp_616_fu_15994_p4 ^ tmp_611_fu_15950_p4);

assign xor_ln1545_45_fu_5905_p2 = (trunc_ln674_13_fu_5535_p1 ^ tmp_82_fu_5593_p4);

assign xor_ln1545_460_fu_16492_p2 = (xor_ln1545_461_fu_16486_p2 ^ xor_ln1545_459_fu_16480_p2);

assign xor_ln1545_461_fu_16486_p2 = (trunc_ln674_151_fu_16014_p1 ^ tmp_625_fu_16072_p4);

assign xor_ln1545_462_fu_16498_p2 = (tmp_631_fu_16120_p4 ^ tmp_629_fu_16106_p4);

assign xor_ln1545_463_fu_16510_p2 = (xor_ln1545_464_fu_16504_p2 ^ xor_ln1545_462_fu_16498_p2);

assign xor_ln1545_464_fu_16504_p2 = (trunc_ln674_156_fu_16184_p1 ^ tmp_636_fu_16164_p4);

assign xor_ln1545_465_fu_16516_p2 = (trunc_ln674_153_fu_16082_p1 ^ tmp_633_fu_16140_p4);

assign xor_ln1545_466_fu_16528_p2 = (xor_ln1545_467_fu_16522_p2 ^ xor_ln1545_465_fu_16516_p2);

assign xor_ln1545_467_fu_16522_p2 = (tmp_640_fu_16198_p4 ^ tmp_635_fu_16154_p4);

assign xor_ln1545_468_fu_16534_p2 = (trunc_ln674_154_fu_16116_p1 ^ tmp_628_fu_16096_p4);

assign xor_ln1545_469_fu_16540_p2 = (tmp_639_fu_16188_p4 ^ tmp_637_fu_16174_p4);

assign xor_ln1545_46_fu_5911_p2 = (tmp_89_fu_5651_p4 ^ tmp_84_fu_5607_p4);

assign xor_ln1545_471_fu_16552_p2 = (tmp_632_fu_16130_p4 ^ tmp_627_fu_16086_p4);

assign xor_ln1545_472_fu_16564_p2 = (xor_ln1545_473_fu_16558_p2 ^ xor_ln1545_471_fu_16552_p2);

assign xor_ln1545_473_fu_16558_p2 = (trunc_ln674_155_fu_16150_p1 ^ tmp_641_fu_16208_p4);

assign xor_ln1545_474_fu_16570_p2 = (tmp_647_fu_16256_p4 ^ tmp_645_fu_16242_p4);

assign xor_ln1545_475_fu_16582_p2 = (xor_ln1545_476_fu_16576_p2 ^ xor_ln1545_474_fu_16570_p2);

assign xor_ln1545_476_fu_16576_p2 = (trunc_ln674_160_fu_16320_p1 ^ tmp_652_fu_16300_p4);

assign xor_ln1545_477_fu_16588_p2 = (trunc_ln674_157_fu_16218_p1 ^ tmp_649_fu_16276_p4);

assign xor_ln1545_478_fu_16594_p2 = (tmp_656_fu_16334_p4 ^ tmp_651_fu_16290_p4);

assign xor_ln1545_480_fu_16606_p2 = (trunc_ln674_158_fu_16252_p1 ^ tmp_644_fu_16232_p4);

assign xor_ln1545_481_fu_16612_p2 = (tmp_655_fu_16324_p4 ^ tmp_653_fu_16310_p4);

assign xor_ln1545_483_fu_16624_p2 = (tmp_648_fu_16266_p4 ^ tmp_643_fu_16222_p4);

assign xor_ln1545_484_fu_16636_p2 = (xor_ln1545_485_fu_16630_p2 ^ xor_ln1545_483_fu_16624_p2);

assign xor_ln1545_485_fu_16630_p2 = (trunc_ln674_159_fu_16286_p1 ^ tmp_657_fu_16344_p4);

assign xor_ln1545_486_fu_17541_p2 = (tmp_662_fu_17035_p4 ^ tmp_660_fu_17021_p4);

assign xor_ln1545_487_fu_17553_p2 = (xor_ln1545_488_fu_17547_p2 ^ xor_ln1545_486_fu_17541_p2);

assign xor_ln1545_488_fu_17547_p2 = (trunc_ln674_164_fu_17099_p1 ^ tmp_667_fu_17079_p4);

assign xor_ln1545_489_fu_17559_p2 = (trunc_ln674_161_fu_16997_p1 ^ tmp_664_fu_17055_p4);

assign xor_ln1545_48_fu_5923_p2 = (trunc_ln674_14_fu_5569_p1 ^ tmp_77_fu_5549_p4);

assign xor_ln1545_490_fu_17571_p2 = (xor_ln1545_491_fu_17565_p2 ^ xor_ln1545_489_fu_17559_p2);

assign xor_ln1545_491_fu_17565_p2 = (tmp_671_fu_17113_p4 ^ tmp_666_fu_17069_p4);

assign xor_ln1545_492_fu_17577_p2 = (trunc_ln674_162_fu_17031_p1 ^ tmp_659_fu_17011_p4);

assign xor_ln1545_493_fu_17589_p2 = (xor_ln1545_494_fu_17583_p2 ^ xor_ln1545_492_fu_17577_p2);

assign xor_ln1545_494_fu_17583_p2 = (tmp_670_fu_17103_p4 ^ tmp_668_fu_17089_p4);

assign xor_ln1545_495_fu_17595_p2 = (tmp_663_fu_17045_p4 ^ tmp_658_fu_17001_p4);

assign xor_ln1545_496_fu_17601_p2 = (trunc_ln674_163_fu_17065_p1 ^ tmp_672_fu_17123_p4);

assign xor_ln1545_498_fu_17613_p2 = (tmp_678_fu_17171_p4 ^ tmp_676_fu_17157_p4);

assign xor_ln1545_499_fu_17625_p2 = (xor_ln1545_500_fu_17619_p2 ^ xor_ln1545_498_fu_17613_p2);

assign xor_ln1545_49_fu_5929_p2 = (tmp_88_fu_5641_p4 ^ tmp_86_fu_5627_p4);

assign xor_ln1545_500_fu_17619_p2 = (trunc_ln674_168_fu_17235_p1 ^ tmp_683_fu_17215_p4);

assign xor_ln1545_501_fu_17631_p2 = (trunc_ln674_165_fu_17133_p1 ^ tmp_680_fu_17191_p4);

assign xor_ln1545_502_fu_17643_p2 = (xor_ln1545_503_fu_17637_p2 ^ xor_ln1545_501_fu_17631_p2);

assign xor_ln1545_503_fu_17637_p2 = (tmp_687_fu_17249_p4 ^ tmp_682_fu_17205_p4);

assign xor_ln1545_504_fu_17649_p2 = (trunc_ln674_166_fu_17167_p1 ^ tmp_675_fu_17147_p4);

assign xor_ln1545_505_fu_17661_p2 = (xor_ln1545_506_fu_17655_p2 ^ xor_ln1545_504_fu_17649_p2);

assign xor_ln1545_506_fu_17655_p2 = (tmp_686_fu_17239_p4 ^ tmp_684_fu_17225_p4);

assign xor_ln1545_507_fu_17667_p2 = (tmp_679_fu_17181_p4 ^ tmp_674_fu_17137_p4);

assign xor_ln1545_508_fu_17679_p2 = (xor_ln1545_509_fu_17673_p2 ^ xor_ln1545_507_fu_17667_p2);

assign xor_ln1545_509_fu_17673_p2 = (trunc_ln674_167_fu_17201_p1 ^ tmp_688_fu_17259_p4);

assign xor_ln1545_510_fu_17685_p2 = (tmp_694_fu_17307_p4 ^ tmp_692_fu_17293_p4);

assign xor_ln1545_511_fu_17697_p2 = (xor_ln1545_512_fu_17691_p2 ^ xor_ln1545_510_fu_17685_p2);

assign xor_ln1545_512_fu_17691_p2 = (trunc_ln674_172_fu_17371_p1 ^ tmp_699_fu_17351_p4);

assign xor_ln1545_513_fu_17703_p2 = (trunc_ln674_169_fu_17269_p1 ^ tmp_696_fu_17327_p4);

assign xor_ln1545_514_fu_17715_p2 = (xor_ln1545_515_fu_17709_p2 ^ xor_ln1545_513_fu_17703_p2);

assign xor_ln1545_515_fu_17709_p2 = (tmp_703_fu_17385_p4 ^ tmp_698_fu_17341_p4);

assign xor_ln1545_516_fu_17721_p2 = (trunc_ln674_170_fu_17303_p1 ^ tmp_691_fu_17283_p4);

assign xor_ln1545_517_fu_17727_p2 = (tmp_702_fu_17375_p4 ^ tmp_700_fu_17361_p4);

assign xor_ln1545_519_fu_17739_p2 = (tmp_695_fu_17317_p4 ^ tmp_690_fu_17273_p4);

assign xor_ln1545_51_fu_5941_p2 = (tmp_81_fu_5583_p4 ^ tmp_76_fu_5539_p4);

assign xor_ln1545_520_fu_17751_p2 = (xor_ln1545_521_fu_17745_p2 ^ xor_ln1545_519_fu_17739_p2);

assign xor_ln1545_521_fu_17745_p2 = (trunc_ln674_171_fu_17337_p1 ^ tmp_704_fu_17395_p4);

assign xor_ln1545_522_fu_17757_p2 = (tmp_710_fu_17443_p4 ^ tmp_708_fu_17429_p4);

assign xor_ln1545_523_fu_17769_p2 = (xor_ln1545_524_fu_17763_p2 ^ xor_ln1545_522_fu_17757_p2);

assign xor_ln1545_524_fu_17763_p2 = (trunc_ln674_176_fu_17507_p1 ^ tmp_715_fu_17487_p4);

assign xor_ln1545_525_fu_17775_p2 = (trunc_ln674_173_fu_17405_p1 ^ tmp_712_fu_17463_p4);

assign xor_ln1545_526_fu_17781_p2 = (tmp_719_fu_17521_p4 ^ tmp_714_fu_17477_p4);

assign xor_ln1545_528_fu_17793_p2 = (trunc_ln674_174_fu_17439_p1 ^ tmp_707_fu_17419_p4);

assign xor_ln1545_529_fu_17799_p2 = (tmp_718_fu_17511_p4 ^ tmp_716_fu_17497_p4);

assign xor_ln1545_52_fu_5953_p2 = (xor_ln1545_53_fu_5947_p2 ^ xor_ln1545_51_fu_5941_p2);

assign xor_ln1545_531_fu_17811_p2 = (tmp_711_fu_17453_p4 ^ tmp_706_fu_17409_p4);

assign xor_ln1545_532_fu_17823_p2 = (xor_ln1545_533_fu_17817_p2 ^ xor_ln1545_531_fu_17811_p2);

assign xor_ln1545_533_fu_17817_p2 = (trunc_ln674_175_fu_17473_p1 ^ tmp_720_fu_17531_p4);

assign xor_ln1545_53_fu_5947_p2 = (trunc_ln674_15_fu_5603_p1 ^ tmp_90_fu_5661_p4);

assign xor_ln1545_54_fu_6858_p2 = (tmp_95_fu_6352_p4 ^ tmp_93_fu_6338_p4);

assign xor_ln1545_55_fu_6870_p2 = (xor_ln1545_56_fu_6864_p2 ^ xor_ln1545_54_fu_6858_p2);

assign xor_ln1545_56_fu_6864_p2 = (trunc_ln674_20_fu_6416_p1 ^ tmp_100_fu_6396_p4);

assign xor_ln1545_57_fu_6876_p2 = (trunc_ln674_17_fu_6314_p1 ^ tmp_97_fu_6372_p4);

assign xor_ln1545_58_fu_6888_p2 = (xor_ln1545_59_fu_6882_p2 ^ xor_ln1545_57_fu_6876_p2);

assign xor_ln1545_59_fu_6882_p2 = (tmp_99_fu_6386_p4 ^ tmp_104_fu_6430_p4);

assign xor_ln1545_60_fu_6894_p2 = (trunc_ln674_18_fu_6348_p1 ^ tmp_92_fu_6328_p4);

assign xor_ln1545_61_fu_6906_p2 = (xor_ln1545_62_fu_6900_p2 ^ xor_ln1545_60_fu_6894_p2);

assign xor_ln1545_62_fu_6900_p2 = (tmp_103_fu_6420_p4 ^ tmp_101_fu_6406_p4);

assign xor_ln1545_63_fu_6912_p2 = (tmp_96_fu_6362_p4 ^ tmp_91_fu_6318_p4);

assign xor_ln1545_64_fu_6918_p2 = (trunc_ln674_19_fu_6382_p1 ^ tmp_105_fu_6440_p4);

assign xor_ln1545_66_fu_6930_p2 = (tmp_111_fu_6488_p4 ^ tmp_109_fu_6474_p4);

assign xor_ln1545_67_fu_6942_p2 = (xor_ln1545_68_fu_6936_p2 ^ xor_ln1545_66_fu_6930_p2);

assign xor_ln1545_68_fu_6936_p2 = (trunc_ln674_24_fu_6552_p1 ^ tmp_116_fu_6532_p4);

assign xor_ln1545_69_fu_6948_p2 = (trunc_ln674_21_fu_6450_p1 ^ tmp_113_fu_6508_p4);

assign xor_ln1545_70_fu_6960_p2 = (xor_ln1545_71_fu_6954_p2 ^ xor_ln1545_69_fu_6948_p2);

assign xor_ln1545_71_fu_6954_p2 = (tmp_120_fu_6566_p4 ^ tmp_115_fu_6522_p4);

assign xor_ln1545_72_fu_6966_p2 = (trunc_ln674_22_fu_6484_p1 ^ tmp_108_fu_6464_p4);

assign xor_ln1545_73_fu_6978_p2 = (xor_ln1545_74_fu_6972_p2 ^ xor_ln1545_72_fu_6966_p2);

assign xor_ln1545_74_fu_6972_p2 = (tmp_119_fu_6556_p4 ^ tmp_117_fu_6542_p4);

assign xor_ln1545_75_fu_6984_p2 = (tmp_112_fu_6498_p4 ^ tmp_107_fu_6454_p4);

assign xor_ln1545_76_fu_6996_p2 = (xor_ln1545_77_fu_6990_p2 ^ xor_ln1545_75_fu_6984_p2);

assign xor_ln1545_77_fu_6990_p2 = (trunc_ln674_23_fu_6518_p1 ^ tmp_121_fu_6576_p4);

assign xor_ln1545_78_fu_7002_p2 = (tmp_127_fu_6624_p4 ^ tmp_125_fu_6610_p4);

assign xor_ln1545_79_fu_7014_p2 = (xor_ln1545_80_fu_7008_p2 ^ xor_ln1545_78_fu_7002_p2);

assign xor_ln1545_7_fu_5683_p2 = (xor_ln1545_fu_5671_p2 ^ xor_ln1545_8_fu_5677_p2);

assign xor_ln1545_80_fu_7008_p2 = (trunc_ln674_28_fu_6688_p1 ^ tmp_132_fu_6668_p4);

assign xor_ln1545_81_fu_7020_p2 = (trunc_ln674_25_fu_6586_p1 ^ tmp_129_fu_6644_p4);

assign xor_ln1545_82_fu_7032_p2 = (xor_ln1545_83_fu_7026_p2 ^ xor_ln1545_81_fu_7020_p2);

assign xor_ln1545_83_fu_7026_p2 = (tmp_136_fu_6702_p4 ^ tmp_131_fu_6658_p4);

assign xor_ln1545_84_fu_7038_p2 = (trunc_ln674_26_fu_6620_p1 ^ tmp_124_fu_6600_p4);

assign xor_ln1545_85_fu_7044_p2 = (tmp_135_fu_6692_p4 ^ tmp_133_fu_6678_p4);

assign xor_ln1545_87_fu_7056_p2 = (tmp_128_fu_6634_p4 ^ tmp_123_fu_6590_p4);

assign xor_ln1545_88_fu_7068_p2 = (xor_ln1545_89_fu_7062_p2 ^ xor_ln1545_87_fu_7056_p2);

assign xor_ln1545_89_fu_7062_p2 = (trunc_ln674_27_fu_6654_p1 ^ tmp_137_fu_6712_p4);

assign xor_ln1545_8_fu_5677_p2 = (trunc_ln674_4_fu_5229_p1 ^ tmp_37_fu_5209_p4);

assign xor_ln1545_90_fu_7074_p2 = (tmp_143_fu_6760_p4 ^ tmp_141_fu_6746_p4);

assign xor_ln1545_91_fu_7086_p2 = (xor_ln1545_92_fu_7080_p2 ^ xor_ln1545_90_fu_7074_p2);

assign xor_ln1545_92_fu_7080_p2 = (trunc_ln674_32_fu_6824_p1 ^ tmp_148_fu_6804_p4);

assign xor_ln1545_93_fu_7092_p2 = (trunc_ln674_29_fu_6722_p1 ^ tmp_145_fu_6780_p4);

assign xor_ln1545_94_fu_7098_p2 = (tmp_152_fu_6838_p4 ^ tmp_147_fu_6794_p4);

assign xor_ln1545_96_fu_7110_p2 = (trunc_ln674_30_fu_6756_p1 ^ tmp_140_fu_6736_p4);

assign xor_ln1545_97_fu_7116_p2 = (tmp_151_fu_6828_p4 ^ tmp_149_fu_6814_p4);

assign xor_ln1545_99_fu_7128_p2 = (tmp_144_fu_6770_p4 ^ tmp_139_fu_6726_p4);

assign xor_ln1545_9_fu_5689_p2 = (trunc_ln674_fu_5127_p1 ^ tmp_34_fu_5185_p4);

assign xor_ln1545_fu_5671_p2 = (tmp_32_fu_5165_p4 ^ tmp_30_fu_5151_p4);

assign zext_ln708_100_fu_8338_p1 = tmp_1_V_2_fu_8291_p2;

assign zext_ln708_101_fu_8343_p1 = tmp_2_1_V_2_fu_8237_p2;

assign zext_ln708_102_fu_8348_p1 = xor_ln1545_124_fu_8183_p2;

assign zext_ln708_103_fu_8353_p1 = xor_ln1545_115_fu_8129_p2;

assign zext_ln708_104_fu_8358_p1 = xor_ln1545_106_fu_8075_p2;

assign zext_ln708_105_fu_8363_p1 = tmp_2_2_V_2_fu_8309_p2;

assign zext_ln708_106_fu_8368_p1 = xor_ln1545_136_fu_8255_p2;

assign zext_ln708_107_fu_8373_p1 = xor_ln1545_127_fu_8201_p2;

assign zext_ln708_108_fu_8378_p1 = xor_ln1545_118_fu_8147_p2;

assign zext_ln708_109_fu_8383_p1 = xor_ln1545_109_fu_8093_p2;

assign zext_ln708_10_fu_4727_p1 = tmp_19_fu_4717_p4;

assign zext_ln708_110_fu_8388_p1 = xor_ln1545_148_fu_8327_p2;

assign zext_ln708_111_fu_8393_p1 = xor_ln1545_139_fu_8273_p2;

assign zext_ln708_112_fu_8398_p1 = xor_ln1545_130_fu_8219_p2;

assign zext_ln708_113_fu_8403_p1 = xor_ln1545_121_fu_8165_p2;

assign zext_ln708_114_fu_8408_p1 = tmp_3_V_2_fu_8111_p2;

assign zext_ln708_115_fu_8458_p1 = trunc_ln708_4_fu_8454_p1;

assign zext_ln708_116_fu_8473_p1 = tmp_220_fu_8463_p4;

assign zext_ln708_117_fu_8488_p1 = tmp_224_fu_8478_p4;

assign zext_ln708_118_fu_8503_p1 = tmp_228_fu_8493_p4;

assign zext_ln708_119_fu_8518_p1 = tmp_232_fu_8508_p4;

assign zext_ln708_11_fu_4742_p1 = tmp_20_fu_4732_p4;

assign zext_ln708_120_fu_8533_p1 = tmp_236_fu_8523_p4;

assign zext_ln708_121_fu_8548_p1 = tmp_240_fu_8538_p4;

assign zext_ln708_122_fu_8563_p1 = tmp_244_fu_8553_p4;

assign zext_ln708_123_fu_8578_p1 = tmp_248_fu_8568_p4;

assign zext_ln708_124_fu_8593_p1 = tmp_252_fu_8583_p4;

assign zext_ln708_125_fu_8608_p1 = tmp_256_fu_8598_p4;

assign zext_ln708_126_fu_8623_p1 = tmp_260_fu_8613_p4;

assign zext_ln708_127_fu_8638_p1 = tmp_264_fu_8628_p4;

assign zext_ln708_128_fu_8653_p1 = tmp_268_fu_8643_p4;

assign zext_ln708_129_fu_8668_p1 = tmp_272_fu_8658_p4;

assign zext_ln708_12_fu_4757_p1 = tmp_21_fu_4747_p4;

assign zext_ln708_130_fu_8683_p1 = tmp_276_fu_8673_p4;

assign zext_ln708_131_fu_9520_p1 = xor_ln1545_151_fu_9244_p2;

assign zext_ln708_132_fu_9525_p1 = tmp_1_V_3_fu_9478_p2;

assign zext_ln708_133_fu_9530_p1 = tmp_2_1_V_3_fu_9424_p2;

assign zext_ln708_134_fu_9535_p1 = xor_ln1545_172_fu_9370_p2;

assign zext_ln708_135_fu_9540_p1 = xor_ln1545_163_fu_9316_p2;

assign zext_ln708_136_fu_9545_p1 = xor_ln1545_154_fu_9262_p2;

assign zext_ln708_137_fu_9550_p1 = tmp_2_2_V_3_fu_9496_p2;

assign zext_ln708_138_fu_9555_p1 = xor_ln1545_184_fu_9442_p2;

assign zext_ln708_139_fu_9560_p1 = xor_ln1545_175_fu_9388_p2;

assign zext_ln708_13_fu_4772_p1 = tmp_22_fu_4762_p4;

assign zext_ln708_140_fu_9565_p1 = xor_ln1545_166_fu_9334_p2;

assign zext_ln708_141_fu_9570_p1 = xor_ln1545_157_fu_9280_p2;

assign zext_ln708_142_fu_9575_p1 = xor_ln1545_196_fu_9514_p2;

assign zext_ln708_143_fu_9580_p1 = xor_ln1545_187_fu_9460_p2;

assign zext_ln708_144_fu_9585_p1 = xor_ln1545_178_fu_9406_p2;

assign zext_ln708_145_fu_9590_p1 = xor_ln1545_169_fu_9352_p2;

assign zext_ln708_146_fu_9595_p1 = tmp_3_V_3_fu_9298_p2;

assign zext_ln708_147_fu_9645_p1 = trunc_ln708_5_fu_9641_p1;

assign zext_ln708_148_fu_9660_p1 = tmp_283_fu_9650_p4;

assign zext_ln708_149_fu_9675_p1 = tmp_287_fu_9665_p4;

assign zext_ln708_14_fu_4787_p1 = tmp_23_fu_4777_p4;

assign zext_ln708_150_fu_9690_p1 = tmp_291_fu_9680_p4;

assign zext_ln708_151_fu_9705_p1 = tmp_295_fu_9695_p4;

assign zext_ln708_152_fu_9720_p1 = tmp_299_fu_9710_p4;

assign zext_ln708_153_fu_9735_p1 = tmp_303_fu_9725_p4;

assign zext_ln708_154_fu_9750_p1 = tmp_307_fu_9740_p4;

assign zext_ln708_155_fu_9765_p1 = tmp_311_fu_9755_p4;

assign zext_ln708_156_fu_9780_p1 = tmp_315_fu_9770_p4;

assign zext_ln708_157_fu_9795_p1 = tmp_319_fu_9785_p4;

assign zext_ln708_158_fu_9810_p1 = tmp_323_fu_9800_p4;

assign zext_ln708_159_fu_9825_p1 = tmp_327_fu_9815_p4;

assign zext_ln708_15_fu_4802_p1 = tmp_24_fu_4792_p4;

assign zext_ln708_160_fu_9840_p1 = tmp_331_fu_9830_p4;

assign zext_ln708_161_fu_9855_p1 = tmp_335_fu_9845_p4;

assign zext_ln708_162_fu_9870_p1 = tmp_339_fu_9860_p4;

assign zext_ln708_163_fu_10707_p1 = xor_ln1545_199_fu_10431_p2;

assign zext_ln708_164_fu_10712_p1 = tmp_1_V_4_fu_10665_p2;

assign zext_ln708_165_fu_10717_p1 = tmp_2_1_V_4_fu_10611_p2;

assign zext_ln708_166_fu_10722_p1 = xor_ln1545_220_fu_10557_p2;

assign zext_ln708_167_fu_10727_p1 = xor_ln1545_211_fu_10503_p2;

assign zext_ln708_168_fu_10732_p1 = xor_ln1545_202_fu_10449_p2;

assign zext_ln708_169_fu_10737_p1 = tmp_2_2_V_4_fu_10683_p2;

assign zext_ln708_16_fu_4817_p1 = tmp_25_fu_4807_p4;

assign zext_ln708_170_fu_10742_p1 = xor_ln1545_232_fu_10629_p2;

assign zext_ln708_171_fu_10747_p1 = xor_ln1545_223_fu_10575_p2;

assign zext_ln708_172_fu_10752_p1 = xor_ln1545_214_fu_10521_p2;

assign zext_ln708_173_fu_10757_p1 = xor_ln1545_205_fu_10467_p2;

assign zext_ln708_174_fu_10762_p1 = xor_ln1545_244_fu_10701_p2;

assign zext_ln708_175_fu_10767_p1 = xor_ln1545_235_fu_10647_p2;

assign zext_ln708_176_fu_10772_p1 = xor_ln1545_226_fu_10593_p2;

assign zext_ln708_177_fu_10777_p1 = xor_ln1545_217_fu_10539_p2;

assign zext_ln708_178_fu_10782_p1 = tmp_3_V_4_fu_10485_p2;

assign zext_ln708_179_fu_10832_p1 = trunc_ln708_6_fu_10828_p1;

assign zext_ln708_17_fu_4832_p1 = tmp_26_fu_4822_p4;

assign zext_ln708_180_fu_10847_p1 = tmp_346_fu_10837_p4;

assign zext_ln708_181_fu_10862_p1 = tmp_350_fu_10852_p4;

assign zext_ln708_182_fu_10877_p1 = tmp_354_fu_10867_p4;

assign zext_ln708_183_fu_10892_p1 = tmp_358_fu_10882_p4;

assign zext_ln708_184_fu_10907_p1 = tmp_362_fu_10897_p4;

assign zext_ln708_185_fu_10922_p1 = tmp_366_fu_10912_p4;

assign zext_ln708_186_fu_10937_p1 = tmp_370_fu_10927_p4;

assign zext_ln708_187_fu_10952_p1 = tmp_374_fu_10942_p4;

assign zext_ln708_188_fu_10967_p1 = tmp_378_fu_10957_p4;

assign zext_ln708_189_fu_10982_p1 = tmp_382_fu_10972_p4;

assign zext_ln708_18_fu_4847_p1 = tmp_27_fu_4837_p4;

assign zext_ln708_190_fu_10997_p1 = tmp_386_fu_10987_p4;

assign zext_ln708_191_fu_11012_p1 = tmp_390_fu_11002_p4;

assign zext_ln708_192_fu_11027_p1 = tmp_394_fu_11017_p4;

assign zext_ln708_193_fu_11042_p1 = tmp_398_fu_11032_p4;

assign zext_ln708_194_fu_11057_p1 = tmp_402_fu_11047_p4;

assign zext_ln708_195_fu_11894_p1 = xor_ln1545_247_fu_11618_p2;

assign zext_ln708_196_fu_11899_p1 = tmp_1_V_5_fu_11852_p2;

assign zext_ln708_197_fu_11904_p1 = tmp_2_1_V_5_fu_11798_p2;

assign zext_ln708_198_fu_11909_p1 = xor_ln1545_268_fu_11744_p2;

assign zext_ln708_199_fu_11914_p1 = xor_ln1545_259_fu_11690_p2;

assign zext_ln708_19_fu_4897_p1 = trunc_ln708_1_fu_4893_p1;

assign zext_ln708_200_fu_11919_p1 = xor_ln1545_250_fu_11636_p2;

assign zext_ln708_201_fu_11924_p1 = tmp_2_2_V_5_fu_11870_p2;

assign zext_ln708_202_fu_11929_p1 = xor_ln1545_280_fu_11816_p2;

assign zext_ln708_203_fu_11934_p1 = xor_ln1545_271_fu_11762_p2;

assign zext_ln708_204_fu_11939_p1 = xor_ln1545_262_fu_11708_p2;

assign zext_ln708_205_fu_11944_p1 = xor_ln1545_253_fu_11654_p2;

assign zext_ln708_206_fu_11949_p1 = xor_ln1545_292_fu_11888_p2;

assign zext_ln708_207_fu_11954_p1 = xor_ln1545_283_fu_11834_p2;

assign zext_ln708_208_fu_11959_p1 = xor_ln1545_274_fu_11780_p2;

assign zext_ln708_209_fu_11964_p1 = xor_ln1545_265_fu_11726_p2;

assign zext_ln708_20_fu_4912_p1 = tmp_31_fu_4902_p4;

assign zext_ln708_210_fu_11969_p1 = tmp_3_V_5_fu_11672_p2;

assign zext_ln708_211_fu_12019_p1 = trunc_ln708_7_fu_12015_p1;

assign zext_ln708_212_fu_12034_p1 = tmp_409_fu_12024_p4;

assign zext_ln708_213_fu_12049_p1 = tmp_413_fu_12039_p4;

assign zext_ln708_214_fu_12064_p1 = tmp_417_fu_12054_p4;

assign zext_ln708_215_fu_12079_p1 = tmp_421_fu_12069_p4;

assign zext_ln708_216_fu_12094_p1 = tmp_425_fu_12084_p4;

assign zext_ln708_217_fu_12109_p1 = tmp_429_fu_12099_p4;

assign zext_ln708_218_fu_12124_p1 = tmp_433_fu_12114_p4;

assign zext_ln708_219_fu_12139_p1 = tmp_437_fu_12129_p4;

assign zext_ln708_21_fu_4927_p1 = tmp_35_fu_4917_p4;

assign zext_ln708_220_fu_12154_p1 = tmp_441_fu_12144_p4;

assign zext_ln708_221_fu_12169_p1 = tmp_445_fu_12159_p4;

assign zext_ln708_222_fu_12184_p1 = tmp_449_fu_12174_p4;

assign zext_ln708_223_fu_12199_p1 = tmp_453_fu_12189_p4;

assign zext_ln708_224_fu_12214_p1 = tmp_457_fu_12204_p4;

assign zext_ln708_225_fu_12229_p1 = tmp_461_fu_12219_p4;

assign zext_ln708_226_fu_12244_p1 = tmp_465_fu_12234_p4;

assign zext_ln708_227_fu_13081_p1 = xor_ln1545_295_fu_12805_p2;

assign zext_ln708_228_fu_13086_p1 = tmp_1_V_6_fu_13039_p2;

assign zext_ln708_229_fu_13091_p1 = tmp_2_1_V_6_fu_12985_p2;

assign zext_ln708_22_fu_4942_p1 = tmp_39_fu_4932_p4;

assign zext_ln708_230_fu_13096_p1 = xor_ln1545_316_fu_12931_p2;

assign zext_ln708_231_fu_13101_p1 = xor_ln1545_307_fu_12877_p2;

assign zext_ln708_232_fu_13106_p1 = xor_ln1545_298_fu_12823_p2;

assign zext_ln708_233_fu_13111_p1 = tmp_2_2_V_6_fu_13057_p2;

assign zext_ln708_234_fu_13116_p1 = xor_ln1545_328_fu_13003_p2;

assign zext_ln708_235_fu_13121_p1 = xor_ln1545_319_fu_12949_p2;

assign zext_ln708_236_fu_13126_p1 = xor_ln1545_310_fu_12895_p2;

assign zext_ln708_237_fu_13131_p1 = xor_ln1545_301_fu_12841_p2;

assign zext_ln708_238_fu_13136_p1 = xor_ln1545_340_fu_13075_p2;

assign zext_ln708_239_fu_13141_p1 = xor_ln1545_331_fu_13021_p2;

assign zext_ln708_23_fu_4957_p1 = tmp_43_fu_4947_p4;

assign zext_ln708_240_fu_13146_p1 = xor_ln1545_322_fu_12967_p2;

assign zext_ln708_241_fu_13151_p1 = xor_ln1545_313_fu_12913_p2;

assign zext_ln708_242_fu_13156_p1 = tmp_3_V_6_fu_12859_p2;

assign zext_ln708_243_fu_13206_p1 = trunc_ln708_8_fu_13202_p1;

assign zext_ln708_244_fu_13221_p1 = tmp_472_fu_13211_p4;

assign zext_ln708_245_fu_13236_p1 = tmp_476_fu_13226_p4;

assign zext_ln708_246_fu_13251_p1 = tmp_480_fu_13241_p4;

assign zext_ln708_247_fu_13266_p1 = tmp_484_fu_13256_p4;

assign zext_ln708_248_fu_13281_p1 = tmp_488_fu_13271_p4;

assign zext_ln708_249_fu_13296_p1 = tmp_492_fu_13286_p4;

assign zext_ln708_24_fu_4972_p1 = tmp_47_fu_4962_p4;

assign zext_ln708_250_fu_13311_p1 = tmp_496_fu_13301_p4;

assign zext_ln708_251_fu_13326_p1 = tmp_500_fu_13316_p4;

assign zext_ln708_252_fu_13341_p1 = tmp_504_fu_13331_p4;

assign zext_ln708_253_fu_13356_p1 = tmp_508_fu_13346_p4;

assign zext_ln708_254_fu_13371_p1 = tmp_512_fu_13361_p4;

assign zext_ln708_255_fu_13386_p1 = tmp_516_fu_13376_p4;

assign zext_ln708_256_fu_13401_p1 = tmp_520_fu_13391_p4;

assign zext_ln708_257_fu_13416_p1 = tmp_524_fu_13406_p4;

assign zext_ln708_258_fu_13431_p1 = tmp_528_fu_13421_p4;

assign zext_ln708_259_fu_14268_p1 = xor_ln1545_343_fu_13992_p2;

assign zext_ln708_25_fu_4987_p1 = tmp_51_fu_4977_p4;

assign zext_ln708_260_fu_14273_p1 = tmp_1_V_7_fu_14226_p2;

assign zext_ln708_261_fu_14278_p1 = tmp_2_1_V_7_fu_14172_p2;

assign zext_ln708_262_fu_14283_p1 = xor_ln1545_364_fu_14118_p2;

assign zext_ln708_263_fu_14288_p1 = xor_ln1545_355_fu_14064_p2;

assign zext_ln708_264_fu_14293_p1 = xor_ln1545_346_fu_14010_p2;

assign zext_ln708_265_fu_14298_p1 = tmp_2_2_V_7_fu_14244_p2;

assign zext_ln708_266_fu_14303_p1 = xor_ln1545_376_fu_14190_p2;

assign zext_ln708_267_fu_14308_p1 = xor_ln1545_367_fu_14136_p2;

assign zext_ln708_268_fu_14313_p1 = xor_ln1545_358_fu_14082_p2;

assign zext_ln708_269_fu_14318_p1 = xor_ln1545_349_fu_14028_p2;

assign zext_ln708_26_fu_5002_p1 = tmp_55_fu_4992_p4;

assign zext_ln708_270_fu_14323_p1 = xor_ln1545_388_fu_14262_p2;

assign zext_ln708_271_fu_14328_p1 = xor_ln1545_379_fu_14208_p2;

assign zext_ln708_272_fu_14333_p1 = xor_ln1545_370_fu_14154_p2;

assign zext_ln708_273_fu_14338_p1 = xor_ln1545_361_fu_14100_p2;

assign zext_ln708_274_fu_14343_p1 = tmp_3_V_7_fu_14046_p2;

assign zext_ln708_275_fu_14393_p1 = trunc_ln708_9_fu_14389_p1;

assign zext_ln708_276_fu_14408_p1 = tmp_535_fu_14398_p4;

assign zext_ln708_277_fu_14423_p1 = tmp_539_fu_14413_p4;

assign zext_ln708_278_fu_14438_p1 = tmp_543_fu_14428_p4;

assign zext_ln708_279_fu_14453_p1 = tmp_547_fu_14443_p4;

assign zext_ln708_27_fu_5017_p1 = tmp_59_fu_5007_p4;

assign zext_ln708_280_fu_14468_p1 = tmp_551_fu_14458_p4;

assign zext_ln708_281_fu_14483_p1 = tmp_555_fu_14473_p4;

assign zext_ln708_282_fu_14498_p1 = tmp_559_fu_14488_p4;

assign zext_ln708_283_fu_14513_p1 = tmp_563_fu_14503_p4;

assign zext_ln708_284_fu_14528_p1 = tmp_567_fu_14518_p4;

assign zext_ln708_285_fu_14543_p1 = tmp_571_fu_14533_p4;

assign zext_ln708_286_fu_14558_p1 = tmp_575_fu_14548_p4;

assign zext_ln708_287_fu_14573_p1 = tmp_579_fu_14563_p4;

assign zext_ln708_288_fu_14588_p1 = tmp_583_fu_14578_p4;

assign zext_ln708_289_fu_14603_p1 = tmp_587_fu_14593_p4;

assign zext_ln708_28_fu_5032_p1 = tmp_63_fu_5022_p4;

assign zext_ln708_290_fu_14618_p1 = tmp_591_fu_14608_p4;

assign zext_ln708_291_fu_15455_p1 = xor_ln1545_391_fu_15179_p2;

assign zext_ln708_292_fu_15460_p1 = tmp_1_V_8_fu_15413_p2;

assign zext_ln708_293_fu_15465_p1 = tmp_2_1_V_8_fu_15359_p2;

assign zext_ln708_294_fu_15470_p1 = xor_ln1545_412_fu_15305_p2;

assign zext_ln708_295_fu_15475_p1 = xor_ln1545_403_fu_15251_p2;

assign zext_ln708_296_fu_15480_p1 = xor_ln1545_394_fu_15197_p2;

assign zext_ln708_297_fu_15485_p1 = tmp_2_2_V_8_fu_15431_p2;

assign zext_ln708_298_fu_15490_p1 = xor_ln1545_424_fu_15377_p2;

assign zext_ln708_299_fu_15495_p1 = xor_ln1545_415_fu_15323_p2;

assign zext_ln708_29_fu_5047_p1 = tmp_67_fu_5037_p4;

assign zext_ln708_300_fu_15500_p1 = xor_ln1545_406_fu_15269_p2;

assign zext_ln708_301_fu_15505_p1 = xor_ln1545_397_fu_15215_p2;

assign zext_ln708_302_fu_15510_p1 = xor_ln1545_436_fu_15449_p2;

assign zext_ln708_303_fu_15515_p1 = xor_ln1545_427_fu_15395_p2;

assign zext_ln708_304_fu_15520_p1 = xor_ln1545_418_fu_15341_p2;

assign zext_ln708_305_fu_15525_p1 = xor_ln1545_409_fu_15287_p2;

assign zext_ln708_306_fu_15530_p1 = tmp_3_V_8_fu_15233_p2;

assign zext_ln708_307_fu_15580_p1 = trunc_ln708_10_fu_15576_p1;

assign zext_ln708_308_fu_15595_p1 = tmp_598_fu_15585_p4;

assign zext_ln708_309_fu_15610_p1 = tmp_602_fu_15600_p4;

assign zext_ln708_30_fu_5062_p1 = tmp_71_fu_5052_p4;

assign zext_ln708_310_fu_15625_p1 = tmp_606_fu_15615_p4;

assign zext_ln708_311_fu_15640_p1 = tmp_610_fu_15630_p4;

assign zext_ln708_312_fu_15655_p1 = tmp_614_fu_15645_p4;

assign zext_ln708_313_fu_15670_p1 = tmp_618_fu_15660_p4;

assign zext_ln708_314_fu_15685_p1 = tmp_622_fu_15675_p4;

assign zext_ln708_315_fu_15700_p1 = tmp_626_fu_15690_p4;

assign zext_ln708_316_fu_15715_p1 = tmp_630_fu_15705_p4;

assign zext_ln708_317_fu_15730_p1 = tmp_634_fu_15720_p4;

assign zext_ln708_318_fu_15745_p1 = tmp_638_fu_15735_p4;

assign zext_ln708_319_fu_15760_p1 = tmp_642_fu_15750_p4;

assign zext_ln708_31_fu_5077_p1 = tmp_75_fu_5067_p4;

assign zext_ln708_320_fu_15775_p1 = tmp_646_fu_15765_p4;

assign zext_ln708_321_fu_15790_p1 = tmp_650_fu_15780_p4;

assign zext_ln708_322_fu_15805_p1 = tmp_654_fu_15795_p4;

assign zext_ln708_323_fu_16642_p1 = xor_ln1545_439_fu_16366_p2;

assign zext_ln708_324_fu_16647_p1 = tmp_1_V_9_fu_16600_p2;

assign zext_ln708_325_fu_16652_p1 = tmp_2_1_V_9_fu_16546_p2;

assign zext_ln708_326_fu_16657_p1 = xor_ln1545_460_fu_16492_p2;

assign zext_ln708_327_fu_16662_p1 = xor_ln1545_451_fu_16438_p2;

assign zext_ln708_328_fu_16667_p1 = xor_ln1545_442_fu_16384_p2;

assign zext_ln708_329_fu_16672_p1 = tmp_2_2_V_9_fu_16618_p2;

assign zext_ln708_32_fu_5092_p1 = tmp_79_fu_5082_p4;

assign zext_ln708_330_fu_16677_p1 = xor_ln1545_472_fu_16564_p2;

assign zext_ln708_331_fu_16682_p1 = xor_ln1545_463_fu_16510_p2;

assign zext_ln708_332_fu_16687_p1 = xor_ln1545_454_fu_16456_p2;

assign zext_ln708_333_fu_16692_p1 = xor_ln1545_445_fu_16402_p2;

assign zext_ln708_334_fu_16697_p1 = xor_ln1545_484_fu_16636_p2;

assign zext_ln708_335_fu_16702_p1 = xor_ln1545_475_fu_16582_p2;

assign zext_ln708_336_fu_16707_p1 = xor_ln1545_466_fu_16528_p2;

assign zext_ln708_337_fu_16712_p1 = xor_ln1545_457_fu_16474_p2;

assign zext_ln708_338_fu_16717_p1 = tmp_3_V_9_fu_16420_p2;

assign zext_ln708_339_fu_16767_p1 = trunc_ln708_11_fu_16763_p1;

assign zext_ln708_33_fu_5107_p1 = tmp_83_fu_5097_p4;

assign zext_ln708_340_fu_16782_p1 = tmp_661_fu_16772_p4;

assign zext_ln708_341_fu_16797_p1 = tmp_665_fu_16787_p4;

assign zext_ln708_342_fu_16812_p1 = tmp_669_fu_16802_p4;

assign zext_ln708_343_fu_16827_p1 = tmp_673_fu_16817_p4;

assign zext_ln708_344_fu_16842_p1 = tmp_677_fu_16832_p4;

assign zext_ln708_345_fu_16857_p1 = tmp_681_fu_16847_p4;

assign zext_ln708_346_fu_16872_p1 = tmp_685_fu_16862_p4;

assign zext_ln708_347_fu_16887_p1 = tmp_689_fu_16877_p4;

assign zext_ln708_348_fu_16902_p1 = tmp_693_fu_16892_p4;

assign zext_ln708_349_fu_16917_p1 = tmp_697_fu_16907_p4;

assign zext_ln708_34_fu_5122_p1 = tmp_87_fu_5112_p4;

assign zext_ln708_350_fu_16932_p1 = tmp_701_fu_16922_p4;

assign zext_ln708_351_fu_16947_p1 = tmp_705_fu_16937_p4;

assign zext_ln708_352_fu_16962_p1 = tmp_709_fu_16952_p4;

assign zext_ln708_353_fu_16977_p1 = tmp_713_fu_16967_p4;

assign zext_ln708_354_fu_16992_p1 = tmp_717_fu_16982_p4;

assign zext_ln708_355_fu_17829_p1 = xor_ln1545_487_fu_17553_p2;

assign zext_ln708_356_fu_17834_p1 = tmp_1_V_10_fu_17787_p2;

assign zext_ln708_357_fu_17839_p1 = tmp_2_1_V_10_fu_17733_p2;

assign zext_ln708_358_fu_17844_p1 = xor_ln1545_508_fu_17679_p2;

assign zext_ln708_359_fu_17849_p1 = xor_ln1545_499_fu_17625_p2;

assign zext_ln708_35_fu_5959_p1 = xor_ln1545_7_fu_5683_p2;

assign zext_ln708_360_fu_17854_p1 = xor_ln1545_490_fu_17571_p2;

assign zext_ln708_361_fu_17859_p1 = tmp_2_2_V_10_fu_17805_p2;

assign zext_ln708_362_fu_17864_p1 = xor_ln1545_520_fu_17751_p2;

assign zext_ln708_363_fu_17869_p1 = xor_ln1545_511_fu_17697_p2;

assign zext_ln708_364_fu_17874_p1 = xor_ln1545_502_fu_17643_p2;

assign zext_ln708_365_fu_17879_p1 = xor_ln1545_493_fu_17589_p2;

assign zext_ln708_366_fu_17884_p1 = xor_ln1545_532_fu_17823_p2;

assign zext_ln708_367_fu_17889_p1 = xor_ln1545_523_fu_17769_p2;

assign zext_ln708_368_fu_17894_p1 = xor_ln1545_514_fu_17715_p2;

assign zext_ln708_369_fu_17899_p1 = xor_ln1545_505_fu_17661_p2;

assign zext_ln708_36_fu_5964_p1 = tmp_1_V_fu_5917_p2;

assign zext_ln708_370_fu_17904_p1 = tmp_3_V_10_fu_17607_p2;

assign zext_ln708_37_fu_5969_p1 = tmp_2_1_V_fu_5863_p2;

assign zext_ln708_38_fu_5974_p1 = xor_ln1545_28_fu_5809_p2;

assign zext_ln708_39_fu_5979_p1 = xor_ln1545_19_fu_5755_p2;

assign zext_ln708_40_fu_5984_p1 = xor_ln1545_10_fu_5701_p2;

assign zext_ln708_41_fu_5989_p1 = tmp_2_2_V_fu_5935_p2;

assign zext_ln708_42_fu_5994_p1 = xor_ln1545_40_fu_5881_p2;

assign zext_ln708_43_fu_5999_p1 = xor_ln1545_31_fu_5827_p2;

assign zext_ln708_44_fu_6004_p1 = xor_ln1545_22_fu_5773_p2;

assign zext_ln708_45_fu_6009_p1 = xor_ln1545_13_fu_5719_p2;

assign zext_ln708_46_fu_6014_p1 = xor_ln1545_52_fu_5953_p2;

assign zext_ln708_47_fu_6019_p1 = xor_ln1545_43_fu_5899_p2;

assign zext_ln708_48_fu_6024_p1 = xor_ln1545_34_fu_5845_p2;

assign zext_ln708_49_fu_6029_p1 = xor_ln1545_25_fu_5791_p2;

assign zext_ln708_4_fu_4637_p1 = tmp_s_fu_4627_p4;

assign zext_ln708_50_fu_6034_p1 = tmp_3_V_fu_5737_p2;

assign zext_ln708_51_fu_6084_p1 = trunc_ln708_2_fu_6080_p1;

assign zext_ln708_52_fu_6099_p1 = tmp_94_fu_6089_p4;

assign zext_ln708_53_fu_6114_p1 = tmp_98_fu_6104_p4;

assign zext_ln708_54_fu_6129_p1 = tmp_102_fu_6119_p4;

assign zext_ln708_55_fu_6144_p1 = tmp_106_fu_6134_p4;

assign zext_ln708_56_fu_6159_p1 = tmp_110_fu_6149_p4;

assign zext_ln708_57_fu_6174_p1 = tmp_114_fu_6164_p4;

assign zext_ln708_58_fu_6189_p1 = tmp_118_fu_6179_p4;

assign zext_ln708_59_fu_6204_p1 = tmp_122_fu_6194_p4;

assign zext_ln708_5_fu_4652_p1 = tmp_14_fu_4642_p4;

assign zext_ln708_60_fu_6219_p1 = tmp_126_fu_6209_p4;

assign zext_ln708_61_fu_6234_p1 = tmp_130_fu_6224_p4;

assign zext_ln708_62_fu_6249_p1 = tmp_134_fu_6239_p4;

assign zext_ln708_63_fu_6264_p1 = tmp_138_fu_6254_p4;

assign zext_ln708_64_fu_6279_p1 = tmp_142_fu_6269_p4;

assign zext_ln708_65_fu_6294_p1 = tmp_146_fu_6284_p4;

assign zext_ln708_66_fu_6309_p1 = tmp_150_fu_6299_p4;

assign zext_ln708_67_fu_7146_p1 = xor_ln1545_55_fu_6870_p2;

assign zext_ln708_68_fu_7151_p1 = tmp_1_V_1_fu_7104_p2;

assign zext_ln708_69_fu_7156_p1 = tmp_2_1_V_1_fu_7050_p2;

assign zext_ln708_6_fu_4667_p1 = tmp_15_fu_4657_p4;

assign zext_ln708_70_fu_7161_p1 = xor_ln1545_76_fu_6996_p2;

assign zext_ln708_71_fu_7166_p1 = xor_ln1545_67_fu_6942_p2;

assign zext_ln708_72_fu_7171_p1 = xor_ln1545_58_fu_6888_p2;

assign zext_ln708_73_fu_7176_p1 = tmp_2_2_V_1_fu_7122_p2;

assign zext_ln708_74_fu_7181_p1 = xor_ln1545_88_fu_7068_p2;

assign zext_ln708_75_fu_7186_p1 = xor_ln1545_79_fu_7014_p2;

assign zext_ln708_76_fu_7191_p1 = xor_ln1545_70_fu_6960_p2;

assign zext_ln708_77_fu_7196_p1 = xor_ln1545_61_fu_6906_p2;

assign zext_ln708_78_fu_7201_p1 = xor_ln1545_100_fu_7140_p2;

assign zext_ln708_79_fu_7206_p1 = xor_ln1545_91_fu_7086_p2;

assign zext_ln708_7_fu_4682_p1 = tmp_16_fu_4672_p4;

assign zext_ln708_80_fu_7211_p1 = xor_ln1545_82_fu_7032_p2;

assign zext_ln708_81_fu_7216_p1 = xor_ln1545_73_fu_6978_p2;

assign zext_ln708_82_fu_7221_p1 = tmp_3_V_1_fu_6924_p2;

assign zext_ln708_83_fu_7271_p1 = trunc_ln708_3_fu_7267_p1;

assign zext_ln708_84_fu_7286_p1 = tmp_157_fu_7276_p4;

assign zext_ln708_85_fu_7301_p1 = tmp_161_fu_7291_p4;

assign zext_ln708_86_fu_7316_p1 = tmp_165_fu_7306_p4;

assign zext_ln708_87_fu_7331_p1 = tmp_169_fu_7321_p4;

assign zext_ln708_88_fu_7346_p1 = tmp_173_fu_7336_p4;

assign zext_ln708_89_fu_7361_p1 = tmp_177_fu_7351_p4;

assign zext_ln708_8_fu_4697_p1 = tmp_17_fu_4687_p4;

assign zext_ln708_90_fu_7376_p1 = tmp_181_fu_7366_p4;

assign zext_ln708_91_fu_7391_p1 = tmp_185_fu_7381_p4;

assign zext_ln708_92_fu_7406_p1 = tmp_189_fu_7396_p4;

assign zext_ln708_93_fu_7421_p1 = tmp_193_fu_7411_p4;

assign zext_ln708_94_fu_7436_p1 = tmp_197_fu_7426_p4;

assign zext_ln708_95_fu_7451_p1 = tmp_201_fu_7441_p4;

assign zext_ln708_96_fu_7466_p1 = tmp_205_fu_7456_p4;

assign zext_ln708_97_fu_7481_p1 = tmp_209_fu_7471_p4;

assign zext_ln708_98_fu_7496_p1 = tmp_213_fu_7486_p4;

assign zext_ln708_99_fu_8333_p1 = xor_ln1545_103_fu_8057_p2;

assign zext_ln708_9_fu_4712_p1 = tmp_18_fu_4702_p4;

assign zext_ln708_fu_4622_p1 = trunc_ln708_fu_4618_p1;

endmodule //testDec_process_r
