// Copyright (C) 2022, Advanced Micro Devices, Inc. All rights reserved.
// SPDX-License-Identifier: MIT
// ==============================================================
// Version: 2022.1.0
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module testDec_process_r (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        p_read,
        p_read1,
        p_read2,
        p_read3,
        p_read4,
        p_read5,
        p_read6,
        p_read7,
        p_read8,
        p_read9,
        p_read10,
        ciphertext,
        ap_return
);

parameter    ap_ST_fsm_pp0_stage0 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [127:0] p_read;
input  [127:0] p_read1;
input  [127:0] p_read2;
input  [127:0] p_read3;
input  [127:0] p_read4;
input  [127:0] p_read5;
input  [127:0] p_read6;
input  [127:0] p_read7;
input  [127:0] p_read8;
input  [127:0] p_read9;
input  [127:0] p_read10;
input  [127:0] ciphertext;
output  [127:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;

(* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg    ap_enable_reg_pp0_iter5;
reg    ap_enable_reg_pp0_iter6;
reg    ap_enable_reg_pp0_iter7;
reg    ap_enable_reg_pp0_iter8;
reg    ap_enable_reg_pp0_iter9;
reg    ap_enable_reg_pp0_iter10;
reg    ap_enable_reg_pp0_iter11;
reg    ap_enable_reg_pp0_iter12;
reg    ap_enable_reg_pp0_iter13;
reg    ap_enable_reg_pp0_iter14;
reg    ap_enable_reg_pp0_iter15;
reg    ap_enable_reg_pp0_iter16;
reg    ap_enable_reg_pp0_iter17;
reg    ap_enable_reg_pp0_iter18;
reg    ap_enable_reg_pp0_iter19;
reg    ap_idle_pp0;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_state4_pp0_stage0_iter3;
wire    ap_block_state5_pp0_stage0_iter4;
wire    ap_block_state6_pp0_stage0_iter5;
wire    ap_block_state7_pp0_stage0_iter6;
wire    ap_block_state8_pp0_stage0_iter7;
wire    ap_block_state9_pp0_stage0_iter8;
wire    ap_block_state10_pp0_stage0_iter9;
wire    ap_block_state11_pp0_stage0_iter10;
wire    ap_block_state12_pp0_stage0_iter11;
wire    ap_block_state13_pp0_stage0_iter12;
wire    ap_block_state14_pp0_stage0_iter13;
wire    ap_block_state15_pp0_stage0_iter14;
wire    ap_block_state16_pp0_stage0_iter15;
wire    ap_block_state17_pp0_stage0_iter16;
wire    ap_block_state18_pp0_stage0_iter17;
wire    ap_block_state19_pp0_stage0_iter18;
wire    ap_block_state20_pp0_stage0_iter19;
wire    ap_block_pp0_stage0_subdone;
wire   [7:0] decipher_0_iibox_address0;
reg    decipher_0_iibox_ce0;
wire   [7:0] decipher_0_iibox_q0;
wire   [7:0] decipher_0_iibox_address1;
reg    decipher_0_iibox_ce1;
wire   [7:0] decipher_0_iibox_q1;
wire   [7:0] decipher_0_iibox_address2;
reg    decipher_0_iibox_ce2;
wire   [7:0] decipher_0_iibox_q2;
wire   [7:0] decipher_0_iibox_address3;
reg    decipher_0_iibox_ce3;
wire   [7:0] decipher_0_iibox_q3;
wire   [7:0] decipher_0_iibox_address4;
reg    decipher_0_iibox_ce4;
wire   [7:0] decipher_0_iibox_q4;
wire   [7:0] decipher_0_iibox_address5;
reg    decipher_0_iibox_ce5;
wire   [7:0] decipher_0_iibox_q5;
wire   [7:0] decipher_0_iibox_address6;
reg    decipher_0_iibox_ce6;
wire   [7:0] decipher_0_iibox_q6;
wire   [7:0] decipher_0_iibox_address7;
reg    decipher_0_iibox_ce7;
wire   [7:0] decipher_0_iibox_q7;
wire   [7:0] decipher_0_iibox_address8;
reg    decipher_0_iibox_ce8;
wire   [7:0] decipher_0_iibox_q8;
wire   [7:0] decipher_0_iibox_address9;
reg    decipher_0_iibox_ce9;
wire   [7:0] decipher_0_iibox_q9;
wire   [7:0] decipher_0_iibox_address10;
reg    decipher_0_iibox_ce10;
wire   [7:0] decipher_0_iibox_q10;
wire   [7:0] decipher_0_iibox_address11;
reg    decipher_0_iibox_ce11;
wire   [7:0] decipher_0_iibox_q11;
wire   [7:0] decipher_0_iibox_address12;
reg    decipher_0_iibox_ce12;
wire   [7:0] decipher_0_iibox_q12;
wire   [7:0] decipher_0_iibox_address13;
reg    decipher_0_iibox_ce13;
wire   [7:0] decipher_0_iibox_q13;
wire   [7:0] decipher_0_iibox_address14;
reg    decipher_0_iibox_ce14;
wire   [7:0] decipher_0_iibox_q14;
wire   [7:0] decipher_0_iibox_address15;
reg    decipher_0_iibox_ce15;
wire   [7:0] decipher_0_iibox_q15;
wire   [7:0] decipher_0_iibox_address16;
reg    decipher_0_iibox_ce16;
wire   [7:0] decipher_0_iibox_q16;
wire   [7:0] decipher_0_iibox_address17;
reg    decipher_0_iibox_ce17;
wire   [7:0] decipher_0_iibox_q17;
wire   [7:0] decipher_0_iibox_address18;
reg    decipher_0_iibox_ce18;
wire   [7:0] decipher_0_iibox_q18;
wire   [7:0] decipher_0_iibox_address19;
reg    decipher_0_iibox_ce19;
wire   [7:0] decipher_0_iibox_q19;
wire   [7:0] decipher_0_iibox_address20;
reg    decipher_0_iibox_ce20;
wire   [7:0] decipher_0_iibox_q20;
wire   [7:0] decipher_0_iibox_address21;
reg    decipher_0_iibox_ce21;
wire   [7:0] decipher_0_iibox_q21;
wire   [7:0] decipher_0_iibox_address22;
reg    decipher_0_iibox_ce22;
wire   [7:0] decipher_0_iibox_q22;
wire   [7:0] decipher_0_iibox_address23;
reg    decipher_0_iibox_ce23;
wire   [7:0] decipher_0_iibox_q23;
wire   [7:0] decipher_0_iibox_address24;
reg    decipher_0_iibox_ce24;
wire   [7:0] decipher_0_iibox_q24;
wire   [7:0] decipher_0_iibox_address25;
reg    decipher_0_iibox_ce25;
wire   [7:0] decipher_0_iibox_q25;
wire   [7:0] decipher_0_iibox_address26;
reg    decipher_0_iibox_ce26;
wire   [7:0] decipher_0_iibox_q26;
wire   [7:0] decipher_0_iibox_address27;
reg    decipher_0_iibox_ce27;
wire   [7:0] decipher_0_iibox_q27;
wire   [7:0] decipher_0_iibox_address28;
reg    decipher_0_iibox_ce28;
wire   [7:0] decipher_0_iibox_q28;
wire   [7:0] decipher_0_iibox_address29;
reg    decipher_0_iibox_ce29;
wire   [7:0] decipher_0_iibox_q29;
wire   [7:0] decipher_0_iibox_address30;
reg    decipher_0_iibox_ce30;
wire   [7:0] decipher_0_iibox_q30;
wire   [7:0] decipher_0_iibox_address31;
reg    decipher_0_iibox_ce31;
wire   [7:0] decipher_0_iibox_q31;
wire   [7:0] decipher_0_iibox_address32;
reg    decipher_0_iibox_ce32;
wire   [7:0] decipher_0_iibox_q32;
wire   [7:0] decipher_0_iibox_address33;
reg    decipher_0_iibox_ce33;
wire   [7:0] decipher_0_iibox_q33;
wire   [7:0] decipher_0_iibox_address34;
reg    decipher_0_iibox_ce34;
wire   [7:0] decipher_0_iibox_q34;
wire   [7:0] decipher_0_iibox_address35;
reg    decipher_0_iibox_ce35;
wire   [7:0] decipher_0_iibox_q35;
wire   [7:0] decipher_0_iibox_address36;
reg    decipher_0_iibox_ce36;
wire   [7:0] decipher_0_iibox_q36;
wire   [7:0] decipher_0_iibox_address37;
reg    decipher_0_iibox_ce37;
wire   [7:0] decipher_0_iibox_q37;
wire   [7:0] decipher_0_iibox_address38;
reg    decipher_0_iibox_ce38;
wire   [7:0] decipher_0_iibox_q38;
wire   [7:0] decipher_0_iibox_address39;
reg    decipher_0_iibox_ce39;
wire   [7:0] decipher_0_iibox_q39;
wire   [7:0] decipher_0_iibox_address40;
reg    decipher_0_iibox_ce40;
wire   [7:0] decipher_0_iibox_q40;
wire   [7:0] decipher_0_iibox_address41;
reg    decipher_0_iibox_ce41;
wire   [7:0] decipher_0_iibox_q41;
wire   [7:0] decipher_0_iibox_address42;
reg    decipher_0_iibox_ce42;
wire   [7:0] decipher_0_iibox_q42;
wire   [7:0] decipher_0_iibox_address43;
reg    decipher_0_iibox_ce43;
wire   [7:0] decipher_0_iibox_q43;
wire   [7:0] decipher_0_iibox_address44;
reg    decipher_0_iibox_ce44;
wire   [7:0] decipher_0_iibox_q44;
wire   [7:0] decipher_0_iibox_address45;
reg    decipher_0_iibox_ce45;
wire   [7:0] decipher_0_iibox_q45;
wire   [7:0] decipher_0_iibox_address46;
reg    decipher_0_iibox_ce46;
wire   [7:0] decipher_0_iibox_q46;
wire   [7:0] decipher_0_iibox_address47;
reg    decipher_0_iibox_ce47;
wire   [7:0] decipher_0_iibox_q47;
wire   [7:0] decipher_0_iibox_address48;
reg    decipher_0_iibox_ce48;
wire   [7:0] decipher_0_iibox_q48;
wire   [7:0] decipher_0_iibox_address49;
reg    decipher_0_iibox_ce49;
wire   [7:0] decipher_0_iibox_q49;
wire   [7:0] decipher_0_iibox_address50;
reg    decipher_0_iibox_ce50;
wire   [7:0] decipher_0_iibox_q50;
wire   [7:0] decipher_0_iibox_address51;
reg    decipher_0_iibox_ce51;
wire   [7:0] decipher_0_iibox_q51;
wire   [7:0] decipher_0_iibox_address52;
reg    decipher_0_iibox_ce52;
wire   [7:0] decipher_0_iibox_q52;
wire   [7:0] decipher_0_iibox_address53;
reg    decipher_0_iibox_ce53;
wire   [7:0] decipher_0_iibox_q53;
wire   [7:0] decipher_0_iibox_address54;
reg    decipher_0_iibox_ce54;
wire   [7:0] decipher_0_iibox_q54;
wire   [7:0] decipher_0_iibox_address55;
reg    decipher_0_iibox_ce55;
wire   [7:0] decipher_0_iibox_q55;
wire   [7:0] decipher_0_iibox_address56;
reg    decipher_0_iibox_ce56;
wire   [7:0] decipher_0_iibox_q56;
wire   [7:0] decipher_0_iibox_address57;
reg    decipher_0_iibox_ce57;
wire   [7:0] decipher_0_iibox_q57;
wire   [7:0] decipher_0_iibox_address58;
reg    decipher_0_iibox_ce58;
wire   [7:0] decipher_0_iibox_q58;
wire   [7:0] decipher_0_iibox_address59;
reg    decipher_0_iibox_ce59;
wire   [7:0] decipher_0_iibox_q59;
wire   [7:0] decipher_0_iibox_address60;
reg    decipher_0_iibox_ce60;
wire   [7:0] decipher_0_iibox_q60;
wire   [7:0] decipher_0_iibox_address61;
reg    decipher_0_iibox_ce61;
wire   [7:0] decipher_0_iibox_q61;
wire   [7:0] decipher_0_iibox_address62;
reg    decipher_0_iibox_ce62;
wire   [7:0] decipher_0_iibox_q62;
wire   [7:0] decipher_0_iibox_address63;
reg    decipher_0_iibox_ce63;
wire   [7:0] decipher_0_iibox_q63;
wire   [7:0] decipher_0_iibox_address64;
reg    decipher_0_iibox_ce64;
wire   [7:0] decipher_0_iibox_q64;
wire   [7:0] decipher_0_iibox_address65;
reg    decipher_0_iibox_ce65;
wire   [7:0] decipher_0_iibox_q65;
wire   [7:0] decipher_0_iibox_address66;
reg    decipher_0_iibox_ce66;
wire   [7:0] decipher_0_iibox_q66;
wire   [7:0] decipher_0_iibox_address67;
reg    decipher_0_iibox_ce67;
wire   [7:0] decipher_0_iibox_q67;
wire   [7:0] decipher_0_iibox_address68;
reg    decipher_0_iibox_ce68;
wire   [7:0] decipher_0_iibox_q68;
wire   [7:0] decipher_0_iibox_address69;
reg    decipher_0_iibox_ce69;
wire   [7:0] decipher_0_iibox_q69;
wire   [7:0] decipher_0_iibox_address70;
reg    decipher_0_iibox_ce70;
wire   [7:0] decipher_0_iibox_q70;
wire   [7:0] decipher_0_iibox_address71;
reg    decipher_0_iibox_ce71;
wire   [7:0] decipher_0_iibox_q71;
wire   [7:0] decipher_0_iibox_address72;
reg    decipher_0_iibox_ce72;
wire   [7:0] decipher_0_iibox_q72;
wire   [7:0] decipher_0_iibox_address73;
reg    decipher_0_iibox_ce73;
wire   [7:0] decipher_0_iibox_q73;
wire   [7:0] decipher_0_iibox_address74;
reg    decipher_0_iibox_ce74;
wire   [7:0] decipher_0_iibox_q74;
wire   [7:0] decipher_0_iibox_address75;
reg    decipher_0_iibox_ce75;
wire   [7:0] decipher_0_iibox_q75;
wire   [7:0] decipher_0_iibox_address76;
reg    decipher_0_iibox_ce76;
wire   [7:0] decipher_0_iibox_q76;
wire   [7:0] decipher_0_iibox_address77;
reg    decipher_0_iibox_ce77;
wire   [7:0] decipher_0_iibox_q77;
wire   [7:0] decipher_0_iibox_address78;
reg    decipher_0_iibox_ce78;
wire   [7:0] decipher_0_iibox_q78;
wire   [7:0] decipher_0_iibox_address79;
reg    decipher_0_iibox_ce79;
wire   [7:0] decipher_0_iibox_q79;
wire   [7:0] decipher_0_iibox_address80;
reg    decipher_0_iibox_ce80;
wire   [7:0] decipher_0_iibox_q80;
wire   [7:0] decipher_0_iibox_address81;
reg    decipher_0_iibox_ce81;
wire   [7:0] decipher_0_iibox_q81;
wire   [7:0] decipher_0_iibox_address82;
reg    decipher_0_iibox_ce82;
wire   [7:0] decipher_0_iibox_q82;
wire   [7:0] decipher_0_iibox_address83;
reg    decipher_0_iibox_ce83;
wire   [7:0] decipher_0_iibox_q83;
wire   [7:0] decipher_0_iibox_address84;
reg    decipher_0_iibox_ce84;
wire   [7:0] decipher_0_iibox_q84;
wire   [7:0] decipher_0_iibox_address85;
reg    decipher_0_iibox_ce85;
wire   [7:0] decipher_0_iibox_q85;
wire   [7:0] decipher_0_iibox_address86;
reg    decipher_0_iibox_ce86;
wire   [7:0] decipher_0_iibox_q86;
wire   [7:0] decipher_0_iibox_address87;
reg    decipher_0_iibox_ce87;
wire   [7:0] decipher_0_iibox_q87;
wire   [7:0] decipher_0_iibox_address88;
reg    decipher_0_iibox_ce88;
wire   [7:0] decipher_0_iibox_q88;
wire   [7:0] decipher_0_iibox_address89;
reg    decipher_0_iibox_ce89;
wire   [7:0] decipher_0_iibox_q89;
wire   [7:0] decipher_0_iibox_address90;
reg    decipher_0_iibox_ce90;
wire   [7:0] decipher_0_iibox_q90;
wire   [7:0] decipher_0_iibox_address91;
reg    decipher_0_iibox_ce91;
wire   [7:0] decipher_0_iibox_q91;
wire   [7:0] decipher_0_iibox_address92;
reg    decipher_0_iibox_ce92;
wire   [7:0] decipher_0_iibox_q92;
wire   [7:0] decipher_0_iibox_address93;
reg    decipher_0_iibox_ce93;
wire   [7:0] decipher_0_iibox_q93;
wire   [7:0] decipher_0_iibox_address94;
reg    decipher_0_iibox_ce94;
wire   [7:0] decipher_0_iibox_q94;
wire   [7:0] decipher_0_iibox_address95;
reg    decipher_0_iibox_ce95;
wire   [7:0] decipher_0_iibox_q95;
wire   [7:0] decipher_0_iibox_address96;
reg    decipher_0_iibox_ce96;
wire   [7:0] decipher_0_iibox_q96;
wire   [7:0] decipher_0_iibox_address97;
reg    decipher_0_iibox_ce97;
wire   [7:0] decipher_0_iibox_q97;
wire   [7:0] decipher_0_iibox_address98;
reg    decipher_0_iibox_ce98;
wire   [7:0] decipher_0_iibox_q98;
wire   [7:0] decipher_0_iibox_address99;
reg    decipher_0_iibox_ce99;
wire   [7:0] decipher_0_iibox_q99;
wire   [7:0] decipher_0_iibox_address100;
reg    decipher_0_iibox_ce100;
wire   [7:0] decipher_0_iibox_q100;
wire   [7:0] decipher_0_iibox_address101;
reg    decipher_0_iibox_ce101;
wire   [7:0] decipher_0_iibox_q101;
wire   [7:0] decipher_0_iibox_address102;
reg    decipher_0_iibox_ce102;
wire   [7:0] decipher_0_iibox_q102;
wire   [7:0] decipher_0_iibox_address103;
reg    decipher_0_iibox_ce103;
wire   [7:0] decipher_0_iibox_q103;
wire   [7:0] decipher_0_iibox_address104;
reg    decipher_0_iibox_ce104;
wire   [7:0] decipher_0_iibox_q104;
wire   [7:0] decipher_0_iibox_address105;
reg    decipher_0_iibox_ce105;
wire   [7:0] decipher_0_iibox_q105;
wire   [7:0] decipher_0_iibox_address106;
reg    decipher_0_iibox_ce106;
wire   [7:0] decipher_0_iibox_q106;
wire   [7:0] decipher_0_iibox_address107;
reg    decipher_0_iibox_ce107;
wire   [7:0] decipher_0_iibox_q107;
wire   [7:0] decipher_0_iibox_address108;
reg    decipher_0_iibox_ce108;
wire   [7:0] decipher_0_iibox_q108;
wire   [7:0] decipher_0_iibox_address109;
reg    decipher_0_iibox_ce109;
wire   [7:0] decipher_0_iibox_q109;
wire   [7:0] decipher_0_iibox_address110;
reg    decipher_0_iibox_ce110;
wire   [7:0] decipher_0_iibox_q110;
wire   [7:0] decipher_0_iibox_address111;
reg    decipher_0_iibox_ce111;
wire   [7:0] decipher_0_iibox_q111;
wire   [7:0] decipher_0_iibox_address112;
reg    decipher_0_iibox_ce112;
wire   [7:0] decipher_0_iibox_q112;
wire   [7:0] decipher_0_iibox_address113;
reg    decipher_0_iibox_ce113;
wire   [7:0] decipher_0_iibox_q113;
wire   [7:0] decipher_0_iibox_address114;
reg    decipher_0_iibox_ce114;
wire   [7:0] decipher_0_iibox_q114;
wire   [7:0] decipher_0_iibox_address115;
reg    decipher_0_iibox_ce115;
wire   [7:0] decipher_0_iibox_q115;
wire   [7:0] decipher_0_iibox_address116;
reg    decipher_0_iibox_ce116;
wire   [7:0] decipher_0_iibox_q116;
wire   [7:0] decipher_0_iibox_address117;
reg    decipher_0_iibox_ce117;
wire   [7:0] decipher_0_iibox_q117;
wire   [7:0] decipher_0_iibox_address118;
reg    decipher_0_iibox_ce118;
wire   [7:0] decipher_0_iibox_q118;
wire   [7:0] decipher_0_iibox_address119;
reg    decipher_0_iibox_ce119;
wire   [7:0] decipher_0_iibox_q119;
wire   [7:0] decipher_0_iibox_address120;
reg    decipher_0_iibox_ce120;
wire   [7:0] decipher_0_iibox_q120;
wire   [7:0] decipher_0_iibox_address121;
reg    decipher_0_iibox_ce121;
wire   [7:0] decipher_0_iibox_q121;
wire   [7:0] decipher_0_iibox_address122;
reg    decipher_0_iibox_ce122;
wire   [7:0] decipher_0_iibox_q122;
wire   [7:0] decipher_0_iibox_address123;
reg    decipher_0_iibox_ce123;
wire   [7:0] decipher_0_iibox_q123;
wire   [7:0] decipher_0_iibox_address124;
reg    decipher_0_iibox_ce124;
wire   [7:0] decipher_0_iibox_q124;
wire   [7:0] decipher_0_iibox_address125;
reg    decipher_0_iibox_ce125;
wire   [7:0] decipher_0_iibox_q125;
wire   [7:0] decipher_0_iibox_address126;
reg    decipher_0_iibox_ce126;
wire   [7:0] decipher_0_iibox_q126;
wire   [7:0] decipher_0_iibox_address127;
reg    decipher_0_iibox_ce127;
wire   [7:0] decipher_0_iibox_q127;
wire   [7:0] decipher_0_iibox_address128;
reg    decipher_0_iibox_ce128;
wire   [7:0] decipher_0_iibox_q128;
wire   [7:0] decipher_0_iibox_address129;
reg    decipher_0_iibox_ce129;
wire   [7:0] decipher_0_iibox_q129;
wire   [7:0] decipher_0_iibox_address130;
reg    decipher_0_iibox_ce130;
wire   [7:0] decipher_0_iibox_q130;
wire   [7:0] decipher_0_iibox_address131;
reg    decipher_0_iibox_ce131;
wire   [7:0] decipher_0_iibox_q131;
wire   [7:0] decipher_0_iibox_address132;
reg    decipher_0_iibox_ce132;
wire   [7:0] decipher_0_iibox_q132;
wire   [7:0] decipher_0_iibox_address133;
reg    decipher_0_iibox_ce133;
wire   [7:0] decipher_0_iibox_q133;
wire   [7:0] decipher_0_iibox_address134;
reg    decipher_0_iibox_ce134;
wire   [7:0] decipher_0_iibox_q134;
wire   [7:0] decipher_0_iibox_address135;
reg    decipher_0_iibox_ce135;
wire   [7:0] decipher_0_iibox_q135;
wire   [7:0] decipher_0_iibox_address136;
reg    decipher_0_iibox_ce136;
wire   [7:0] decipher_0_iibox_q136;
wire   [7:0] decipher_0_iibox_address137;
reg    decipher_0_iibox_ce137;
wire   [7:0] decipher_0_iibox_q137;
wire   [7:0] decipher_0_iibox_address138;
reg    decipher_0_iibox_ce138;
wire   [7:0] decipher_0_iibox_q138;
wire   [7:0] decipher_0_iibox_address139;
reg    decipher_0_iibox_ce139;
wire   [7:0] decipher_0_iibox_q139;
wire   [7:0] decipher_0_iibox_address140;
reg    decipher_0_iibox_ce140;
wire   [7:0] decipher_0_iibox_q140;
wire   [7:0] decipher_0_iibox_address141;
reg    decipher_0_iibox_ce141;
wire   [7:0] decipher_0_iibox_q141;
wire   [7:0] decipher_0_iibox_address142;
reg    decipher_0_iibox_ce142;
wire   [7:0] decipher_0_iibox_q142;
wire   [7:0] decipher_0_iibox_address143;
reg    decipher_0_iibox_ce143;
wire   [7:0] decipher_0_iibox_q143;
wire   [7:0] decipher_0_iibox_address144;
reg    decipher_0_iibox_ce144;
wire   [7:0] decipher_0_iibox_q144;
wire   [7:0] decipher_0_iibox_address145;
reg    decipher_0_iibox_ce145;
wire   [7:0] decipher_0_iibox_q145;
wire   [7:0] decipher_0_iibox_address146;
reg    decipher_0_iibox_ce146;
wire   [7:0] decipher_0_iibox_q146;
wire   [7:0] decipher_0_iibox_address147;
reg    decipher_0_iibox_ce147;
wire   [7:0] decipher_0_iibox_q147;
wire   [7:0] decipher_0_iibox_address148;
reg    decipher_0_iibox_ce148;
wire   [7:0] decipher_0_iibox_q148;
wire   [7:0] decipher_0_iibox_address149;
reg    decipher_0_iibox_ce149;
wire   [7:0] decipher_0_iibox_q149;
wire   [7:0] decipher_0_iibox_address150;
reg    decipher_0_iibox_ce150;
wire   [7:0] decipher_0_iibox_q150;
wire   [7:0] decipher_0_iibox_address151;
reg    decipher_0_iibox_ce151;
wire   [7:0] decipher_0_iibox_q151;
wire   [7:0] decipher_0_iibox_address152;
reg    decipher_0_iibox_ce152;
wire   [7:0] decipher_0_iibox_q152;
wire   [7:0] decipher_0_iibox_address153;
reg    decipher_0_iibox_ce153;
wire   [7:0] decipher_0_iibox_q153;
wire   [7:0] decipher_0_iibox_address154;
reg    decipher_0_iibox_ce154;
wire   [7:0] decipher_0_iibox_q154;
wire   [7:0] decipher_0_iibox_address155;
reg    decipher_0_iibox_ce155;
wire   [7:0] decipher_0_iibox_q155;
wire   [7:0] decipher_0_iibox_address156;
reg    decipher_0_iibox_ce156;
wire   [7:0] decipher_0_iibox_q156;
wire   [7:0] decipher_0_iibox_address157;
reg    decipher_0_iibox_ce157;
wire   [7:0] decipher_0_iibox_q157;
wire   [7:0] decipher_0_iibox_address158;
reg    decipher_0_iibox_ce158;
wire   [7:0] decipher_0_iibox_q158;
wire   [7:0] decipher_0_iibox_address159;
reg    decipher_0_iibox_ce159;
wire   [7:0] decipher_0_iibox_q159;
wire   [7:0] decipher_0_i32box_address0;
reg    decipher_0_i32box_ce0;
wire   [31:0] decipher_0_i32box_q0;
wire   [7:0] decipher_0_i32box_address1;
reg    decipher_0_i32box_ce1;
wire   [31:0] decipher_0_i32box_q1;
wire   [7:0] decipher_0_i32box_address2;
reg    decipher_0_i32box_ce2;
wire   [31:0] decipher_0_i32box_q2;
wire   [7:0] decipher_0_i32box_address3;
reg    decipher_0_i32box_ce3;
wire   [31:0] decipher_0_i32box_q3;
wire   [7:0] decipher_0_i32box_address4;
reg    decipher_0_i32box_ce4;
wire   [31:0] decipher_0_i32box_q4;
wire   [7:0] decipher_0_i32box_address5;
reg    decipher_0_i32box_ce5;
wire   [31:0] decipher_0_i32box_q5;
wire   [7:0] decipher_0_i32box_address6;
reg    decipher_0_i32box_ce6;
wire   [31:0] decipher_0_i32box_q6;
wire   [7:0] decipher_0_i32box_address7;
reg    decipher_0_i32box_ce7;
wire   [31:0] decipher_0_i32box_q7;
wire   [7:0] decipher_0_i32box_address8;
reg    decipher_0_i32box_ce8;
wire   [31:0] decipher_0_i32box_q8;
wire   [7:0] decipher_0_i32box_address9;
reg    decipher_0_i32box_ce9;
wire   [31:0] decipher_0_i32box_q9;
wire   [7:0] decipher_0_i32box_address10;
reg    decipher_0_i32box_ce10;
wire   [31:0] decipher_0_i32box_q10;
wire   [7:0] decipher_0_i32box_address11;
reg    decipher_0_i32box_ce11;
wire   [31:0] decipher_0_i32box_q11;
wire   [7:0] decipher_0_i32box_address12;
reg    decipher_0_i32box_ce12;
wire   [31:0] decipher_0_i32box_q12;
wire   [7:0] decipher_0_i32box_address13;
reg    decipher_0_i32box_ce13;
wire   [31:0] decipher_0_i32box_q13;
wire   [7:0] decipher_0_i32box_address14;
reg    decipher_0_i32box_ce14;
wire   [31:0] decipher_0_i32box_q14;
wire   [7:0] decipher_0_i32box_address15;
reg    decipher_0_i32box_ce15;
wire   [31:0] decipher_0_i32box_q15;
wire   [7:0] decipher_0_i32box_address16;
reg    decipher_0_i32box_ce16;
wire   [31:0] decipher_0_i32box_q16;
wire   [7:0] decipher_0_i32box_address17;
reg    decipher_0_i32box_ce17;
wire   [31:0] decipher_0_i32box_q17;
wire   [7:0] decipher_0_i32box_address18;
reg    decipher_0_i32box_ce18;
wire   [31:0] decipher_0_i32box_q18;
wire   [7:0] decipher_0_i32box_address19;
reg    decipher_0_i32box_ce19;
wire   [31:0] decipher_0_i32box_q19;
wire   [7:0] decipher_0_i32box_address20;
reg    decipher_0_i32box_ce20;
wire   [31:0] decipher_0_i32box_q20;
wire   [7:0] decipher_0_i32box_address21;
reg    decipher_0_i32box_ce21;
wire   [31:0] decipher_0_i32box_q21;
wire   [7:0] decipher_0_i32box_address22;
reg    decipher_0_i32box_ce22;
wire   [31:0] decipher_0_i32box_q22;
wire   [7:0] decipher_0_i32box_address23;
reg    decipher_0_i32box_ce23;
wire   [31:0] decipher_0_i32box_q23;
wire   [7:0] decipher_0_i32box_address24;
reg    decipher_0_i32box_ce24;
wire   [31:0] decipher_0_i32box_q24;
wire   [7:0] decipher_0_i32box_address25;
reg    decipher_0_i32box_ce25;
wire   [31:0] decipher_0_i32box_q25;
wire   [7:0] decipher_0_i32box_address26;
reg    decipher_0_i32box_ce26;
wire   [31:0] decipher_0_i32box_q26;
wire   [7:0] decipher_0_i32box_address27;
reg    decipher_0_i32box_ce27;
wire   [31:0] decipher_0_i32box_q27;
wire   [7:0] decipher_0_i32box_address28;
reg    decipher_0_i32box_ce28;
wire   [31:0] decipher_0_i32box_q28;
wire   [7:0] decipher_0_i32box_address29;
reg    decipher_0_i32box_ce29;
wire   [31:0] decipher_0_i32box_q29;
wire   [7:0] decipher_0_i32box_address30;
reg    decipher_0_i32box_ce30;
wire   [31:0] decipher_0_i32box_q30;
wire   [7:0] decipher_0_i32box_address31;
reg    decipher_0_i32box_ce31;
wire   [31:0] decipher_0_i32box_q31;
wire   [7:0] decipher_0_i32box_address32;
reg    decipher_0_i32box_ce32;
wire   [31:0] decipher_0_i32box_q32;
wire   [7:0] decipher_0_i32box_address33;
reg    decipher_0_i32box_ce33;
wire   [31:0] decipher_0_i32box_q33;
wire   [7:0] decipher_0_i32box_address34;
reg    decipher_0_i32box_ce34;
wire   [31:0] decipher_0_i32box_q34;
wire   [7:0] decipher_0_i32box_address35;
reg    decipher_0_i32box_ce35;
wire   [31:0] decipher_0_i32box_q35;
wire   [7:0] decipher_0_i32box_address36;
reg    decipher_0_i32box_ce36;
wire   [31:0] decipher_0_i32box_q36;
wire   [7:0] decipher_0_i32box_address37;
reg    decipher_0_i32box_ce37;
wire   [31:0] decipher_0_i32box_q37;
wire   [7:0] decipher_0_i32box_address38;
reg    decipher_0_i32box_ce38;
wire   [31:0] decipher_0_i32box_q38;
wire   [7:0] decipher_0_i32box_address39;
reg    decipher_0_i32box_ce39;
wire   [31:0] decipher_0_i32box_q39;
wire   [7:0] decipher_0_i32box_address40;
reg    decipher_0_i32box_ce40;
wire   [31:0] decipher_0_i32box_q40;
wire   [7:0] decipher_0_i32box_address41;
reg    decipher_0_i32box_ce41;
wire   [31:0] decipher_0_i32box_q41;
wire   [7:0] decipher_0_i32box_address42;
reg    decipher_0_i32box_ce42;
wire   [31:0] decipher_0_i32box_q42;
wire   [7:0] decipher_0_i32box_address43;
reg    decipher_0_i32box_ce43;
wire   [31:0] decipher_0_i32box_q43;
wire   [7:0] decipher_0_i32box_address44;
reg    decipher_0_i32box_ce44;
wire   [31:0] decipher_0_i32box_q44;
wire   [7:0] decipher_0_i32box_address45;
reg    decipher_0_i32box_ce45;
wire   [31:0] decipher_0_i32box_q45;
wire   [7:0] decipher_0_i32box_address46;
reg    decipher_0_i32box_ce46;
wire   [31:0] decipher_0_i32box_q46;
wire   [7:0] decipher_0_i32box_address47;
reg    decipher_0_i32box_ce47;
wire   [31:0] decipher_0_i32box_q47;
wire   [7:0] decipher_0_i32box_address48;
reg    decipher_0_i32box_ce48;
wire   [31:0] decipher_0_i32box_q48;
wire   [7:0] decipher_0_i32box_address49;
reg    decipher_0_i32box_ce49;
wire   [31:0] decipher_0_i32box_q49;
wire   [7:0] decipher_0_i32box_address50;
reg    decipher_0_i32box_ce50;
wire   [31:0] decipher_0_i32box_q50;
wire   [7:0] decipher_0_i32box_address51;
reg    decipher_0_i32box_ce51;
wire   [31:0] decipher_0_i32box_q51;
wire   [7:0] decipher_0_i32box_address52;
reg    decipher_0_i32box_ce52;
wire   [31:0] decipher_0_i32box_q52;
wire   [7:0] decipher_0_i32box_address53;
reg    decipher_0_i32box_ce53;
wire   [31:0] decipher_0_i32box_q53;
wire   [7:0] decipher_0_i32box_address54;
reg    decipher_0_i32box_ce54;
wire   [31:0] decipher_0_i32box_q54;
wire   [7:0] decipher_0_i32box_address55;
reg    decipher_0_i32box_ce55;
wire   [31:0] decipher_0_i32box_q55;
wire   [7:0] decipher_0_i32box_address56;
reg    decipher_0_i32box_ce56;
wire   [31:0] decipher_0_i32box_q56;
wire   [7:0] decipher_0_i32box_address57;
reg    decipher_0_i32box_ce57;
wire   [31:0] decipher_0_i32box_q57;
wire   [7:0] decipher_0_i32box_address58;
reg    decipher_0_i32box_ce58;
wire   [31:0] decipher_0_i32box_q58;
wire   [7:0] decipher_0_i32box_address59;
reg    decipher_0_i32box_ce59;
wire   [31:0] decipher_0_i32box_q59;
wire   [7:0] decipher_0_i32box_address60;
reg    decipher_0_i32box_ce60;
wire   [31:0] decipher_0_i32box_q60;
wire   [7:0] decipher_0_i32box_address61;
reg    decipher_0_i32box_ce61;
wire   [31:0] decipher_0_i32box_q61;
wire   [7:0] decipher_0_i32box_address62;
reg    decipher_0_i32box_ce62;
wire   [31:0] decipher_0_i32box_q62;
wire   [7:0] decipher_0_i32box_address63;
reg    decipher_0_i32box_ce63;
wire   [31:0] decipher_0_i32box_q63;
wire   [7:0] decipher_0_i32box_address64;
reg    decipher_0_i32box_ce64;
wire   [31:0] decipher_0_i32box_q64;
wire   [7:0] decipher_0_i32box_address65;
reg    decipher_0_i32box_ce65;
wire   [31:0] decipher_0_i32box_q65;
wire   [7:0] decipher_0_i32box_address66;
reg    decipher_0_i32box_ce66;
wire   [31:0] decipher_0_i32box_q66;
wire   [7:0] decipher_0_i32box_address67;
reg    decipher_0_i32box_ce67;
wire   [31:0] decipher_0_i32box_q67;
wire   [7:0] decipher_0_i32box_address68;
reg    decipher_0_i32box_ce68;
wire   [31:0] decipher_0_i32box_q68;
wire   [7:0] decipher_0_i32box_address69;
reg    decipher_0_i32box_ce69;
wire   [31:0] decipher_0_i32box_q69;
wire   [7:0] decipher_0_i32box_address70;
reg    decipher_0_i32box_ce70;
wire   [31:0] decipher_0_i32box_q70;
wire   [7:0] decipher_0_i32box_address71;
reg    decipher_0_i32box_ce71;
wire   [31:0] decipher_0_i32box_q71;
wire   [7:0] decipher_0_i32box_address72;
reg    decipher_0_i32box_ce72;
wire   [31:0] decipher_0_i32box_q72;
wire   [7:0] decipher_0_i32box_address73;
reg    decipher_0_i32box_ce73;
wire   [31:0] decipher_0_i32box_q73;
wire   [7:0] decipher_0_i32box_address74;
reg    decipher_0_i32box_ce74;
wire   [31:0] decipher_0_i32box_q74;
wire   [7:0] decipher_0_i32box_address75;
reg    decipher_0_i32box_ce75;
wire   [31:0] decipher_0_i32box_q75;
wire   [7:0] decipher_0_i32box_address76;
reg    decipher_0_i32box_ce76;
wire   [31:0] decipher_0_i32box_q76;
wire   [7:0] decipher_0_i32box_address77;
reg    decipher_0_i32box_ce77;
wire   [31:0] decipher_0_i32box_q77;
wire   [7:0] decipher_0_i32box_address78;
reg    decipher_0_i32box_ce78;
wire   [31:0] decipher_0_i32box_q78;
wire   [7:0] decipher_0_i32box_address79;
reg    decipher_0_i32box_ce79;
wire   [31:0] decipher_0_i32box_q79;
wire   [7:0] decipher_0_i32box_address80;
reg    decipher_0_i32box_ce80;
wire   [31:0] decipher_0_i32box_q80;
wire   [7:0] decipher_0_i32box_address81;
reg    decipher_0_i32box_ce81;
wire   [31:0] decipher_0_i32box_q81;
wire   [7:0] decipher_0_i32box_address82;
reg    decipher_0_i32box_ce82;
wire   [31:0] decipher_0_i32box_q82;
wire   [7:0] decipher_0_i32box_address83;
reg    decipher_0_i32box_ce83;
wire   [31:0] decipher_0_i32box_q83;
wire   [7:0] decipher_0_i32box_address84;
reg    decipher_0_i32box_ce84;
wire   [31:0] decipher_0_i32box_q84;
wire   [7:0] decipher_0_i32box_address85;
reg    decipher_0_i32box_ce85;
wire   [31:0] decipher_0_i32box_q85;
wire   [7:0] decipher_0_i32box_address86;
reg    decipher_0_i32box_ce86;
wire   [31:0] decipher_0_i32box_q86;
wire   [7:0] decipher_0_i32box_address87;
reg    decipher_0_i32box_ce87;
wire   [31:0] decipher_0_i32box_q87;
wire   [7:0] decipher_0_i32box_address88;
reg    decipher_0_i32box_ce88;
wire   [31:0] decipher_0_i32box_q88;
wire   [7:0] decipher_0_i32box_address89;
reg    decipher_0_i32box_ce89;
wire   [31:0] decipher_0_i32box_q89;
wire   [7:0] decipher_0_i32box_address90;
reg    decipher_0_i32box_ce90;
wire   [31:0] decipher_0_i32box_q90;
wire   [7:0] decipher_0_i32box_address91;
reg    decipher_0_i32box_ce91;
wire   [31:0] decipher_0_i32box_q91;
wire   [7:0] decipher_0_i32box_address92;
reg    decipher_0_i32box_ce92;
wire   [31:0] decipher_0_i32box_q92;
wire   [7:0] decipher_0_i32box_address93;
reg    decipher_0_i32box_ce93;
wire   [31:0] decipher_0_i32box_q93;
wire   [7:0] decipher_0_i32box_address94;
reg    decipher_0_i32box_ce94;
wire   [31:0] decipher_0_i32box_q94;
wire   [7:0] decipher_0_i32box_address95;
reg    decipher_0_i32box_ce95;
wire   [31:0] decipher_0_i32box_q95;
wire   [7:0] decipher_0_i32box_address96;
reg    decipher_0_i32box_ce96;
wire   [31:0] decipher_0_i32box_q96;
wire   [7:0] decipher_0_i32box_address97;
reg    decipher_0_i32box_ce97;
wire   [31:0] decipher_0_i32box_q97;
wire   [7:0] decipher_0_i32box_address98;
reg    decipher_0_i32box_ce98;
wire   [31:0] decipher_0_i32box_q98;
wire   [7:0] decipher_0_i32box_address99;
reg    decipher_0_i32box_ce99;
wire   [31:0] decipher_0_i32box_q99;
wire   [7:0] decipher_0_i32box_address100;
reg    decipher_0_i32box_ce100;
wire   [31:0] decipher_0_i32box_q100;
wire   [7:0] decipher_0_i32box_address101;
reg    decipher_0_i32box_ce101;
wire   [31:0] decipher_0_i32box_q101;
wire   [7:0] decipher_0_i32box_address102;
reg    decipher_0_i32box_ce102;
wire   [31:0] decipher_0_i32box_q102;
wire   [7:0] decipher_0_i32box_address103;
reg    decipher_0_i32box_ce103;
wire   [31:0] decipher_0_i32box_q103;
wire   [7:0] decipher_0_i32box_address104;
reg    decipher_0_i32box_ce104;
wire   [31:0] decipher_0_i32box_q104;
wire   [7:0] decipher_0_i32box_address105;
reg    decipher_0_i32box_ce105;
wire   [31:0] decipher_0_i32box_q105;
wire   [7:0] decipher_0_i32box_address106;
reg    decipher_0_i32box_ce106;
wire   [31:0] decipher_0_i32box_q106;
wire   [7:0] decipher_0_i32box_address107;
reg    decipher_0_i32box_ce107;
wire   [31:0] decipher_0_i32box_q107;
wire   [7:0] decipher_0_i32box_address108;
reg    decipher_0_i32box_ce108;
wire   [31:0] decipher_0_i32box_q108;
wire   [7:0] decipher_0_i32box_address109;
reg    decipher_0_i32box_ce109;
wire   [31:0] decipher_0_i32box_q109;
wire   [7:0] decipher_0_i32box_address110;
reg    decipher_0_i32box_ce110;
wire   [31:0] decipher_0_i32box_q110;
wire   [7:0] decipher_0_i32box_address111;
reg    decipher_0_i32box_ce111;
wire   [31:0] decipher_0_i32box_q111;
wire   [7:0] decipher_0_i32box_address112;
reg    decipher_0_i32box_ce112;
wire   [31:0] decipher_0_i32box_q112;
wire   [7:0] decipher_0_i32box_address113;
reg    decipher_0_i32box_ce113;
wire   [31:0] decipher_0_i32box_q113;
wire   [7:0] decipher_0_i32box_address114;
reg    decipher_0_i32box_ce114;
wire   [31:0] decipher_0_i32box_q114;
wire   [7:0] decipher_0_i32box_address115;
reg    decipher_0_i32box_ce115;
wire   [31:0] decipher_0_i32box_q115;
wire   [7:0] decipher_0_i32box_address116;
reg    decipher_0_i32box_ce116;
wire   [31:0] decipher_0_i32box_q116;
wire   [7:0] decipher_0_i32box_address117;
reg    decipher_0_i32box_ce117;
wire   [31:0] decipher_0_i32box_q117;
wire   [7:0] decipher_0_i32box_address118;
reg    decipher_0_i32box_ce118;
wire   [31:0] decipher_0_i32box_q118;
wire   [7:0] decipher_0_i32box_address119;
reg    decipher_0_i32box_ce119;
wire   [31:0] decipher_0_i32box_q119;
wire   [7:0] decipher_0_i32box_address120;
reg    decipher_0_i32box_ce120;
wire   [31:0] decipher_0_i32box_q120;
wire   [7:0] decipher_0_i32box_address121;
reg    decipher_0_i32box_ce121;
wire   [31:0] decipher_0_i32box_q121;
wire   [7:0] decipher_0_i32box_address122;
reg    decipher_0_i32box_ce122;
wire   [31:0] decipher_0_i32box_q122;
wire   [7:0] decipher_0_i32box_address123;
reg    decipher_0_i32box_ce123;
wire   [31:0] decipher_0_i32box_q123;
wire   [7:0] decipher_0_i32box_address124;
reg    decipher_0_i32box_ce124;
wire   [31:0] decipher_0_i32box_q124;
wire   [7:0] decipher_0_i32box_address125;
reg    decipher_0_i32box_ce125;
wire   [31:0] decipher_0_i32box_q125;
wire   [7:0] decipher_0_i32box_address126;
reg    decipher_0_i32box_ce126;
wire   [31:0] decipher_0_i32box_q126;
wire   [7:0] decipher_0_i32box_address127;
reg    decipher_0_i32box_ce127;
wire   [31:0] decipher_0_i32box_q127;
wire   [7:0] decipher_0_i32box_address128;
reg    decipher_0_i32box_ce128;
wire   [31:0] decipher_0_i32box_q128;
wire   [7:0] decipher_0_i32box_address129;
reg    decipher_0_i32box_ce129;
wire   [31:0] decipher_0_i32box_q129;
wire   [7:0] decipher_0_i32box_address130;
reg    decipher_0_i32box_ce130;
wire   [31:0] decipher_0_i32box_q130;
wire   [7:0] decipher_0_i32box_address131;
reg    decipher_0_i32box_ce131;
wire   [31:0] decipher_0_i32box_q131;
wire   [7:0] decipher_0_i32box_address132;
reg    decipher_0_i32box_ce132;
wire   [31:0] decipher_0_i32box_q132;
wire   [7:0] decipher_0_i32box_address133;
reg    decipher_0_i32box_ce133;
wire   [31:0] decipher_0_i32box_q133;
wire   [7:0] decipher_0_i32box_address134;
reg    decipher_0_i32box_ce134;
wire   [31:0] decipher_0_i32box_q134;
wire   [7:0] decipher_0_i32box_address135;
reg    decipher_0_i32box_ce135;
wire   [31:0] decipher_0_i32box_q135;
wire   [7:0] decipher_0_i32box_address136;
reg    decipher_0_i32box_ce136;
wire   [31:0] decipher_0_i32box_q136;
wire   [7:0] decipher_0_i32box_address137;
reg    decipher_0_i32box_ce137;
wire   [31:0] decipher_0_i32box_q137;
wire   [7:0] decipher_0_i32box_address138;
reg    decipher_0_i32box_ce138;
wire   [31:0] decipher_0_i32box_q138;
wire   [7:0] decipher_0_i32box_address139;
reg    decipher_0_i32box_ce139;
wire   [31:0] decipher_0_i32box_q139;
wire   [7:0] decipher_0_i32box_address140;
reg    decipher_0_i32box_ce140;
wire   [31:0] decipher_0_i32box_q140;
wire   [7:0] decipher_0_i32box_address141;
reg    decipher_0_i32box_ce141;
wire   [31:0] decipher_0_i32box_q141;
wire   [7:0] decipher_0_i32box_address142;
reg    decipher_0_i32box_ce142;
wire   [31:0] decipher_0_i32box_q142;
wire   [7:0] decipher_0_i32box_address143;
reg    decipher_0_i32box_ce143;
wire   [31:0] decipher_0_i32box_q143;
reg   [127:0] p_read_2_reg_14792;
wire    ap_block_pp0_stage0_11001;
reg   [127:0] p_read_3_reg_14797;
reg   [127:0] p_read_3_reg_14797_pp0_iter1_reg;
reg   [127:0] p_read_3_reg_14797_pp0_iter2_reg;
reg   [127:0] p_read_4_reg_14802;
reg   [127:0] p_read_4_reg_14802_pp0_iter1_reg;
reg   [127:0] p_read_4_reg_14802_pp0_iter2_reg;
reg   [127:0] p_read_4_reg_14802_pp0_iter3_reg;
reg   [127:0] p_read_4_reg_14802_pp0_iter4_reg;
reg   [127:0] p_read_5_reg_14807;
reg   [127:0] p_read_5_reg_14807_pp0_iter1_reg;
reg   [127:0] p_read_5_reg_14807_pp0_iter2_reg;
reg   [127:0] p_read_5_reg_14807_pp0_iter3_reg;
reg   [127:0] p_read_5_reg_14807_pp0_iter4_reg;
reg   [127:0] p_read_5_reg_14807_pp0_iter5_reg;
reg   [127:0] p_read_5_reg_14807_pp0_iter6_reg;
reg   [127:0] p_read_6_reg_14812;
reg   [127:0] p_read_6_reg_14812_pp0_iter1_reg;
reg   [127:0] p_read_6_reg_14812_pp0_iter2_reg;
reg   [127:0] p_read_6_reg_14812_pp0_iter3_reg;
reg   [127:0] p_read_6_reg_14812_pp0_iter4_reg;
reg   [127:0] p_read_6_reg_14812_pp0_iter5_reg;
reg   [127:0] p_read_6_reg_14812_pp0_iter6_reg;
reg   [127:0] p_read_6_reg_14812_pp0_iter7_reg;
reg   [127:0] p_read_6_reg_14812_pp0_iter8_reg;
reg   [127:0] p_read_7_reg_14817;
reg   [127:0] p_read_7_reg_14817_pp0_iter1_reg;
reg   [127:0] p_read_7_reg_14817_pp0_iter2_reg;
reg   [127:0] p_read_7_reg_14817_pp0_iter3_reg;
reg   [127:0] p_read_7_reg_14817_pp0_iter4_reg;
reg   [127:0] p_read_7_reg_14817_pp0_iter5_reg;
reg   [127:0] p_read_7_reg_14817_pp0_iter6_reg;
reg   [127:0] p_read_7_reg_14817_pp0_iter7_reg;
reg   [127:0] p_read_7_reg_14817_pp0_iter8_reg;
reg   [127:0] p_read_7_reg_14817_pp0_iter9_reg;
reg   [127:0] p_read_7_reg_14817_pp0_iter10_reg;
reg   [127:0] p_read_8_reg_14822;
reg   [127:0] p_read_8_reg_14822_pp0_iter1_reg;
reg   [127:0] p_read_8_reg_14822_pp0_iter2_reg;
reg   [127:0] p_read_8_reg_14822_pp0_iter3_reg;
reg   [127:0] p_read_8_reg_14822_pp0_iter4_reg;
reg   [127:0] p_read_8_reg_14822_pp0_iter5_reg;
reg   [127:0] p_read_8_reg_14822_pp0_iter6_reg;
reg   [127:0] p_read_8_reg_14822_pp0_iter7_reg;
reg   [127:0] p_read_8_reg_14822_pp0_iter8_reg;
reg   [127:0] p_read_8_reg_14822_pp0_iter9_reg;
reg   [127:0] p_read_8_reg_14822_pp0_iter10_reg;
reg   [127:0] p_read_8_reg_14822_pp0_iter11_reg;
reg   [127:0] p_read_8_reg_14822_pp0_iter12_reg;
reg   [127:0] p_read_9_reg_14827;
reg   [127:0] p_read_9_reg_14827_pp0_iter1_reg;
reg   [127:0] p_read_9_reg_14827_pp0_iter2_reg;
reg   [127:0] p_read_9_reg_14827_pp0_iter3_reg;
reg   [127:0] p_read_9_reg_14827_pp0_iter4_reg;
reg   [127:0] p_read_9_reg_14827_pp0_iter5_reg;
reg   [127:0] p_read_9_reg_14827_pp0_iter6_reg;
reg   [127:0] p_read_9_reg_14827_pp0_iter7_reg;
reg   [127:0] p_read_9_reg_14827_pp0_iter8_reg;
reg   [127:0] p_read_9_reg_14827_pp0_iter9_reg;
reg   [127:0] p_read_9_reg_14827_pp0_iter10_reg;
reg   [127:0] p_read_9_reg_14827_pp0_iter11_reg;
reg   [127:0] p_read_9_reg_14827_pp0_iter12_reg;
reg   [127:0] p_read_9_reg_14827_pp0_iter13_reg;
reg   [127:0] p_read_9_reg_14827_pp0_iter14_reg;
reg   [127:0] p_read_10_reg_14832;
reg   [127:0] p_read_10_reg_14832_pp0_iter1_reg;
reg   [127:0] p_read_10_reg_14832_pp0_iter2_reg;
reg   [127:0] p_read_10_reg_14832_pp0_iter3_reg;
reg   [127:0] p_read_10_reg_14832_pp0_iter4_reg;
reg   [127:0] p_read_10_reg_14832_pp0_iter5_reg;
reg   [127:0] p_read_10_reg_14832_pp0_iter6_reg;
reg   [127:0] p_read_10_reg_14832_pp0_iter7_reg;
reg   [127:0] p_read_10_reg_14832_pp0_iter8_reg;
reg   [127:0] p_read_10_reg_14832_pp0_iter9_reg;
reg   [127:0] p_read_10_reg_14832_pp0_iter10_reg;
reg   [127:0] p_read_10_reg_14832_pp0_iter11_reg;
reg   [127:0] p_read_10_reg_14832_pp0_iter12_reg;
reg   [127:0] p_read_10_reg_14832_pp0_iter13_reg;
reg   [127:0] p_read_10_reg_14832_pp0_iter14_reg;
reg   [127:0] p_read_10_reg_14832_pp0_iter15_reg;
reg   [127:0] p_read_10_reg_14832_pp0_iter16_reg;
reg   [127:0] p_read11_reg_14837;
reg   [127:0] p_read11_reg_14837_pp0_iter1_reg;
reg   [127:0] p_read11_reg_14837_pp0_iter2_reg;
reg   [127:0] p_read11_reg_14837_pp0_iter3_reg;
reg   [127:0] p_read11_reg_14837_pp0_iter4_reg;
reg   [127:0] p_read11_reg_14837_pp0_iter5_reg;
reg   [127:0] p_read11_reg_14837_pp0_iter6_reg;
reg   [127:0] p_read11_reg_14837_pp0_iter7_reg;
reg   [127:0] p_read11_reg_14837_pp0_iter8_reg;
reg   [127:0] p_read11_reg_14837_pp0_iter9_reg;
reg   [127:0] p_read11_reg_14837_pp0_iter10_reg;
reg   [127:0] p_read11_reg_14837_pp0_iter11_reg;
reg   [127:0] p_read11_reg_14837_pp0_iter12_reg;
reg   [127:0] p_read11_reg_14837_pp0_iter13_reg;
reg   [127:0] p_read11_reg_14837_pp0_iter14_reg;
reg   [127:0] p_read11_reg_14837_pp0_iter15_reg;
reg   [127:0] p_read11_reg_14837_pp0_iter16_reg;
reg   [127:0] p_read11_reg_14837_pp0_iter17_reg;
reg   [127:0] p_read11_reg_14837_pp0_iter18_reg;
wire   [63:0] zext_ln708_fu_3838_p1;
wire    ap_block_pp0_stage0;
wire   [63:0] zext_ln708_4_fu_3853_p1;
wire   [63:0] zext_ln708_5_fu_3868_p1;
wire   [63:0] zext_ln708_6_fu_3883_p1;
wire   [63:0] zext_ln708_7_fu_3898_p1;
wire   [63:0] zext_ln708_8_fu_3913_p1;
wire   [63:0] zext_ln708_9_fu_3928_p1;
wire   [63:0] zext_ln708_10_fu_3943_p1;
wire   [63:0] zext_ln708_11_fu_3958_p1;
wire   [63:0] zext_ln708_12_fu_3973_p1;
wire   [63:0] zext_ln708_13_fu_3988_p1;
wire   [63:0] zext_ln708_14_fu_4003_p1;
wire   [63:0] zext_ln708_15_fu_4018_p1;
wire   [63:0] zext_ln708_16_fu_4033_p1;
wire   [63:0] zext_ln708_17_fu_4048_p1;
wire   [63:0] zext_ln708_18_fu_4063_p1;
wire   [63:0] zext_ln708_19_fu_4113_p1;
wire   [63:0] zext_ln708_20_fu_4128_p1;
wire   [63:0] zext_ln708_21_fu_4143_p1;
wire   [63:0] zext_ln708_22_fu_4158_p1;
wire   [63:0] zext_ln708_23_fu_4173_p1;
wire   [63:0] zext_ln708_24_fu_4188_p1;
wire   [63:0] zext_ln708_25_fu_4203_p1;
wire   [63:0] zext_ln708_26_fu_4218_p1;
wire   [63:0] zext_ln708_27_fu_4233_p1;
wire   [63:0] zext_ln708_28_fu_4248_p1;
wire   [63:0] zext_ln708_29_fu_4263_p1;
wire   [63:0] zext_ln708_30_fu_4278_p1;
wire   [63:0] zext_ln708_31_fu_4293_p1;
wire   [63:0] zext_ln708_32_fu_4308_p1;
wire   [63:0] zext_ln708_33_fu_4323_p1;
wire   [63:0] zext_ln708_34_fu_4338_p1;
wire   [63:0] zext_ln708_35_fu_5175_p1;
wire   [63:0] zext_ln708_36_fu_5180_p1;
wire   [63:0] zext_ln708_37_fu_5185_p1;
wire   [63:0] zext_ln708_38_fu_5190_p1;
wire   [63:0] zext_ln708_39_fu_5195_p1;
wire   [63:0] zext_ln708_40_fu_5200_p1;
wire   [63:0] zext_ln708_41_fu_5205_p1;
wire   [63:0] zext_ln708_42_fu_5210_p1;
wire   [63:0] zext_ln708_43_fu_5215_p1;
wire   [63:0] zext_ln708_44_fu_5220_p1;
wire   [63:0] zext_ln708_45_fu_5225_p1;
wire   [63:0] zext_ln708_46_fu_5230_p1;
wire   [63:0] zext_ln708_47_fu_5235_p1;
wire   [63:0] zext_ln708_48_fu_5240_p1;
wire   [63:0] zext_ln708_49_fu_5245_p1;
wire   [63:0] zext_ln708_50_fu_5250_p1;
wire   [63:0] zext_ln708_51_fu_5300_p1;
wire   [63:0] zext_ln708_52_fu_5315_p1;
wire   [63:0] zext_ln708_53_fu_5330_p1;
wire   [63:0] zext_ln708_54_fu_5345_p1;
wire   [63:0] zext_ln708_55_fu_5360_p1;
wire   [63:0] zext_ln708_56_fu_5375_p1;
wire   [63:0] zext_ln708_57_fu_5390_p1;
wire   [63:0] zext_ln708_58_fu_5405_p1;
wire   [63:0] zext_ln708_59_fu_5420_p1;
wire   [63:0] zext_ln708_60_fu_5435_p1;
wire   [63:0] zext_ln708_61_fu_5450_p1;
wire   [63:0] zext_ln708_62_fu_5465_p1;
wire   [63:0] zext_ln708_63_fu_5480_p1;
wire   [63:0] zext_ln708_64_fu_5495_p1;
wire   [63:0] zext_ln708_65_fu_5510_p1;
wire   [63:0] zext_ln708_66_fu_5525_p1;
wire   [63:0] zext_ln708_67_fu_6362_p1;
wire   [63:0] zext_ln708_68_fu_6367_p1;
wire   [63:0] zext_ln708_69_fu_6372_p1;
wire   [63:0] zext_ln708_70_fu_6377_p1;
wire   [63:0] zext_ln708_71_fu_6382_p1;
wire   [63:0] zext_ln708_72_fu_6387_p1;
wire   [63:0] zext_ln708_73_fu_6392_p1;
wire   [63:0] zext_ln708_74_fu_6397_p1;
wire   [63:0] zext_ln708_75_fu_6402_p1;
wire   [63:0] zext_ln708_76_fu_6407_p1;
wire   [63:0] zext_ln708_77_fu_6412_p1;
wire   [63:0] zext_ln708_78_fu_6417_p1;
wire   [63:0] zext_ln708_79_fu_6422_p1;
wire   [63:0] zext_ln708_80_fu_6427_p1;
wire   [63:0] zext_ln708_81_fu_6432_p1;
wire   [63:0] zext_ln708_82_fu_6437_p1;
wire   [63:0] zext_ln708_83_fu_6487_p1;
wire   [63:0] zext_ln708_84_fu_6502_p1;
wire   [63:0] zext_ln708_85_fu_6517_p1;
wire   [63:0] zext_ln708_86_fu_6532_p1;
wire   [63:0] zext_ln708_87_fu_6547_p1;
wire   [63:0] zext_ln708_88_fu_6562_p1;
wire   [63:0] zext_ln708_89_fu_6577_p1;
wire   [63:0] zext_ln708_90_fu_6592_p1;
wire   [63:0] zext_ln708_91_fu_6607_p1;
wire   [63:0] zext_ln708_92_fu_6622_p1;
wire   [63:0] zext_ln708_93_fu_6637_p1;
wire   [63:0] zext_ln708_94_fu_6652_p1;
wire   [63:0] zext_ln708_95_fu_6667_p1;
wire   [63:0] zext_ln708_96_fu_6682_p1;
wire   [63:0] zext_ln708_97_fu_6697_p1;
wire   [63:0] zext_ln708_98_fu_6712_p1;
wire   [63:0] zext_ln708_99_fu_7549_p1;
wire   [63:0] zext_ln708_100_fu_7554_p1;
wire   [63:0] zext_ln708_101_fu_7559_p1;
wire   [63:0] zext_ln708_102_fu_7564_p1;
wire   [63:0] zext_ln708_103_fu_7569_p1;
wire   [63:0] zext_ln708_104_fu_7574_p1;
wire   [63:0] zext_ln708_105_fu_7579_p1;
wire   [63:0] zext_ln708_106_fu_7584_p1;
wire   [63:0] zext_ln708_107_fu_7589_p1;
wire   [63:0] zext_ln708_108_fu_7594_p1;
wire   [63:0] zext_ln708_109_fu_7599_p1;
wire   [63:0] zext_ln708_110_fu_7604_p1;
wire   [63:0] zext_ln708_111_fu_7609_p1;
wire   [63:0] zext_ln708_112_fu_7614_p1;
wire   [63:0] zext_ln708_113_fu_7619_p1;
wire   [63:0] zext_ln708_114_fu_7624_p1;
wire   [63:0] zext_ln708_115_fu_7674_p1;
wire   [63:0] zext_ln708_116_fu_7689_p1;
wire   [63:0] zext_ln708_117_fu_7704_p1;
wire   [63:0] zext_ln708_118_fu_7719_p1;
wire   [63:0] zext_ln708_119_fu_7734_p1;
wire   [63:0] zext_ln708_120_fu_7749_p1;
wire   [63:0] zext_ln708_121_fu_7764_p1;
wire   [63:0] zext_ln708_122_fu_7779_p1;
wire   [63:0] zext_ln708_123_fu_7794_p1;
wire   [63:0] zext_ln708_124_fu_7809_p1;
wire   [63:0] zext_ln708_125_fu_7824_p1;
wire   [63:0] zext_ln708_126_fu_7839_p1;
wire   [63:0] zext_ln708_127_fu_7854_p1;
wire   [63:0] zext_ln708_128_fu_7869_p1;
wire   [63:0] zext_ln708_129_fu_7884_p1;
wire   [63:0] zext_ln708_130_fu_7899_p1;
wire   [63:0] zext_ln708_131_fu_8736_p1;
wire   [63:0] zext_ln708_132_fu_8741_p1;
wire   [63:0] zext_ln708_133_fu_8746_p1;
wire   [63:0] zext_ln708_134_fu_8751_p1;
wire   [63:0] zext_ln708_135_fu_8756_p1;
wire   [63:0] zext_ln708_136_fu_8761_p1;
wire   [63:0] zext_ln708_137_fu_8766_p1;
wire   [63:0] zext_ln708_138_fu_8771_p1;
wire   [63:0] zext_ln708_139_fu_8776_p1;
wire   [63:0] zext_ln708_140_fu_8781_p1;
wire   [63:0] zext_ln708_141_fu_8786_p1;
wire   [63:0] zext_ln708_142_fu_8791_p1;
wire   [63:0] zext_ln708_143_fu_8796_p1;
wire   [63:0] zext_ln708_144_fu_8801_p1;
wire   [63:0] zext_ln708_145_fu_8806_p1;
wire   [63:0] zext_ln708_146_fu_8811_p1;
wire   [63:0] zext_ln708_147_fu_8861_p1;
wire   [63:0] zext_ln708_148_fu_8876_p1;
wire   [63:0] zext_ln708_149_fu_8891_p1;
wire   [63:0] zext_ln708_150_fu_8906_p1;
wire   [63:0] zext_ln708_151_fu_8921_p1;
wire   [63:0] zext_ln708_152_fu_8936_p1;
wire   [63:0] zext_ln708_153_fu_8951_p1;
wire   [63:0] zext_ln708_154_fu_8966_p1;
wire   [63:0] zext_ln708_155_fu_8981_p1;
wire   [63:0] zext_ln708_156_fu_8996_p1;
wire   [63:0] zext_ln708_157_fu_9011_p1;
wire   [63:0] zext_ln708_158_fu_9026_p1;
wire   [63:0] zext_ln708_159_fu_9041_p1;
wire   [63:0] zext_ln708_160_fu_9056_p1;
wire   [63:0] zext_ln708_161_fu_9071_p1;
wire   [63:0] zext_ln708_162_fu_9086_p1;
wire   [63:0] zext_ln708_163_fu_9923_p1;
wire   [63:0] zext_ln708_164_fu_9928_p1;
wire   [63:0] zext_ln708_165_fu_9933_p1;
wire   [63:0] zext_ln708_166_fu_9938_p1;
wire   [63:0] zext_ln708_167_fu_9943_p1;
wire   [63:0] zext_ln708_168_fu_9948_p1;
wire   [63:0] zext_ln708_169_fu_9953_p1;
wire   [63:0] zext_ln708_170_fu_9958_p1;
wire   [63:0] zext_ln708_171_fu_9963_p1;
wire   [63:0] zext_ln708_172_fu_9968_p1;
wire   [63:0] zext_ln708_173_fu_9973_p1;
wire   [63:0] zext_ln708_174_fu_9978_p1;
wire   [63:0] zext_ln708_175_fu_9983_p1;
wire   [63:0] zext_ln708_176_fu_9988_p1;
wire   [63:0] zext_ln708_177_fu_9993_p1;
wire   [63:0] zext_ln708_178_fu_9998_p1;
wire   [63:0] zext_ln708_179_fu_10048_p1;
wire   [63:0] zext_ln708_180_fu_10063_p1;
wire   [63:0] zext_ln708_181_fu_10078_p1;
wire   [63:0] zext_ln708_182_fu_10093_p1;
wire   [63:0] zext_ln708_183_fu_10108_p1;
wire   [63:0] zext_ln708_184_fu_10123_p1;
wire   [63:0] zext_ln708_185_fu_10138_p1;
wire   [63:0] zext_ln708_186_fu_10153_p1;
wire   [63:0] zext_ln708_187_fu_10168_p1;
wire   [63:0] zext_ln708_188_fu_10183_p1;
wire   [63:0] zext_ln708_189_fu_10198_p1;
wire   [63:0] zext_ln708_190_fu_10213_p1;
wire   [63:0] zext_ln708_191_fu_10228_p1;
wire   [63:0] zext_ln708_192_fu_10243_p1;
wire   [63:0] zext_ln708_193_fu_10258_p1;
wire   [63:0] zext_ln708_194_fu_10273_p1;
wire   [63:0] zext_ln708_195_fu_11110_p1;
wire   [63:0] zext_ln708_196_fu_11115_p1;
wire   [63:0] zext_ln708_197_fu_11120_p1;
wire   [63:0] zext_ln708_198_fu_11125_p1;
wire   [63:0] zext_ln708_199_fu_11130_p1;
wire   [63:0] zext_ln708_200_fu_11135_p1;
wire   [63:0] zext_ln708_201_fu_11140_p1;
wire   [63:0] zext_ln708_202_fu_11145_p1;
wire   [63:0] zext_ln708_203_fu_11150_p1;
wire   [63:0] zext_ln708_204_fu_11155_p1;
wire   [63:0] zext_ln708_205_fu_11160_p1;
wire   [63:0] zext_ln708_206_fu_11165_p1;
wire   [63:0] zext_ln708_207_fu_11170_p1;
wire   [63:0] zext_ln708_208_fu_11175_p1;
wire   [63:0] zext_ln708_209_fu_11180_p1;
wire   [63:0] zext_ln708_210_fu_11185_p1;
wire   [63:0] zext_ln708_211_fu_11235_p1;
wire   [63:0] zext_ln708_212_fu_11250_p1;
wire   [63:0] zext_ln708_213_fu_11265_p1;
wire   [63:0] zext_ln708_214_fu_11280_p1;
wire   [63:0] zext_ln708_215_fu_11295_p1;
wire   [63:0] zext_ln708_216_fu_11310_p1;
wire   [63:0] zext_ln708_217_fu_11325_p1;
wire   [63:0] zext_ln708_218_fu_11340_p1;
wire   [63:0] zext_ln708_219_fu_11355_p1;
wire   [63:0] zext_ln708_220_fu_11370_p1;
wire   [63:0] zext_ln708_221_fu_11385_p1;
wire   [63:0] zext_ln708_222_fu_11400_p1;
wire   [63:0] zext_ln708_223_fu_11415_p1;
wire   [63:0] zext_ln708_224_fu_11430_p1;
wire   [63:0] zext_ln708_225_fu_11445_p1;
wire   [63:0] zext_ln708_226_fu_11460_p1;
wire   [63:0] zext_ln708_227_fu_12297_p1;
wire   [63:0] zext_ln708_228_fu_12302_p1;
wire   [63:0] zext_ln708_229_fu_12307_p1;
wire   [63:0] zext_ln708_230_fu_12312_p1;
wire   [63:0] zext_ln708_231_fu_12317_p1;
wire   [63:0] zext_ln708_232_fu_12322_p1;
wire   [63:0] zext_ln708_233_fu_12327_p1;
wire   [63:0] zext_ln708_234_fu_12332_p1;
wire   [63:0] zext_ln708_235_fu_12337_p1;
wire   [63:0] zext_ln708_236_fu_12342_p1;
wire   [63:0] zext_ln708_237_fu_12347_p1;
wire   [63:0] zext_ln708_238_fu_12352_p1;
wire   [63:0] zext_ln708_239_fu_12357_p1;
wire   [63:0] zext_ln708_240_fu_12362_p1;
wire   [63:0] zext_ln708_241_fu_12367_p1;
wire   [63:0] zext_ln708_242_fu_12372_p1;
wire   [63:0] zext_ln708_243_fu_12422_p1;
wire   [63:0] zext_ln708_244_fu_12437_p1;
wire   [63:0] zext_ln708_245_fu_12452_p1;
wire   [63:0] zext_ln708_246_fu_12467_p1;
wire   [63:0] zext_ln708_247_fu_12482_p1;
wire   [63:0] zext_ln708_248_fu_12497_p1;
wire   [63:0] zext_ln708_249_fu_12512_p1;
wire   [63:0] zext_ln708_250_fu_12527_p1;
wire   [63:0] zext_ln708_251_fu_12542_p1;
wire   [63:0] zext_ln708_252_fu_12557_p1;
wire   [63:0] zext_ln708_253_fu_12572_p1;
wire   [63:0] zext_ln708_254_fu_12587_p1;
wire   [63:0] zext_ln708_255_fu_12602_p1;
wire   [63:0] zext_ln708_256_fu_12617_p1;
wire   [63:0] zext_ln708_257_fu_12632_p1;
wire   [63:0] zext_ln708_258_fu_12647_p1;
wire   [63:0] zext_ln708_259_fu_13484_p1;
wire   [63:0] zext_ln708_260_fu_13489_p1;
wire   [63:0] zext_ln708_261_fu_13494_p1;
wire   [63:0] zext_ln708_262_fu_13499_p1;
wire   [63:0] zext_ln708_263_fu_13504_p1;
wire   [63:0] zext_ln708_264_fu_13509_p1;
wire   [63:0] zext_ln708_265_fu_13514_p1;
wire   [63:0] zext_ln708_266_fu_13519_p1;
wire   [63:0] zext_ln708_267_fu_13524_p1;
wire   [63:0] zext_ln708_268_fu_13529_p1;
wire   [63:0] zext_ln708_269_fu_13534_p1;
wire   [63:0] zext_ln708_270_fu_13539_p1;
wire   [63:0] zext_ln708_271_fu_13544_p1;
wire   [63:0] zext_ln708_272_fu_13549_p1;
wire   [63:0] zext_ln708_273_fu_13554_p1;
wire   [63:0] zext_ln708_274_fu_13559_p1;
wire   [63:0] zext_ln708_275_fu_13609_p1;
wire   [63:0] zext_ln708_276_fu_13624_p1;
wire   [63:0] zext_ln708_277_fu_13639_p1;
wire   [63:0] zext_ln708_278_fu_13654_p1;
wire   [63:0] zext_ln708_279_fu_13669_p1;
wire   [63:0] zext_ln708_280_fu_13684_p1;
wire   [63:0] zext_ln708_281_fu_13699_p1;
wire   [63:0] zext_ln708_282_fu_13714_p1;
wire   [63:0] zext_ln708_283_fu_13729_p1;
wire   [63:0] zext_ln708_284_fu_13744_p1;
wire   [63:0] zext_ln708_285_fu_13759_p1;
wire   [63:0] zext_ln708_286_fu_13774_p1;
wire   [63:0] zext_ln708_287_fu_13789_p1;
wire   [63:0] zext_ln708_288_fu_13804_p1;
wire   [63:0] zext_ln708_289_fu_13819_p1;
wire   [63:0] zext_ln708_290_fu_13834_p1;
wire   [63:0] zext_ln708_291_fu_14671_p1;
wire   [63:0] zext_ln708_292_fu_14676_p1;
wire   [63:0] zext_ln708_293_fu_14681_p1;
wire   [63:0] zext_ln708_294_fu_14686_p1;
wire   [63:0] zext_ln708_295_fu_14691_p1;
wire   [63:0] zext_ln708_296_fu_14696_p1;
wire   [63:0] zext_ln708_297_fu_14701_p1;
wire   [63:0] zext_ln708_298_fu_14706_p1;
wire   [63:0] zext_ln708_299_fu_14711_p1;
wire   [63:0] zext_ln708_300_fu_14716_p1;
wire   [63:0] zext_ln708_301_fu_14721_p1;
wire   [63:0] zext_ln708_302_fu_14726_p1;
wire   [63:0] zext_ln708_303_fu_14731_p1;
wire   [63:0] zext_ln708_304_fu_14736_p1;
wire   [63:0] zext_ln708_305_fu_14741_p1;
wire   [63:0] zext_ln708_306_fu_14746_p1;
wire   [127:0] ret_V_fu_3828_p2;
wire   [7:0] trunc_ln708_fu_3834_p1;
wire   [7:0] tmp_1_fu_3843_p4;
wire   [7:0] tmp_2_fu_3858_p4;
wire   [7:0] tmp_3_fu_3873_p4;
wire   [7:0] tmp_s_fu_3888_p4;
wire   [7:0] tmp_5_fu_3903_p4;
wire   [7:0] tmp_6_fu_3918_p4;
wire   [7:0] tmp_7_fu_3933_p4;
wire   [7:0] tmp_4_fu_3948_p4;
wire   [7:0] tmp_9_fu_3963_p4;
wire   [7:0] tmp_8_fu_3978_p4;
wire   [7:0] tmp_10_fu_3993_p4;
wire   [7:0] tmp_11_fu_4008_p4;
wire   [7:0] tmp_12_fu_4023_p4;
wire   [7:0] tmp_13_fu_4038_p4;
wire   [7:0] tmp_14_fu_4053_p4;
wire   [127:0] p_Result_s_fu_4068_p17;
wire   [127:0] state_V_20_fu_4104_p2;
wire   [7:0] trunc_ln708_1_fu_4109_p1;
wire   [7:0] tmp_18_fu_4118_p4;
wire   [7:0] tmp_22_fu_4133_p4;
wire   [7:0] tmp_26_fu_4148_p4;
wire   [7:0] tmp_30_fu_4163_p4;
wire   [7:0] tmp_34_fu_4178_p4;
wire   [7:0] tmp_38_fu_4193_p4;
wire   [7:0] tmp_42_fu_4208_p4;
wire   [7:0] tmp_46_fu_4223_p4;
wire   [7:0] tmp_50_fu_4238_p4;
wire   [7:0] tmp_54_fu_4253_p4;
wire   [7:0] tmp_58_fu_4268_p4;
wire   [7:0] tmp_62_fu_4283_p4;
wire   [7:0] tmp_66_fu_4298_p4;
wire   [7:0] tmp_70_fu_4313_p4;
wire   [7:0] tmp_74_fu_4328_p4;
wire   [7:0] tmp_19_fu_4381_p4;
wire   [7:0] tmp_17_fu_4367_p4;
wire   [7:0] tmp_24_fu_4425_p4;
wire   [7:0] trunc_ln674_3_fu_4445_p1;
wire   [7:0] xor_ln1545_6_fu_4893_p2;
wire   [7:0] xor_ln1545_fu_4887_p2;
wire   [7:0] tmp_21_fu_4401_p4;
wire   [7:0] trunc_ln674_fu_4343_p1;
wire   [7:0] tmp_23_fu_4415_p4;
wire   [7:0] tmp_28_fu_4459_p4;
wire   [7:0] xor_ln1545_9_fu_4911_p2;
wire   [7:0] xor_ln1545_7_fu_4905_p2;
wire   [7:0] trunc_ln674_1_fu_4377_p1;
wire   [7:0] tmp_16_fu_4357_p4;
wire   [7:0] tmp_25_fu_4435_p4;
wire   [7:0] tmp_27_fu_4449_p4;
wire   [7:0] xor_ln1545_12_fu_4929_p2;
wire   [7:0] xor_ln1545_10_fu_4923_p2;
wire   [7:0] tmp_20_fu_4391_p4;
wire   [7:0] tmp_15_fu_4347_p4;
wire   [7:0] trunc_ln674_2_fu_4411_p1;
wire   [7:0] tmp_29_fu_4469_p4;
wire   [7:0] xor_ln1545_14_fu_4947_p2;
wire   [7:0] xor_ln1545_13_fu_4941_p2;
wire   [7:0] tmp_35_fu_4517_p4;
wire   [7:0] tmp_33_fu_4503_p4;
wire   [7:0] tmp_40_fu_4561_p4;
wire   [7:0] trunc_ln674_7_fu_4581_p1;
wire   [7:0] xor_ln1545_18_fu_4965_p2;
wire   [7:0] xor_ln1545_16_fu_4959_p2;
wire   [7:0] tmp_37_fu_4537_p4;
wire   [7:0] trunc_ln674_4_fu_4479_p1;
wire   [7:0] tmp_39_fu_4551_p4;
wire   [7:0] tmp_44_fu_4595_p4;
wire   [7:0] xor_ln1545_21_fu_4983_p2;
wire   [7:0] xor_ln1545_19_fu_4977_p2;
wire   [7:0] trunc_ln674_5_fu_4513_p1;
wire   [7:0] tmp_32_fu_4493_p4;
wire   [7:0] tmp_41_fu_4571_p4;
wire   [7:0] tmp_43_fu_4585_p4;
wire   [7:0] xor_ln1545_24_fu_5001_p2;
wire   [7:0] xor_ln1545_22_fu_4995_p2;
wire   [7:0] tmp_36_fu_4527_p4;
wire   [7:0] tmp_31_fu_4483_p4;
wire   [7:0] trunc_ln674_6_fu_4547_p1;
wire   [7:0] tmp_45_fu_4605_p4;
wire   [7:0] xor_ln1545_27_fu_5019_p2;
wire   [7:0] xor_ln1545_25_fu_5013_p2;
wire   [7:0] tmp_51_fu_4653_p4;
wire   [7:0] tmp_49_fu_4639_p4;
wire   [7:0] tmp_56_fu_4697_p4;
wire   [7:0] trunc_ln674_11_fu_4717_p1;
wire   [7:0] xor_ln1545_30_fu_5037_p2;
wire   [7:0] xor_ln1545_28_fu_5031_p2;
wire   [7:0] tmp_53_fu_4673_p4;
wire   [7:0] trunc_ln674_8_fu_4615_p1;
wire   [7:0] tmp_55_fu_4687_p4;
wire   [7:0] tmp_60_fu_4731_p4;
wire   [7:0] xor_ln1545_33_fu_5055_p2;
wire   [7:0] xor_ln1545_31_fu_5049_p2;
wire   [7:0] trunc_ln674_9_fu_4649_p1;
wire   [7:0] tmp_48_fu_4629_p4;
wire   [7:0] tmp_57_fu_4707_p4;
wire   [7:0] tmp_59_fu_4721_p4;
wire   [7:0] xor_ln1545_35_fu_5073_p2;
wire   [7:0] xor_ln1545_34_fu_5067_p2;
wire   [7:0] tmp_52_fu_4663_p4;
wire   [7:0] tmp_47_fu_4619_p4;
wire   [7:0] trunc_ln674_10_fu_4683_p1;
wire   [7:0] tmp_61_fu_4741_p4;
wire   [7:0] xor_ln1545_39_fu_5091_p2;
wire   [7:0] xor_ln1545_37_fu_5085_p2;
wire   [7:0] tmp_67_fu_4789_p4;
wire   [7:0] tmp_65_fu_4775_p4;
wire   [7:0] tmp_72_fu_4833_p4;
wire   [7:0] trunc_ln674_15_fu_4853_p1;
wire   [7:0] xor_ln1545_42_fu_5109_p2;
wire   [7:0] xor_ln1545_40_fu_5103_p2;
wire   [7:0] tmp_69_fu_4809_p4;
wire   [7:0] trunc_ln674_12_fu_4751_p1;
wire   [7:0] tmp_71_fu_4823_p4;
wire   [7:0] tmp_76_fu_4867_p4;
wire   [7:0] xor_ln1545_44_fu_5127_p2;
wire   [7:0] xor_ln1545_43_fu_5121_p2;
wire   [7:0] trunc_ln674_13_fu_4785_p1;
wire   [7:0] tmp_64_fu_4765_p4;
wire   [7:0] tmp_73_fu_4843_p4;
wire   [7:0] tmp_75_fu_4857_p4;
wire   [7:0] xor_ln1545_47_fu_5145_p2;
wire   [7:0] xor_ln1545_46_fu_5139_p2;
wire   [7:0] tmp_68_fu_4799_p4;
wire   [7:0] tmp_63_fu_4755_p4;
wire   [7:0] trunc_ln674_14_fu_4819_p1;
wire   [7:0] tmp_77_fu_4877_p4;
wire   [7:0] xor_ln1545_51_fu_5163_p2;
wire   [7:0] xor_ln1545_49_fu_5157_p2;
wire   [7:0] xor_ln1545_5_fu_4899_p2;
wire   [7:0] tmp_1_V_fu_5133_p2;
wire   [7:0] tmp_2_1_V_fu_5079_p2;
wire   [7:0] xor_ln1545_26_fu_5025_p2;
wire   [7:0] xor_ln1545_17_fu_4971_p2;
wire   [7:0] xor_ln1545_8_fu_4917_p2;
wire   [7:0] tmp_2_2_V_fu_5151_p2;
wire   [7:0] xor_ln1545_38_fu_5097_p2;
wire   [7:0] xor_ln1545_29_fu_5043_p2;
wire   [7:0] xor_ln1545_20_fu_4989_p2;
wire   [7:0] xor_ln1545_11_fu_4935_p2;
wire   [7:0] xor_ln1545_50_fu_5169_p2;
wire   [7:0] xor_ln1545_41_fu_5115_p2;
wire   [7:0] xor_ln1545_32_fu_5061_p2;
wire   [7:0] xor_ln1545_23_fu_5007_p2;
wire   [7:0] tmp_3_V_fu_4953_p2;
wire   [127:0] p_Result_2_fu_5255_p17;
wire   [127:0] state_V_21_fu_5291_p2;
wire   [7:0] trunc_ln708_2_fu_5296_p1;
wire   [7:0] tmp_81_fu_5305_p4;
wire   [7:0] tmp_85_fu_5320_p4;
wire   [7:0] tmp_89_fu_5335_p4;
wire   [7:0] tmp_93_fu_5350_p4;
wire   [7:0] tmp_97_fu_5365_p4;
wire   [7:0] tmp_101_fu_5380_p4;
wire   [7:0] tmp_105_fu_5395_p4;
wire   [7:0] tmp_109_fu_5410_p4;
wire   [7:0] tmp_113_fu_5425_p4;
wire   [7:0] tmp_117_fu_5440_p4;
wire   [7:0] tmp_121_fu_5455_p4;
wire   [7:0] tmp_125_fu_5470_p4;
wire   [7:0] tmp_129_fu_5485_p4;
wire   [7:0] tmp_133_fu_5500_p4;
wire   [7:0] tmp_137_fu_5515_p4;
wire   [7:0] tmp_82_fu_5568_p4;
wire   [7:0] tmp_80_fu_5554_p4;
wire   [7:0] tmp_87_fu_5612_p4;
wire   [7:0] trunc_ln674_19_fu_5632_p1;
wire   [7:0] xor_ln1545_54_fu_6080_p2;
wire   [7:0] xor_ln1545_52_fu_6074_p2;
wire   [7:0] tmp_84_fu_5588_p4;
wire   [7:0] trunc_ln674_16_fu_5530_p1;
wire   [7:0] tmp_86_fu_5602_p4;
wire   [7:0] tmp_91_fu_5646_p4;
wire   [7:0] xor_ln1545_57_fu_6098_p2;
wire   [7:0] xor_ln1545_55_fu_6092_p2;
wire   [7:0] trunc_ln674_17_fu_5564_p1;
wire   [7:0] tmp_79_fu_5544_p4;
wire   [7:0] tmp_88_fu_5622_p4;
wire   [7:0] tmp_90_fu_5636_p4;
wire   [7:0] xor_ln1545_60_fu_6116_p2;
wire   [7:0] xor_ln1545_58_fu_6110_p2;
wire   [7:0] tmp_83_fu_5578_p4;
wire   [7:0] tmp_78_fu_5534_p4;
wire   [7:0] trunc_ln674_18_fu_5598_p1;
wire   [7:0] tmp_92_fu_5656_p4;
wire   [7:0] xor_ln1545_62_fu_6134_p2;
wire   [7:0] xor_ln1545_61_fu_6128_p2;
wire   [7:0] tmp_98_fu_5704_p4;
wire   [7:0] tmp_96_fu_5690_p4;
wire   [7:0] tmp_103_fu_5748_p4;
wire   [7:0] trunc_ln674_23_fu_5768_p1;
wire   [7:0] xor_ln1545_66_fu_6152_p2;
wire   [7:0] xor_ln1545_64_fu_6146_p2;
wire   [7:0] tmp_100_fu_5724_p4;
wire   [7:0] trunc_ln674_20_fu_5666_p1;
wire   [7:0] tmp_102_fu_5738_p4;
wire   [7:0] tmp_107_fu_5782_p4;
wire   [7:0] xor_ln1545_69_fu_6170_p2;
wire   [7:0] xor_ln1545_67_fu_6164_p2;
wire   [7:0] trunc_ln674_21_fu_5700_p1;
wire   [7:0] tmp_95_fu_5680_p4;
wire   [7:0] tmp_104_fu_5758_p4;
wire   [7:0] tmp_106_fu_5772_p4;
wire   [7:0] xor_ln1545_72_fu_6188_p2;
wire   [7:0] xor_ln1545_70_fu_6182_p2;
wire   [7:0] tmp_99_fu_5714_p4;
wire   [7:0] tmp_94_fu_5670_p4;
wire   [7:0] trunc_ln674_22_fu_5734_p1;
wire   [7:0] tmp_108_fu_5792_p4;
wire   [7:0] xor_ln1545_75_fu_6206_p2;
wire   [7:0] xor_ln1545_73_fu_6200_p2;
wire   [7:0] tmp_114_fu_5840_p4;
wire   [7:0] tmp_112_fu_5826_p4;
wire   [7:0] tmp_119_fu_5884_p4;
wire   [7:0] trunc_ln674_27_fu_5904_p1;
wire   [7:0] xor_ln1545_78_fu_6224_p2;
wire   [7:0] xor_ln1545_76_fu_6218_p2;
wire   [7:0] tmp_116_fu_5860_p4;
wire   [7:0] trunc_ln674_24_fu_5802_p1;
wire   [7:0] tmp_118_fu_5874_p4;
wire   [7:0] tmp_123_fu_5918_p4;
wire   [7:0] xor_ln1545_81_fu_6242_p2;
wire   [7:0] xor_ln1545_79_fu_6236_p2;
wire   [7:0] trunc_ln674_25_fu_5836_p1;
wire   [7:0] tmp_111_fu_5816_p4;
wire   [7:0] tmp_120_fu_5894_p4;
wire   [7:0] tmp_122_fu_5908_p4;
wire   [7:0] xor_ln1545_83_fu_6260_p2;
wire   [7:0] xor_ln1545_82_fu_6254_p2;
wire   [7:0] tmp_115_fu_5850_p4;
wire   [7:0] tmp_110_fu_5806_p4;
wire   [7:0] trunc_ln674_26_fu_5870_p1;
wire   [7:0] tmp_124_fu_5928_p4;
wire   [7:0] xor_ln1545_87_fu_6278_p2;
wire   [7:0] xor_ln1545_85_fu_6272_p2;
wire   [7:0] tmp_130_fu_5976_p4;
wire   [7:0] tmp_128_fu_5962_p4;
wire   [7:0] tmp_135_fu_6020_p4;
wire   [7:0] trunc_ln674_31_fu_6040_p1;
wire   [7:0] xor_ln1545_90_fu_6296_p2;
wire   [7:0] xor_ln1545_88_fu_6290_p2;
wire   [7:0] tmp_132_fu_5996_p4;
wire   [7:0] trunc_ln674_28_fu_5938_p1;
wire   [7:0] tmp_134_fu_6010_p4;
wire   [7:0] tmp_139_fu_6054_p4;
wire   [7:0] xor_ln1545_92_fu_6314_p2;
wire   [7:0] xor_ln1545_91_fu_6308_p2;
wire   [7:0] trunc_ln674_29_fu_5972_p1;
wire   [7:0] tmp_127_fu_5952_p4;
wire   [7:0] tmp_136_fu_6030_p4;
wire   [7:0] tmp_138_fu_6044_p4;
wire   [7:0] xor_ln1545_95_fu_6332_p2;
wire   [7:0] xor_ln1545_94_fu_6326_p2;
wire   [7:0] tmp_131_fu_5986_p4;
wire   [7:0] tmp_126_fu_5942_p4;
wire   [7:0] trunc_ln674_30_fu_6006_p1;
wire   [7:0] tmp_140_fu_6064_p4;
wire   [7:0] xor_ln1545_99_fu_6350_p2;
wire   [7:0] xor_ln1545_97_fu_6344_p2;
wire   [7:0] xor_ln1545_53_fu_6086_p2;
wire   [7:0] tmp_1_V_1_fu_6320_p2;
wire   [7:0] tmp_2_1_V_1_fu_6266_p2;
wire   [7:0] xor_ln1545_74_fu_6212_p2;
wire   [7:0] xor_ln1545_65_fu_6158_p2;
wire   [7:0] xor_ln1545_56_fu_6104_p2;
wire   [7:0] tmp_2_2_V_1_fu_6338_p2;
wire   [7:0] xor_ln1545_86_fu_6284_p2;
wire   [7:0] xor_ln1545_77_fu_6230_p2;
wire   [7:0] xor_ln1545_68_fu_6176_p2;
wire   [7:0] xor_ln1545_59_fu_6122_p2;
wire   [7:0] xor_ln1545_98_fu_6356_p2;
wire   [7:0] xor_ln1545_89_fu_6302_p2;
wire   [7:0] xor_ln1545_80_fu_6248_p2;
wire   [7:0] xor_ln1545_71_fu_6194_p2;
wire   [7:0] tmp_3_V_1_fu_6140_p2;
wire   [127:0] p_Result_3_fu_6442_p17;
wire   [127:0] state_V_22_fu_6478_p2;
wire   [7:0] trunc_ln708_3_fu_6483_p1;
wire   [7:0] tmp_144_fu_6492_p4;
wire   [7:0] tmp_148_fu_6507_p4;
wire   [7:0] tmp_152_fu_6522_p4;
wire   [7:0] tmp_156_fu_6537_p4;
wire   [7:0] tmp_160_fu_6552_p4;
wire   [7:0] tmp_164_fu_6567_p4;
wire   [7:0] tmp_168_fu_6582_p4;
wire   [7:0] tmp_172_fu_6597_p4;
wire   [7:0] tmp_176_fu_6612_p4;
wire   [7:0] tmp_180_fu_6627_p4;
wire   [7:0] tmp_184_fu_6642_p4;
wire   [7:0] tmp_188_fu_6657_p4;
wire   [7:0] tmp_192_fu_6672_p4;
wire   [7:0] tmp_196_fu_6687_p4;
wire   [7:0] tmp_200_fu_6702_p4;
wire   [7:0] tmp_145_fu_6755_p4;
wire   [7:0] tmp_143_fu_6741_p4;
wire   [7:0] tmp_150_fu_6799_p4;
wire   [7:0] trunc_ln674_35_fu_6819_p1;
wire   [7:0] xor_ln1545_102_fu_7267_p2;
wire   [7:0] xor_ln1545_100_fu_7261_p2;
wire   [7:0] tmp_147_fu_6775_p4;
wire   [7:0] trunc_ln674_32_fu_6717_p1;
wire   [7:0] tmp_149_fu_6789_p4;
wire   [7:0] tmp_154_fu_6833_p4;
wire   [7:0] xor_ln1545_105_fu_7285_p2;
wire   [7:0] xor_ln1545_103_fu_7279_p2;
wire   [7:0] trunc_ln674_33_fu_6751_p1;
wire   [7:0] tmp_142_fu_6731_p4;
wire   [7:0] tmp_151_fu_6809_p4;
wire   [7:0] tmp_153_fu_6823_p4;
wire   [7:0] xor_ln1545_108_fu_7303_p2;
wire   [7:0] xor_ln1545_106_fu_7297_p2;
wire   [7:0] tmp_146_fu_6765_p4;
wire   [7:0] tmp_141_fu_6721_p4;
wire   [7:0] trunc_ln674_34_fu_6785_p1;
wire   [7:0] tmp_155_fu_6843_p4;
wire   [7:0] xor_ln1545_110_fu_7321_p2;
wire   [7:0] xor_ln1545_109_fu_7315_p2;
wire   [7:0] tmp_161_fu_6891_p4;
wire   [7:0] tmp_159_fu_6877_p4;
wire   [7:0] tmp_166_fu_6935_p4;
wire   [7:0] trunc_ln674_39_fu_6955_p1;
wire   [7:0] xor_ln1545_114_fu_7339_p2;
wire   [7:0] xor_ln1545_112_fu_7333_p2;
wire   [7:0] tmp_163_fu_6911_p4;
wire   [7:0] trunc_ln674_36_fu_6853_p1;
wire   [7:0] tmp_165_fu_6925_p4;
wire   [7:0] tmp_170_fu_6969_p4;
wire   [7:0] xor_ln1545_117_fu_7357_p2;
wire   [7:0] xor_ln1545_115_fu_7351_p2;
wire   [7:0] trunc_ln674_37_fu_6887_p1;
wire   [7:0] tmp_158_fu_6867_p4;
wire   [7:0] tmp_167_fu_6945_p4;
wire   [7:0] tmp_169_fu_6959_p4;
wire   [7:0] xor_ln1545_120_fu_7375_p2;
wire   [7:0] xor_ln1545_118_fu_7369_p2;
wire   [7:0] tmp_162_fu_6901_p4;
wire   [7:0] tmp_157_fu_6857_p4;
wire   [7:0] trunc_ln674_38_fu_6921_p1;
wire   [7:0] tmp_171_fu_6979_p4;
wire   [7:0] xor_ln1545_123_fu_7393_p2;
wire   [7:0] xor_ln1545_121_fu_7387_p2;
wire   [7:0] tmp_177_fu_7027_p4;
wire   [7:0] tmp_175_fu_7013_p4;
wire   [7:0] tmp_182_fu_7071_p4;
wire   [7:0] trunc_ln674_43_fu_7091_p1;
wire   [7:0] xor_ln1545_126_fu_7411_p2;
wire   [7:0] xor_ln1545_124_fu_7405_p2;
wire   [7:0] tmp_179_fu_7047_p4;
wire   [7:0] trunc_ln674_40_fu_6989_p1;
wire   [7:0] tmp_181_fu_7061_p4;
wire   [7:0] tmp_186_fu_7105_p4;
wire   [7:0] xor_ln1545_129_fu_7429_p2;
wire   [7:0] xor_ln1545_127_fu_7423_p2;
wire   [7:0] trunc_ln674_41_fu_7023_p1;
wire   [7:0] tmp_174_fu_7003_p4;
wire   [7:0] tmp_183_fu_7081_p4;
wire   [7:0] tmp_185_fu_7095_p4;
wire   [7:0] xor_ln1545_131_fu_7447_p2;
wire   [7:0] xor_ln1545_130_fu_7441_p2;
wire   [7:0] tmp_178_fu_7037_p4;
wire   [7:0] tmp_173_fu_6993_p4;
wire   [7:0] trunc_ln674_42_fu_7057_p1;
wire   [7:0] tmp_187_fu_7115_p4;
wire   [7:0] xor_ln1545_135_fu_7465_p2;
wire   [7:0] xor_ln1545_133_fu_7459_p2;
wire   [7:0] tmp_193_fu_7163_p4;
wire   [7:0] tmp_191_fu_7149_p4;
wire   [7:0] tmp_198_fu_7207_p4;
wire   [7:0] trunc_ln674_47_fu_7227_p1;
wire   [7:0] xor_ln1545_138_fu_7483_p2;
wire   [7:0] xor_ln1545_136_fu_7477_p2;
wire   [7:0] tmp_195_fu_7183_p4;
wire   [7:0] trunc_ln674_44_fu_7125_p1;
wire   [7:0] tmp_197_fu_7197_p4;
wire   [7:0] tmp_202_fu_7241_p4;
wire   [7:0] xor_ln1545_140_fu_7501_p2;
wire   [7:0] xor_ln1545_139_fu_7495_p2;
wire   [7:0] trunc_ln674_45_fu_7159_p1;
wire   [7:0] tmp_190_fu_7139_p4;
wire   [7:0] tmp_199_fu_7217_p4;
wire   [7:0] tmp_201_fu_7231_p4;
wire   [7:0] xor_ln1545_143_fu_7519_p2;
wire   [7:0] xor_ln1545_142_fu_7513_p2;
wire   [7:0] tmp_194_fu_7173_p4;
wire   [7:0] tmp_189_fu_7129_p4;
wire   [7:0] trunc_ln674_46_fu_7193_p1;
wire   [7:0] tmp_203_fu_7251_p4;
wire   [7:0] xor_ln1545_147_fu_7537_p2;
wire   [7:0] xor_ln1545_145_fu_7531_p2;
wire   [7:0] xor_ln1545_101_fu_7273_p2;
wire   [7:0] tmp_1_V_2_fu_7507_p2;
wire   [7:0] tmp_2_1_V_2_fu_7453_p2;
wire   [7:0] xor_ln1545_122_fu_7399_p2;
wire   [7:0] xor_ln1545_113_fu_7345_p2;
wire   [7:0] xor_ln1545_104_fu_7291_p2;
wire   [7:0] tmp_2_2_V_2_fu_7525_p2;
wire   [7:0] xor_ln1545_134_fu_7471_p2;
wire   [7:0] xor_ln1545_125_fu_7417_p2;
wire   [7:0] xor_ln1545_116_fu_7363_p2;
wire   [7:0] xor_ln1545_107_fu_7309_p2;
wire   [7:0] xor_ln1545_146_fu_7543_p2;
wire   [7:0] xor_ln1545_137_fu_7489_p2;
wire   [7:0] xor_ln1545_128_fu_7435_p2;
wire   [7:0] xor_ln1545_119_fu_7381_p2;
wire   [7:0] tmp_3_V_2_fu_7327_p2;
wire   [127:0] p_Result_4_fu_7629_p17;
wire   [127:0] state_V_23_fu_7665_p2;
wire   [7:0] trunc_ln708_4_fu_7670_p1;
wire   [7:0] tmp_207_fu_7679_p4;
wire   [7:0] tmp_211_fu_7694_p4;
wire   [7:0] tmp_215_fu_7709_p4;
wire   [7:0] tmp_219_fu_7724_p4;
wire   [7:0] tmp_223_fu_7739_p4;
wire   [7:0] tmp_227_fu_7754_p4;
wire   [7:0] tmp_231_fu_7769_p4;
wire   [7:0] tmp_235_fu_7784_p4;
wire   [7:0] tmp_239_fu_7799_p4;
wire   [7:0] tmp_243_fu_7814_p4;
wire   [7:0] tmp_247_fu_7829_p4;
wire   [7:0] tmp_251_fu_7844_p4;
wire   [7:0] tmp_255_fu_7859_p4;
wire   [7:0] tmp_259_fu_7874_p4;
wire   [7:0] tmp_263_fu_7889_p4;
wire   [7:0] tmp_208_fu_7942_p4;
wire   [7:0] tmp_206_fu_7928_p4;
wire   [7:0] tmp_213_fu_7986_p4;
wire   [7:0] trunc_ln674_51_fu_8006_p1;
wire   [7:0] xor_ln1545_150_fu_8454_p2;
wire   [7:0] xor_ln1545_148_fu_8448_p2;
wire   [7:0] tmp_210_fu_7962_p4;
wire   [7:0] trunc_ln674_48_fu_7904_p1;
wire   [7:0] tmp_212_fu_7976_p4;
wire   [7:0] tmp_217_fu_8020_p4;
wire   [7:0] xor_ln1545_153_fu_8472_p2;
wire   [7:0] xor_ln1545_151_fu_8466_p2;
wire   [7:0] trunc_ln674_49_fu_7938_p1;
wire   [7:0] tmp_205_fu_7918_p4;
wire   [7:0] tmp_214_fu_7996_p4;
wire   [7:0] tmp_216_fu_8010_p4;
wire   [7:0] xor_ln1545_156_fu_8490_p2;
wire   [7:0] xor_ln1545_154_fu_8484_p2;
wire   [7:0] tmp_209_fu_7952_p4;
wire   [7:0] tmp_204_fu_7908_p4;
wire   [7:0] trunc_ln674_50_fu_7972_p1;
wire   [7:0] tmp_218_fu_8030_p4;
wire   [7:0] xor_ln1545_158_fu_8508_p2;
wire   [7:0] xor_ln1545_157_fu_8502_p2;
wire   [7:0] tmp_224_fu_8078_p4;
wire   [7:0] tmp_222_fu_8064_p4;
wire   [7:0] tmp_229_fu_8122_p4;
wire   [7:0] trunc_ln674_55_fu_8142_p1;
wire   [7:0] xor_ln1545_162_fu_8526_p2;
wire   [7:0] xor_ln1545_160_fu_8520_p2;
wire   [7:0] tmp_226_fu_8098_p4;
wire   [7:0] trunc_ln674_52_fu_8040_p1;
wire   [7:0] tmp_228_fu_8112_p4;
wire   [7:0] tmp_233_fu_8156_p4;
wire   [7:0] xor_ln1545_165_fu_8544_p2;
wire   [7:0] xor_ln1545_163_fu_8538_p2;
wire   [7:0] trunc_ln674_53_fu_8074_p1;
wire   [7:0] tmp_221_fu_8054_p4;
wire   [7:0] tmp_230_fu_8132_p4;
wire   [7:0] tmp_232_fu_8146_p4;
wire   [7:0] xor_ln1545_168_fu_8562_p2;
wire   [7:0] xor_ln1545_166_fu_8556_p2;
wire   [7:0] tmp_225_fu_8088_p4;
wire   [7:0] tmp_220_fu_8044_p4;
wire   [7:0] trunc_ln674_54_fu_8108_p1;
wire   [7:0] tmp_234_fu_8166_p4;
wire   [7:0] xor_ln1545_171_fu_8580_p2;
wire   [7:0] xor_ln1545_169_fu_8574_p2;
wire   [7:0] tmp_240_fu_8214_p4;
wire   [7:0] tmp_238_fu_8200_p4;
wire   [7:0] tmp_245_fu_8258_p4;
wire   [7:0] trunc_ln674_59_fu_8278_p1;
wire   [7:0] xor_ln1545_174_fu_8598_p2;
wire   [7:0] xor_ln1545_172_fu_8592_p2;
wire   [7:0] tmp_242_fu_8234_p4;
wire   [7:0] trunc_ln674_56_fu_8176_p1;
wire   [7:0] tmp_244_fu_8248_p4;
wire   [7:0] tmp_249_fu_8292_p4;
wire   [7:0] xor_ln1545_177_fu_8616_p2;
wire   [7:0] xor_ln1545_175_fu_8610_p2;
wire   [7:0] trunc_ln674_57_fu_8210_p1;
wire   [7:0] tmp_237_fu_8190_p4;
wire   [7:0] tmp_246_fu_8268_p4;
wire   [7:0] tmp_248_fu_8282_p4;
wire   [7:0] xor_ln1545_179_fu_8634_p2;
wire   [7:0] xor_ln1545_178_fu_8628_p2;
wire   [7:0] tmp_241_fu_8224_p4;
wire   [7:0] tmp_236_fu_8180_p4;
wire   [7:0] trunc_ln674_58_fu_8244_p1;
wire   [7:0] tmp_250_fu_8302_p4;
wire   [7:0] xor_ln1545_183_fu_8652_p2;
wire   [7:0] xor_ln1545_181_fu_8646_p2;
wire   [7:0] tmp_256_fu_8350_p4;
wire   [7:0] tmp_254_fu_8336_p4;
wire   [7:0] tmp_261_fu_8394_p4;
wire   [7:0] trunc_ln674_63_fu_8414_p1;
wire   [7:0] xor_ln1545_186_fu_8670_p2;
wire   [7:0] xor_ln1545_184_fu_8664_p2;
wire   [7:0] tmp_258_fu_8370_p4;
wire   [7:0] trunc_ln674_60_fu_8312_p1;
wire   [7:0] tmp_260_fu_8384_p4;
wire   [7:0] tmp_265_fu_8428_p4;
wire   [7:0] xor_ln1545_188_fu_8688_p2;
wire   [7:0] xor_ln1545_187_fu_8682_p2;
wire   [7:0] trunc_ln674_61_fu_8346_p1;
wire   [7:0] tmp_253_fu_8326_p4;
wire   [7:0] tmp_262_fu_8404_p4;
wire   [7:0] tmp_264_fu_8418_p4;
wire   [7:0] xor_ln1545_191_fu_8706_p2;
wire   [7:0] xor_ln1545_190_fu_8700_p2;
wire   [7:0] tmp_257_fu_8360_p4;
wire   [7:0] tmp_252_fu_8316_p4;
wire   [7:0] trunc_ln674_62_fu_8380_p1;
wire   [7:0] tmp_266_fu_8438_p4;
wire   [7:0] xor_ln1545_195_fu_8724_p2;
wire   [7:0] xor_ln1545_193_fu_8718_p2;
wire   [7:0] xor_ln1545_149_fu_8460_p2;
wire   [7:0] tmp_1_V_3_fu_8694_p2;
wire   [7:0] tmp_2_1_V_3_fu_8640_p2;
wire   [7:0] xor_ln1545_170_fu_8586_p2;
wire   [7:0] xor_ln1545_161_fu_8532_p2;
wire   [7:0] xor_ln1545_152_fu_8478_p2;
wire   [7:0] tmp_2_2_V_3_fu_8712_p2;
wire   [7:0] xor_ln1545_182_fu_8658_p2;
wire   [7:0] xor_ln1545_173_fu_8604_p2;
wire   [7:0] xor_ln1545_164_fu_8550_p2;
wire   [7:0] xor_ln1545_155_fu_8496_p2;
wire   [7:0] xor_ln1545_194_fu_8730_p2;
wire   [7:0] xor_ln1545_185_fu_8676_p2;
wire   [7:0] xor_ln1545_176_fu_8622_p2;
wire   [7:0] xor_ln1545_167_fu_8568_p2;
wire   [7:0] tmp_3_V_3_fu_8514_p2;
wire   [127:0] p_Result_5_fu_8816_p17;
wire   [127:0] state_V_24_fu_8852_p2;
wire   [7:0] trunc_ln708_5_fu_8857_p1;
wire   [7:0] tmp_270_fu_8866_p4;
wire   [7:0] tmp_274_fu_8881_p4;
wire   [7:0] tmp_278_fu_8896_p4;
wire   [7:0] tmp_282_fu_8911_p4;
wire   [7:0] tmp_286_fu_8926_p4;
wire   [7:0] tmp_290_fu_8941_p4;
wire   [7:0] tmp_294_fu_8956_p4;
wire   [7:0] tmp_298_fu_8971_p4;
wire   [7:0] tmp_302_fu_8986_p4;
wire   [7:0] tmp_306_fu_9001_p4;
wire   [7:0] tmp_310_fu_9016_p4;
wire   [7:0] tmp_314_fu_9031_p4;
wire   [7:0] tmp_318_fu_9046_p4;
wire   [7:0] tmp_322_fu_9061_p4;
wire   [7:0] tmp_326_fu_9076_p4;
wire   [7:0] tmp_271_fu_9129_p4;
wire   [7:0] tmp_269_fu_9115_p4;
wire   [7:0] tmp_276_fu_9173_p4;
wire   [7:0] trunc_ln674_67_fu_9193_p1;
wire   [7:0] xor_ln1545_198_fu_9641_p2;
wire   [7:0] xor_ln1545_196_fu_9635_p2;
wire   [7:0] tmp_273_fu_9149_p4;
wire   [7:0] trunc_ln674_64_fu_9091_p1;
wire   [7:0] tmp_275_fu_9163_p4;
wire   [7:0] tmp_280_fu_9207_p4;
wire   [7:0] xor_ln1545_201_fu_9659_p2;
wire   [7:0] xor_ln1545_199_fu_9653_p2;
wire   [7:0] trunc_ln674_65_fu_9125_p1;
wire   [7:0] tmp_268_fu_9105_p4;
wire   [7:0] tmp_277_fu_9183_p4;
wire   [7:0] tmp_279_fu_9197_p4;
wire   [7:0] xor_ln1545_204_fu_9677_p2;
wire   [7:0] xor_ln1545_202_fu_9671_p2;
wire   [7:0] tmp_272_fu_9139_p4;
wire   [7:0] tmp_267_fu_9095_p4;
wire   [7:0] trunc_ln674_66_fu_9159_p1;
wire   [7:0] tmp_281_fu_9217_p4;
wire   [7:0] xor_ln1545_206_fu_9695_p2;
wire   [7:0] xor_ln1545_205_fu_9689_p2;
wire   [7:0] tmp_287_fu_9265_p4;
wire   [7:0] tmp_285_fu_9251_p4;
wire   [7:0] tmp_292_fu_9309_p4;
wire   [7:0] trunc_ln674_71_fu_9329_p1;
wire   [7:0] xor_ln1545_210_fu_9713_p2;
wire   [7:0] xor_ln1545_208_fu_9707_p2;
wire   [7:0] tmp_289_fu_9285_p4;
wire   [7:0] trunc_ln674_68_fu_9227_p1;
wire   [7:0] tmp_291_fu_9299_p4;
wire   [7:0] tmp_296_fu_9343_p4;
wire   [7:0] xor_ln1545_213_fu_9731_p2;
wire   [7:0] xor_ln1545_211_fu_9725_p2;
wire   [7:0] trunc_ln674_69_fu_9261_p1;
wire   [7:0] tmp_284_fu_9241_p4;
wire   [7:0] tmp_293_fu_9319_p4;
wire   [7:0] tmp_295_fu_9333_p4;
wire   [7:0] xor_ln1545_216_fu_9749_p2;
wire   [7:0] xor_ln1545_214_fu_9743_p2;
wire   [7:0] tmp_288_fu_9275_p4;
wire   [7:0] tmp_283_fu_9231_p4;
wire   [7:0] trunc_ln674_70_fu_9295_p1;
wire   [7:0] tmp_297_fu_9353_p4;
wire   [7:0] xor_ln1545_219_fu_9767_p2;
wire   [7:0] xor_ln1545_217_fu_9761_p2;
wire   [7:0] tmp_303_fu_9401_p4;
wire   [7:0] tmp_301_fu_9387_p4;
wire   [7:0] tmp_308_fu_9445_p4;
wire   [7:0] trunc_ln674_75_fu_9465_p1;
wire   [7:0] xor_ln1545_222_fu_9785_p2;
wire   [7:0] xor_ln1545_220_fu_9779_p2;
wire   [7:0] tmp_305_fu_9421_p4;
wire   [7:0] trunc_ln674_72_fu_9363_p1;
wire   [7:0] tmp_307_fu_9435_p4;
wire   [7:0] tmp_312_fu_9479_p4;
wire   [7:0] xor_ln1545_225_fu_9803_p2;
wire   [7:0] xor_ln1545_223_fu_9797_p2;
wire   [7:0] trunc_ln674_73_fu_9397_p1;
wire   [7:0] tmp_300_fu_9377_p4;
wire   [7:0] tmp_309_fu_9455_p4;
wire   [7:0] tmp_311_fu_9469_p4;
wire   [7:0] xor_ln1545_227_fu_9821_p2;
wire   [7:0] xor_ln1545_226_fu_9815_p2;
wire   [7:0] tmp_304_fu_9411_p4;
wire   [7:0] tmp_299_fu_9367_p4;
wire   [7:0] trunc_ln674_74_fu_9431_p1;
wire   [7:0] tmp_313_fu_9489_p4;
wire   [7:0] xor_ln1545_231_fu_9839_p2;
wire   [7:0] xor_ln1545_229_fu_9833_p2;
wire   [7:0] tmp_319_fu_9537_p4;
wire   [7:0] tmp_317_fu_9523_p4;
wire   [7:0] tmp_324_fu_9581_p4;
wire   [7:0] trunc_ln674_79_fu_9601_p1;
wire   [7:0] xor_ln1545_234_fu_9857_p2;
wire   [7:0] xor_ln1545_232_fu_9851_p2;
wire   [7:0] tmp_321_fu_9557_p4;
wire   [7:0] trunc_ln674_76_fu_9499_p1;
wire   [7:0] tmp_323_fu_9571_p4;
wire   [7:0] tmp_328_fu_9615_p4;
wire   [7:0] xor_ln1545_236_fu_9875_p2;
wire   [7:0] xor_ln1545_235_fu_9869_p2;
wire   [7:0] trunc_ln674_77_fu_9533_p1;
wire   [7:0] tmp_316_fu_9513_p4;
wire   [7:0] tmp_325_fu_9591_p4;
wire   [7:0] tmp_327_fu_9605_p4;
wire   [7:0] xor_ln1545_239_fu_9893_p2;
wire   [7:0] xor_ln1545_238_fu_9887_p2;
wire   [7:0] tmp_320_fu_9547_p4;
wire   [7:0] tmp_315_fu_9503_p4;
wire   [7:0] trunc_ln674_78_fu_9567_p1;
wire   [7:0] tmp_329_fu_9625_p4;
wire   [7:0] xor_ln1545_243_fu_9911_p2;
wire   [7:0] xor_ln1545_241_fu_9905_p2;
wire   [7:0] xor_ln1545_197_fu_9647_p2;
wire   [7:0] tmp_1_V_4_fu_9881_p2;
wire   [7:0] tmp_2_1_V_4_fu_9827_p2;
wire   [7:0] xor_ln1545_218_fu_9773_p2;
wire   [7:0] xor_ln1545_209_fu_9719_p2;
wire   [7:0] xor_ln1545_200_fu_9665_p2;
wire   [7:0] tmp_2_2_V_4_fu_9899_p2;
wire   [7:0] xor_ln1545_230_fu_9845_p2;
wire   [7:0] xor_ln1545_221_fu_9791_p2;
wire   [7:0] xor_ln1545_212_fu_9737_p2;
wire   [7:0] xor_ln1545_203_fu_9683_p2;
wire   [7:0] xor_ln1545_242_fu_9917_p2;
wire   [7:0] xor_ln1545_233_fu_9863_p2;
wire   [7:0] xor_ln1545_224_fu_9809_p2;
wire   [7:0] xor_ln1545_215_fu_9755_p2;
wire   [7:0] tmp_3_V_4_fu_9701_p2;
wire   [127:0] p_Result_6_fu_10003_p17;
wire   [127:0] state_V_25_fu_10039_p2;
wire   [7:0] trunc_ln708_6_fu_10044_p1;
wire   [7:0] tmp_333_fu_10053_p4;
wire   [7:0] tmp_337_fu_10068_p4;
wire   [7:0] tmp_341_fu_10083_p4;
wire   [7:0] tmp_345_fu_10098_p4;
wire   [7:0] tmp_349_fu_10113_p4;
wire   [7:0] tmp_353_fu_10128_p4;
wire   [7:0] tmp_357_fu_10143_p4;
wire   [7:0] tmp_361_fu_10158_p4;
wire   [7:0] tmp_365_fu_10173_p4;
wire   [7:0] tmp_369_fu_10188_p4;
wire   [7:0] tmp_373_fu_10203_p4;
wire   [7:0] tmp_377_fu_10218_p4;
wire   [7:0] tmp_381_fu_10233_p4;
wire   [7:0] tmp_385_fu_10248_p4;
wire   [7:0] tmp_389_fu_10263_p4;
wire   [7:0] tmp_334_fu_10316_p4;
wire   [7:0] tmp_332_fu_10302_p4;
wire   [7:0] tmp_339_fu_10360_p4;
wire   [7:0] trunc_ln674_83_fu_10380_p1;
wire   [7:0] xor_ln1545_246_fu_10828_p2;
wire   [7:0] xor_ln1545_244_fu_10822_p2;
wire   [7:0] tmp_336_fu_10336_p4;
wire   [7:0] trunc_ln674_80_fu_10278_p1;
wire   [7:0] tmp_338_fu_10350_p4;
wire   [7:0] tmp_343_fu_10394_p4;
wire   [7:0] xor_ln1545_249_fu_10846_p2;
wire   [7:0] xor_ln1545_247_fu_10840_p2;
wire   [7:0] trunc_ln674_81_fu_10312_p1;
wire   [7:0] tmp_331_fu_10292_p4;
wire   [7:0] tmp_340_fu_10370_p4;
wire   [7:0] tmp_342_fu_10384_p4;
wire   [7:0] xor_ln1545_252_fu_10864_p2;
wire   [7:0] xor_ln1545_250_fu_10858_p2;
wire   [7:0] tmp_335_fu_10326_p4;
wire   [7:0] tmp_330_fu_10282_p4;
wire   [7:0] trunc_ln674_82_fu_10346_p1;
wire   [7:0] tmp_344_fu_10404_p4;
wire   [7:0] xor_ln1545_254_fu_10882_p2;
wire   [7:0] xor_ln1545_253_fu_10876_p2;
wire   [7:0] tmp_350_fu_10452_p4;
wire   [7:0] tmp_348_fu_10438_p4;
wire   [7:0] tmp_355_fu_10496_p4;
wire   [7:0] trunc_ln674_87_fu_10516_p1;
wire   [7:0] xor_ln1545_258_fu_10900_p2;
wire   [7:0] xor_ln1545_256_fu_10894_p2;
wire   [7:0] tmp_352_fu_10472_p4;
wire   [7:0] trunc_ln674_84_fu_10414_p1;
wire   [7:0] tmp_354_fu_10486_p4;
wire   [7:0] tmp_359_fu_10530_p4;
wire   [7:0] xor_ln1545_261_fu_10918_p2;
wire   [7:0] xor_ln1545_259_fu_10912_p2;
wire   [7:0] trunc_ln674_85_fu_10448_p1;
wire   [7:0] tmp_347_fu_10428_p4;
wire   [7:0] tmp_356_fu_10506_p4;
wire   [7:0] tmp_358_fu_10520_p4;
wire   [7:0] xor_ln1545_264_fu_10936_p2;
wire   [7:0] xor_ln1545_262_fu_10930_p2;
wire   [7:0] tmp_351_fu_10462_p4;
wire   [7:0] tmp_346_fu_10418_p4;
wire   [7:0] trunc_ln674_86_fu_10482_p1;
wire   [7:0] tmp_360_fu_10540_p4;
wire   [7:0] xor_ln1545_267_fu_10954_p2;
wire   [7:0] xor_ln1545_265_fu_10948_p2;
wire   [7:0] tmp_366_fu_10588_p4;
wire   [7:0] tmp_364_fu_10574_p4;
wire   [7:0] tmp_371_fu_10632_p4;
wire   [7:0] trunc_ln674_91_fu_10652_p1;
wire   [7:0] xor_ln1545_270_fu_10972_p2;
wire   [7:0] xor_ln1545_268_fu_10966_p2;
wire   [7:0] tmp_368_fu_10608_p4;
wire   [7:0] trunc_ln674_88_fu_10550_p1;
wire   [7:0] tmp_370_fu_10622_p4;
wire   [7:0] tmp_375_fu_10666_p4;
wire   [7:0] xor_ln1545_273_fu_10990_p2;
wire   [7:0] xor_ln1545_271_fu_10984_p2;
wire   [7:0] trunc_ln674_89_fu_10584_p1;
wire   [7:0] tmp_363_fu_10564_p4;
wire   [7:0] tmp_372_fu_10642_p4;
wire   [7:0] tmp_374_fu_10656_p4;
wire   [7:0] xor_ln1545_275_fu_11008_p2;
wire   [7:0] xor_ln1545_274_fu_11002_p2;
wire   [7:0] tmp_367_fu_10598_p4;
wire   [7:0] tmp_362_fu_10554_p4;
wire   [7:0] trunc_ln674_90_fu_10618_p1;
wire   [7:0] tmp_376_fu_10676_p4;
wire   [7:0] xor_ln1545_279_fu_11026_p2;
wire   [7:0] xor_ln1545_277_fu_11020_p2;
wire   [7:0] tmp_382_fu_10724_p4;
wire   [7:0] tmp_380_fu_10710_p4;
wire   [7:0] tmp_387_fu_10768_p4;
wire   [7:0] trunc_ln674_95_fu_10788_p1;
wire   [7:0] xor_ln1545_282_fu_11044_p2;
wire   [7:0] xor_ln1545_280_fu_11038_p2;
wire   [7:0] tmp_384_fu_10744_p4;
wire   [7:0] trunc_ln674_92_fu_10686_p1;
wire   [7:0] tmp_386_fu_10758_p4;
wire   [7:0] tmp_391_fu_10802_p4;
wire   [7:0] xor_ln1545_284_fu_11062_p2;
wire   [7:0] xor_ln1545_283_fu_11056_p2;
wire   [7:0] trunc_ln674_93_fu_10720_p1;
wire   [7:0] tmp_379_fu_10700_p4;
wire   [7:0] tmp_388_fu_10778_p4;
wire   [7:0] tmp_390_fu_10792_p4;
wire   [7:0] xor_ln1545_287_fu_11080_p2;
wire   [7:0] xor_ln1545_286_fu_11074_p2;
wire   [7:0] tmp_383_fu_10734_p4;
wire   [7:0] tmp_378_fu_10690_p4;
wire   [7:0] trunc_ln674_94_fu_10754_p1;
wire   [7:0] tmp_392_fu_10812_p4;
wire   [7:0] xor_ln1545_291_fu_11098_p2;
wire   [7:0] xor_ln1545_289_fu_11092_p2;
wire   [7:0] xor_ln1545_245_fu_10834_p2;
wire   [7:0] tmp_1_V_5_fu_11068_p2;
wire   [7:0] tmp_2_1_V_5_fu_11014_p2;
wire   [7:0] xor_ln1545_266_fu_10960_p2;
wire   [7:0] xor_ln1545_257_fu_10906_p2;
wire   [7:0] xor_ln1545_248_fu_10852_p2;
wire   [7:0] tmp_2_2_V_5_fu_11086_p2;
wire   [7:0] xor_ln1545_278_fu_11032_p2;
wire   [7:0] xor_ln1545_269_fu_10978_p2;
wire   [7:0] xor_ln1545_260_fu_10924_p2;
wire   [7:0] xor_ln1545_251_fu_10870_p2;
wire   [7:0] xor_ln1545_290_fu_11104_p2;
wire   [7:0] xor_ln1545_281_fu_11050_p2;
wire   [7:0] xor_ln1545_272_fu_10996_p2;
wire   [7:0] xor_ln1545_263_fu_10942_p2;
wire   [7:0] tmp_3_V_5_fu_10888_p2;
wire   [127:0] p_Result_7_fu_11190_p17;
wire   [127:0] state_V_fu_11226_p2;
wire   [7:0] trunc_ln708_7_fu_11231_p1;
wire   [7:0] tmp_396_fu_11240_p4;
wire   [7:0] tmp_400_fu_11255_p4;
wire   [7:0] tmp_404_fu_11270_p4;
wire   [7:0] tmp_408_fu_11285_p4;
wire   [7:0] tmp_412_fu_11300_p4;
wire   [7:0] tmp_416_fu_11315_p4;
wire   [7:0] tmp_420_fu_11330_p4;
wire   [7:0] tmp_424_fu_11345_p4;
wire   [7:0] tmp_428_fu_11360_p4;
wire   [7:0] tmp_432_fu_11375_p4;
wire   [7:0] tmp_436_fu_11390_p4;
wire   [7:0] tmp_440_fu_11405_p4;
wire   [7:0] tmp_444_fu_11420_p4;
wire   [7:0] tmp_448_fu_11435_p4;
wire   [7:0] tmp_452_fu_11450_p4;
wire   [7:0] tmp_397_fu_11503_p4;
wire   [7:0] tmp_395_fu_11489_p4;
wire   [7:0] tmp_402_fu_11547_p4;
wire   [7:0] trunc_ln674_99_fu_11567_p1;
wire   [7:0] xor_ln1545_294_fu_12015_p2;
wire   [7:0] xor_ln1545_292_fu_12009_p2;
wire   [7:0] tmp_399_fu_11523_p4;
wire   [7:0] trunc_ln674_96_fu_11465_p1;
wire   [7:0] tmp_401_fu_11537_p4;
wire   [7:0] tmp_406_fu_11581_p4;
wire   [7:0] xor_ln1545_297_fu_12033_p2;
wire   [7:0] xor_ln1545_295_fu_12027_p2;
wire   [7:0] trunc_ln674_97_fu_11499_p1;
wire   [7:0] tmp_394_fu_11479_p4;
wire   [7:0] tmp_403_fu_11557_p4;
wire   [7:0] tmp_405_fu_11571_p4;
wire   [7:0] xor_ln1545_300_fu_12051_p2;
wire   [7:0] xor_ln1545_298_fu_12045_p2;
wire   [7:0] tmp_398_fu_11513_p4;
wire   [7:0] tmp_393_fu_11469_p4;
wire   [7:0] trunc_ln674_98_fu_11533_p1;
wire   [7:0] tmp_407_fu_11591_p4;
wire   [7:0] xor_ln1545_302_fu_12069_p2;
wire   [7:0] xor_ln1545_301_fu_12063_p2;
wire   [7:0] tmp_413_fu_11639_p4;
wire   [7:0] tmp_411_fu_11625_p4;
wire   [7:0] tmp_418_fu_11683_p4;
wire   [7:0] trunc_ln674_103_fu_11703_p1;
wire   [7:0] xor_ln1545_306_fu_12087_p2;
wire   [7:0] xor_ln1545_304_fu_12081_p2;
wire   [7:0] tmp_415_fu_11659_p4;
wire   [7:0] trunc_ln674_100_fu_11601_p1;
wire   [7:0] tmp_417_fu_11673_p4;
wire   [7:0] tmp_422_fu_11717_p4;
wire   [7:0] xor_ln1545_309_fu_12105_p2;
wire   [7:0] xor_ln1545_307_fu_12099_p2;
wire   [7:0] trunc_ln674_101_fu_11635_p1;
wire   [7:0] tmp_410_fu_11615_p4;
wire   [7:0] tmp_419_fu_11693_p4;
wire   [7:0] tmp_421_fu_11707_p4;
wire   [7:0] xor_ln1545_312_fu_12123_p2;
wire   [7:0] xor_ln1545_310_fu_12117_p2;
wire   [7:0] tmp_414_fu_11649_p4;
wire   [7:0] tmp_409_fu_11605_p4;
wire   [7:0] trunc_ln674_102_fu_11669_p1;
wire   [7:0] tmp_423_fu_11727_p4;
wire   [7:0] xor_ln1545_315_fu_12141_p2;
wire   [7:0] xor_ln1545_313_fu_12135_p2;
wire   [7:0] tmp_429_fu_11775_p4;
wire   [7:0] tmp_427_fu_11761_p4;
wire   [7:0] tmp_434_fu_11819_p4;
wire   [7:0] trunc_ln674_107_fu_11839_p1;
wire   [7:0] xor_ln1545_318_fu_12159_p2;
wire   [7:0] xor_ln1545_316_fu_12153_p2;
wire   [7:0] tmp_431_fu_11795_p4;
wire   [7:0] trunc_ln674_104_fu_11737_p1;
wire   [7:0] tmp_433_fu_11809_p4;
wire   [7:0] tmp_438_fu_11853_p4;
wire   [7:0] xor_ln1545_321_fu_12177_p2;
wire   [7:0] xor_ln1545_319_fu_12171_p2;
wire   [7:0] trunc_ln674_105_fu_11771_p1;
wire   [7:0] tmp_426_fu_11751_p4;
wire   [7:0] tmp_435_fu_11829_p4;
wire   [7:0] tmp_437_fu_11843_p4;
wire   [7:0] xor_ln1545_323_fu_12195_p2;
wire   [7:0] xor_ln1545_322_fu_12189_p2;
wire   [7:0] tmp_430_fu_11785_p4;
wire   [7:0] tmp_425_fu_11741_p4;
wire   [7:0] trunc_ln674_106_fu_11805_p1;
wire   [7:0] tmp_439_fu_11863_p4;
wire   [7:0] xor_ln1545_327_fu_12213_p2;
wire   [7:0] xor_ln1545_325_fu_12207_p2;
wire   [7:0] tmp_445_fu_11911_p4;
wire   [7:0] tmp_443_fu_11897_p4;
wire   [7:0] tmp_450_fu_11955_p4;
wire   [7:0] trunc_ln674_111_fu_11975_p1;
wire   [7:0] xor_ln1545_330_fu_12231_p2;
wire   [7:0] xor_ln1545_328_fu_12225_p2;
wire   [7:0] tmp_447_fu_11931_p4;
wire   [7:0] trunc_ln674_108_fu_11873_p1;
wire   [7:0] tmp_449_fu_11945_p4;
wire   [7:0] tmp_454_fu_11989_p4;
wire   [7:0] xor_ln1545_332_fu_12249_p2;
wire   [7:0] xor_ln1545_331_fu_12243_p2;
wire   [7:0] trunc_ln674_109_fu_11907_p1;
wire   [7:0] tmp_442_fu_11887_p4;
wire   [7:0] tmp_451_fu_11965_p4;
wire   [7:0] tmp_453_fu_11979_p4;
wire   [7:0] xor_ln1545_335_fu_12267_p2;
wire   [7:0] xor_ln1545_334_fu_12261_p2;
wire   [7:0] tmp_446_fu_11921_p4;
wire   [7:0] tmp_441_fu_11877_p4;
wire   [7:0] trunc_ln674_110_fu_11941_p1;
wire   [7:0] tmp_455_fu_11999_p4;
wire   [7:0] xor_ln1545_339_fu_12285_p2;
wire   [7:0] xor_ln1545_337_fu_12279_p2;
wire   [7:0] xor_ln1545_293_fu_12021_p2;
wire   [7:0] tmp_1_V_6_fu_12255_p2;
wire   [7:0] tmp_2_1_V_6_fu_12201_p2;
wire   [7:0] xor_ln1545_314_fu_12147_p2;
wire   [7:0] xor_ln1545_305_fu_12093_p2;
wire   [7:0] xor_ln1545_296_fu_12039_p2;
wire   [7:0] tmp_2_2_V_6_fu_12273_p2;
wire   [7:0] xor_ln1545_326_fu_12219_p2;
wire   [7:0] xor_ln1545_317_fu_12165_p2;
wire   [7:0] xor_ln1545_308_fu_12111_p2;
wire   [7:0] xor_ln1545_299_fu_12057_p2;
wire   [7:0] xor_ln1545_338_fu_12291_p2;
wire   [7:0] xor_ln1545_329_fu_12237_p2;
wire   [7:0] xor_ln1545_320_fu_12183_p2;
wire   [7:0] xor_ln1545_311_fu_12129_p2;
wire   [7:0] tmp_3_V_6_fu_12075_p2;
wire   [127:0] p_Result_8_fu_12377_p17;
wire   [127:0] state_V_26_fu_12413_p2;
wire   [7:0] trunc_ln708_8_fu_12418_p1;
wire   [7:0] tmp_459_fu_12427_p4;
wire   [7:0] tmp_463_fu_12442_p4;
wire   [7:0] tmp_467_fu_12457_p4;
wire   [7:0] tmp_471_fu_12472_p4;
wire   [7:0] tmp_475_fu_12487_p4;
wire   [7:0] tmp_479_fu_12502_p4;
wire   [7:0] tmp_483_fu_12517_p4;
wire   [7:0] tmp_487_fu_12532_p4;
wire   [7:0] tmp_491_fu_12547_p4;
wire   [7:0] tmp_495_fu_12562_p4;
wire   [7:0] tmp_499_fu_12577_p4;
wire   [7:0] tmp_503_fu_12592_p4;
wire   [7:0] tmp_507_fu_12607_p4;
wire   [7:0] tmp_511_fu_12622_p4;
wire   [7:0] tmp_515_fu_12637_p4;
wire   [7:0] tmp_460_fu_12690_p4;
wire   [7:0] tmp_458_fu_12676_p4;
wire   [7:0] tmp_465_fu_12734_p4;
wire   [7:0] trunc_ln674_115_fu_12754_p1;
wire   [7:0] xor_ln1545_342_fu_13202_p2;
wire   [7:0] xor_ln1545_340_fu_13196_p2;
wire   [7:0] tmp_462_fu_12710_p4;
wire   [7:0] trunc_ln674_112_fu_12652_p1;
wire   [7:0] tmp_464_fu_12724_p4;
wire   [7:0] tmp_469_fu_12768_p4;
wire   [7:0] xor_ln1545_345_fu_13220_p2;
wire   [7:0] xor_ln1545_343_fu_13214_p2;
wire   [7:0] trunc_ln674_113_fu_12686_p1;
wire   [7:0] tmp_457_fu_12666_p4;
wire   [7:0] tmp_466_fu_12744_p4;
wire   [7:0] tmp_468_fu_12758_p4;
wire   [7:0] xor_ln1545_348_fu_13238_p2;
wire   [7:0] xor_ln1545_346_fu_13232_p2;
wire   [7:0] tmp_461_fu_12700_p4;
wire   [7:0] tmp_456_fu_12656_p4;
wire   [7:0] trunc_ln674_114_fu_12720_p1;
wire   [7:0] tmp_470_fu_12778_p4;
wire   [7:0] xor_ln1545_350_fu_13256_p2;
wire   [7:0] xor_ln1545_349_fu_13250_p2;
wire   [7:0] tmp_476_fu_12826_p4;
wire   [7:0] tmp_474_fu_12812_p4;
wire   [7:0] tmp_481_fu_12870_p4;
wire   [7:0] trunc_ln674_119_fu_12890_p1;
wire   [7:0] xor_ln1545_354_fu_13274_p2;
wire   [7:0] xor_ln1545_352_fu_13268_p2;
wire   [7:0] tmp_478_fu_12846_p4;
wire   [7:0] trunc_ln674_116_fu_12788_p1;
wire   [7:0] tmp_480_fu_12860_p4;
wire   [7:0] tmp_485_fu_12904_p4;
wire   [7:0] xor_ln1545_357_fu_13292_p2;
wire   [7:0] xor_ln1545_355_fu_13286_p2;
wire   [7:0] trunc_ln674_117_fu_12822_p1;
wire   [7:0] tmp_473_fu_12802_p4;
wire   [7:0] tmp_482_fu_12880_p4;
wire   [7:0] tmp_484_fu_12894_p4;
wire   [7:0] xor_ln1545_360_fu_13310_p2;
wire   [7:0] xor_ln1545_358_fu_13304_p2;
wire   [7:0] tmp_477_fu_12836_p4;
wire   [7:0] tmp_472_fu_12792_p4;
wire   [7:0] trunc_ln674_118_fu_12856_p1;
wire   [7:0] tmp_486_fu_12914_p4;
wire   [7:0] xor_ln1545_363_fu_13328_p2;
wire   [7:0] xor_ln1545_361_fu_13322_p2;
wire   [7:0] tmp_492_fu_12962_p4;
wire   [7:0] tmp_490_fu_12948_p4;
wire   [7:0] tmp_497_fu_13006_p4;
wire   [7:0] trunc_ln674_123_fu_13026_p1;
wire   [7:0] xor_ln1545_366_fu_13346_p2;
wire   [7:0] xor_ln1545_364_fu_13340_p2;
wire   [7:0] tmp_494_fu_12982_p4;
wire   [7:0] trunc_ln674_120_fu_12924_p1;
wire   [7:0] tmp_496_fu_12996_p4;
wire   [7:0] tmp_501_fu_13040_p4;
wire   [7:0] xor_ln1545_369_fu_13364_p2;
wire   [7:0] xor_ln1545_367_fu_13358_p2;
wire   [7:0] trunc_ln674_121_fu_12958_p1;
wire   [7:0] tmp_489_fu_12938_p4;
wire   [7:0] tmp_498_fu_13016_p4;
wire   [7:0] tmp_500_fu_13030_p4;
wire   [7:0] xor_ln1545_371_fu_13382_p2;
wire   [7:0] xor_ln1545_370_fu_13376_p2;
wire   [7:0] tmp_493_fu_12972_p4;
wire   [7:0] tmp_488_fu_12928_p4;
wire   [7:0] trunc_ln674_122_fu_12992_p1;
wire   [7:0] tmp_502_fu_13050_p4;
wire   [7:0] xor_ln1545_375_fu_13400_p2;
wire   [7:0] xor_ln1545_373_fu_13394_p2;
wire   [7:0] tmp_508_fu_13098_p4;
wire   [7:0] tmp_506_fu_13084_p4;
wire   [7:0] tmp_513_fu_13142_p4;
wire   [7:0] trunc_ln674_127_fu_13162_p1;
wire   [7:0] xor_ln1545_378_fu_13418_p2;
wire   [7:0] xor_ln1545_376_fu_13412_p2;
wire   [7:0] tmp_510_fu_13118_p4;
wire   [7:0] trunc_ln674_124_fu_13060_p1;
wire   [7:0] tmp_512_fu_13132_p4;
wire   [7:0] tmp_517_fu_13176_p4;
wire   [7:0] xor_ln1545_380_fu_13436_p2;
wire   [7:0] xor_ln1545_379_fu_13430_p2;
wire   [7:0] trunc_ln674_125_fu_13094_p1;
wire   [7:0] tmp_505_fu_13074_p4;
wire   [7:0] tmp_514_fu_13152_p4;
wire   [7:0] tmp_516_fu_13166_p4;
wire   [7:0] xor_ln1545_383_fu_13454_p2;
wire   [7:0] xor_ln1545_382_fu_13448_p2;
wire   [7:0] tmp_509_fu_13108_p4;
wire   [7:0] tmp_504_fu_13064_p4;
wire   [7:0] trunc_ln674_126_fu_13128_p1;
wire   [7:0] tmp_518_fu_13186_p4;
wire   [7:0] xor_ln1545_387_fu_13472_p2;
wire   [7:0] xor_ln1545_385_fu_13466_p2;
wire   [7:0] xor_ln1545_341_fu_13208_p2;
wire   [7:0] tmp_1_V_7_fu_13442_p2;
wire   [7:0] tmp_2_1_V_7_fu_13388_p2;
wire   [7:0] xor_ln1545_362_fu_13334_p2;
wire   [7:0] xor_ln1545_353_fu_13280_p2;
wire   [7:0] xor_ln1545_344_fu_13226_p2;
wire   [7:0] tmp_2_2_V_7_fu_13460_p2;
wire   [7:0] xor_ln1545_374_fu_13406_p2;
wire   [7:0] xor_ln1545_365_fu_13352_p2;
wire   [7:0] xor_ln1545_356_fu_13298_p2;
wire   [7:0] xor_ln1545_347_fu_13244_p2;
wire   [7:0] xor_ln1545_386_fu_13478_p2;
wire   [7:0] xor_ln1545_377_fu_13424_p2;
wire   [7:0] xor_ln1545_368_fu_13370_p2;
wire   [7:0] xor_ln1545_359_fu_13316_p2;
wire   [7:0] tmp_3_V_7_fu_13262_p2;
wire   [127:0] p_Result_9_fu_13564_p17;
wire   [127:0] state_V_27_fu_13600_p2;
wire   [7:0] trunc_ln708_9_fu_13605_p1;
wire   [7:0] tmp_522_fu_13614_p4;
wire   [7:0] tmp_526_fu_13629_p4;
wire   [7:0] tmp_530_fu_13644_p4;
wire   [7:0] tmp_534_fu_13659_p4;
wire   [7:0] tmp_538_fu_13674_p4;
wire   [7:0] tmp_542_fu_13689_p4;
wire   [7:0] tmp_546_fu_13704_p4;
wire   [7:0] tmp_550_fu_13719_p4;
wire   [7:0] tmp_554_fu_13734_p4;
wire   [7:0] tmp_558_fu_13749_p4;
wire   [7:0] tmp_562_fu_13764_p4;
wire   [7:0] tmp_566_fu_13779_p4;
wire   [7:0] tmp_570_fu_13794_p4;
wire   [7:0] tmp_574_fu_13809_p4;
wire   [7:0] tmp_578_fu_13824_p4;
wire   [7:0] tmp_523_fu_13877_p4;
wire   [7:0] tmp_521_fu_13863_p4;
wire   [7:0] tmp_528_fu_13921_p4;
wire   [7:0] trunc_ln674_131_fu_13941_p1;
wire   [7:0] xor_ln1545_390_fu_14389_p2;
wire   [7:0] xor_ln1545_388_fu_14383_p2;
wire   [7:0] tmp_525_fu_13897_p4;
wire   [7:0] trunc_ln674_128_fu_13839_p1;
wire   [7:0] tmp_527_fu_13911_p4;
wire   [7:0] tmp_532_fu_13955_p4;
wire   [7:0] xor_ln1545_393_fu_14407_p2;
wire   [7:0] xor_ln1545_391_fu_14401_p2;
wire   [7:0] trunc_ln674_129_fu_13873_p1;
wire   [7:0] tmp_520_fu_13853_p4;
wire   [7:0] tmp_529_fu_13931_p4;
wire   [7:0] tmp_531_fu_13945_p4;
wire   [7:0] xor_ln1545_396_fu_14425_p2;
wire   [7:0] xor_ln1545_394_fu_14419_p2;
wire   [7:0] tmp_524_fu_13887_p4;
wire   [7:0] tmp_519_fu_13843_p4;
wire   [7:0] trunc_ln674_130_fu_13907_p1;
wire   [7:0] tmp_533_fu_13965_p4;
wire   [7:0] xor_ln1545_398_fu_14443_p2;
wire   [7:0] xor_ln1545_397_fu_14437_p2;
wire   [7:0] tmp_539_fu_14013_p4;
wire   [7:0] tmp_537_fu_13999_p4;
wire   [7:0] tmp_544_fu_14057_p4;
wire   [7:0] trunc_ln674_135_fu_14077_p1;
wire   [7:0] xor_ln1545_402_fu_14461_p2;
wire   [7:0] xor_ln1545_400_fu_14455_p2;
wire   [7:0] tmp_541_fu_14033_p4;
wire   [7:0] trunc_ln674_132_fu_13975_p1;
wire   [7:0] tmp_543_fu_14047_p4;
wire   [7:0] tmp_548_fu_14091_p4;
wire   [7:0] xor_ln1545_405_fu_14479_p2;
wire   [7:0] xor_ln1545_403_fu_14473_p2;
wire   [7:0] trunc_ln674_133_fu_14009_p1;
wire   [7:0] tmp_536_fu_13989_p4;
wire   [7:0] tmp_545_fu_14067_p4;
wire   [7:0] tmp_547_fu_14081_p4;
wire   [7:0] xor_ln1545_408_fu_14497_p2;
wire   [7:0] xor_ln1545_406_fu_14491_p2;
wire   [7:0] tmp_540_fu_14023_p4;
wire   [7:0] tmp_535_fu_13979_p4;
wire   [7:0] trunc_ln674_134_fu_14043_p1;
wire   [7:0] tmp_549_fu_14101_p4;
wire   [7:0] xor_ln1545_411_fu_14515_p2;
wire   [7:0] xor_ln1545_409_fu_14509_p2;
wire   [7:0] tmp_555_fu_14149_p4;
wire   [7:0] tmp_553_fu_14135_p4;
wire   [7:0] tmp_560_fu_14193_p4;
wire   [7:0] trunc_ln674_139_fu_14213_p1;
wire   [7:0] xor_ln1545_414_fu_14533_p2;
wire   [7:0] xor_ln1545_412_fu_14527_p2;
wire   [7:0] tmp_557_fu_14169_p4;
wire   [7:0] trunc_ln674_136_fu_14111_p1;
wire   [7:0] tmp_559_fu_14183_p4;
wire   [7:0] tmp_564_fu_14227_p4;
wire   [7:0] xor_ln1545_417_fu_14551_p2;
wire   [7:0] xor_ln1545_415_fu_14545_p2;
wire   [7:0] trunc_ln674_137_fu_14145_p1;
wire   [7:0] tmp_552_fu_14125_p4;
wire   [7:0] tmp_561_fu_14203_p4;
wire   [7:0] tmp_563_fu_14217_p4;
wire   [7:0] xor_ln1545_419_fu_14569_p2;
wire   [7:0] xor_ln1545_418_fu_14563_p2;
wire   [7:0] tmp_556_fu_14159_p4;
wire   [7:0] tmp_551_fu_14115_p4;
wire   [7:0] trunc_ln674_138_fu_14179_p1;
wire   [7:0] tmp_565_fu_14237_p4;
wire   [7:0] xor_ln1545_423_fu_14587_p2;
wire   [7:0] xor_ln1545_421_fu_14581_p2;
wire   [7:0] tmp_571_fu_14285_p4;
wire   [7:0] tmp_569_fu_14271_p4;
wire   [7:0] tmp_576_fu_14329_p4;
wire   [7:0] trunc_ln674_143_fu_14349_p1;
wire   [7:0] xor_ln1545_426_fu_14605_p2;
wire   [7:0] xor_ln1545_424_fu_14599_p2;
wire   [7:0] tmp_573_fu_14305_p4;
wire   [7:0] trunc_ln674_140_fu_14247_p1;
wire   [7:0] tmp_575_fu_14319_p4;
wire   [7:0] tmp_580_fu_14363_p4;
wire   [7:0] xor_ln1545_428_fu_14623_p2;
wire   [7:0] xor_ln1545_427_fu_14617_p2;
wire   [7:0] trunc_ln674_141_fu_14281_p1;
wire   [7:0] tmp_568_fu_14261_p4;
wire   [7:0] tmp_577_fu_14339_p4;
wire   [7:0] tmp_579_fu_14353_p4;
wire   [7:0] xor_ln1545_431_fu_14641_p2;
wire   [7:0] xor_ln1545_430_fu_14635_p2;
wire   [7:0] tmp_572_fu_14295_p4;
wire   [7:0] tmp_567_fu_14251_p4;
wire   [7:0] trunc_ln674_142_fu_14315_p1;
wire   [7:0] tmp_581_fu_14373_p4;
wire   [7:0] xor_ln1545_435_fu_14659_p2;
wire   [7:0] xor_ln1545_433_fu_14653_p2;
wire   [7:0] xor_ln1545_389_fu_14395_p2;
wire   [7:0] tmp_1_V_8_fu_14629_p2;
wire   [7:0] tmp_2_1_V_8_fu_14575_p2;
wire   [7:0] xor_ln1545_410_fu_14521_p2;
wire   [7:0] xor_ln1545_401_fu_14467_p2;
wire   [7:0] xor_ln1545_392_fu_14413_p2;
wire   [7:0] tmp_2_2_V_8_fu_14647_p2;
wire   [7:0] xor_ln1545_422_fu_14593_p2;
wire   [7:0] xor_ln1545_413_fu_14539_p2;
wire   [7:0] xor_ln1545_404_fu_14485_p2;
wire   [7:0] xor_ln1545_395_fu_14431_p2;
wire   [7:0] xor_ln1545_434_fu_14665_p2;
wire   [7:0] xor_ln1545_425_fu_14611_p2;
wire   [7:0] xor_ln1545_416_fu_14557_p2;
wire   [7:0] xor_ln1545_407_fu_14503_p2;
wire   [7:0] tmp_3_V_8_fu_14449_p2;
wire   [127:0] p_Result_10_fu_14751_p17;
reg   [0:0] ap_NS_fsm;
reg    ap_idle_pp0_0to18;
reg    ap_reset_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 1'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter5 = 1'b0;
#0 ap_enable_reg_pp0_iter6 = 1'b0;
#0 ap_enable_reg_pp0_iter7 = 1'b0;
#0 ap_enable_reg_pp0_iter8 = 1'b0;
#0 ap_enable_reg_pp0_iter9 = 1'b0;
#0 ap_enable_reg_pp0_iter10 = 1'b0;
#0 ap_enable_reg_pp0_iter11 = 1'b0;
#0 ap_enable_reg_pp0_iter12 = 1'b0;
#0 ap_enable_reg_pp0_iter13 = 1'b0;
#0 ap_enable_reg_pp0_iter14 = 1'b0;
#0 ap_enable_reg_pp0_iter15 = 1'b0;
#0 ap_enable_reg_pp0_iter16 = 1'b0;
#0 ap_enable_reg_pp0_iter17 = 1'b0;
#0 ap_enable_reg_pp0_iter18 = 1'b0;
#0 ap_enable_reg_pp0_iter19 = 1'b0;
end

testDec_process_r_decipher_0_iibox_ROM_NP_LUTRAM_1R #(
    .DataWidth( 8 ),
    .AddressRange( 256 ),
    .AddressWidth( 8 ))
decipher_0_iibox_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(decipher_0_iibox_address0),
    .ce0(decipher_0_iibox_ce0),
    .q0(decipher_0_iibox_q0),
    .address1(decipher_0_iibox_address1),
    .ce1(decipher_0_iibox_ce1),
    .q1(decipher_0_iibox_q1),
    .address2(decipher_0_iibox_address2),
    .ce2(decipher_0_iibox_ce2),
    .q2(decipher_0_iibox_q2),
    .address3(decipher_0_iibox_address3),
    .ce3(decipher_0_iibox_ce3),
    .q3(decipher_0_iibox_q3),
    .address4(decipher_0_iibox_address4),
    .ce4(decipher_0_iibox_ce4),
    .q4(decipher_0_iibox_q4),
    .address5(decipher_0_iibox_address5),
    .ce5(decipher_0_iibox_ce5),
    .q5(decipher_0_iibox_q5),
    .address6(decipher_0_iibox_address6),
    .ce6(decipher_0_iibox_ce6),
    .q6(decipher_0_iibox_q6),
    .address7(decipher_0_iibox_address7),
    .ce7(decipher_0_iibox_ce7),
    .q7(decipher_0_iibox_q7),
    .address8(decipher_0_iibox_address8),
    .ce8(decipher_0_iibox_ce8),
    .q8(decipher_0_iibox_q8),
    .address9(decipher_0_iibox_address9),
    .ce9(decipher_0_iibox_ce9),
    .q9(decipher_0_iibox_q9),
    .address10(decipher_0_iibox_address10),
    .ce10(decipher_0_iibox_ce10),
    .q10(decipher_0_iibox_q10),
    .address11(decipher_0_iibox_address11),
    .ce11(decipher_0_iibox_ce11),
    .q11(decipher_0_iibox_q11),
    .address12(decipher_0_iibox_address12),
    .ce12(decipher_0_iibox_ce12),
    .q12(decipher_0_iibox_q12),
    .address13(decipher_0_iibox_address13),
    .ce13(decipher_0_iibox_ce13),
    .q13(decipher_0_iibox_q13),
    .address14(decipher_0_iibox_address14),
    .ce14(decipher_0_iibox_ce14),
    .q14(decipher_0_iibox_q14),
    .address15(decipher_0_iibox_address15),
    .ce15(decipher_0_iibox_ce15),
    .q15(decipher_0_iibox_q15),
    .address16(decipher_0_iibox_address16),
    .ce16(decipher_0_iibox_ce16),
    .q16(decipher_0_iibox_q16),
    .address17(decipher_0_iibox_address17),
    .ce17(decipher_0_iibox_ce17),
    .q17(decipher_0_iibox_q17),
    .address18(decipher_0_iibox_address18),
    .ce18(decipher_0_iibox_ce18),
    .q18(decipher_0_iibox_q18),
    .address19(decipher_0_iibox_address19),
    .ce19(decipher_0_iibox_ce19),
    .q19(decipher_0_iibox_q19),
    .address20(decipher_0_iibox_address20),
    .ce20(decipher_0_iibox_ce20),
    .q20(decipher_0_iibox_q20),
    .address21(decipher_0_iibox_address21),
    .ce21(decipher_0_iibox_ce21),
    .q21(decipher_0_iibox_q21),
    .address22(decipher_0_iibox_address22),
    .ce22(decipher_0_iibox_ce22),
    .q22(decipher_0_iibox_q22),
    .address23(decipher_0_iibox_address23),
    .ce23(decipher_0_iibox_ce23),
    .q23(decipher_0_iibox_q23),
    .address24(decipher_0_iibox_address24),
    .ce24(decipher_0_iibox_ce24),
    .q24(decipher_0_iibox_q24),
    .address25(decipher_0_iibox_address25),
    .ce25(decipher_0_iibox_ce25),
    .q25(decipher_0_iibox_q25),
    .address26(decipher_0_iibox_address26),
    .ce26(decipher_0_iibox_ce26),
    .q26(decipher_0_iibox_q26),
    .address27(decipher_0_iibox_address27),
    .ce27(decipher_0_iibox_ce27),
    .q27(decipher_0_iibox_q27),
    .address28(decipher_0_iibox_address28),
    .ce28(decipher_0_iibox_ce28),
    .q28(decipher_0_iibox_q28),
    .address29(decipher_0_iibox_address29),
    .ce29(decipher_0_iibox_ce29),
    .q29(decipher_0_iibox_q29),
    .address30(decipher_0_iibox_address30),
    .ce30(decipher_0_iibox_ce30),
    .q30(decipher_0_iibox_q30),
    .address31(decipher_0_iibox_address31),
    .ce31(decipher_0_iibox_ce31),
    .q31(decipher_0_iibox_q31),
    .address32(decipher_0_iibox_address32),
    .ce32(decipher_0_iibox_ce32),
    .q32(decipher_0_iibox_q32),
    .address33(decipher_0_iibox_address33),
    .ce33(decipher_0_iibox_ce33),
    .q33(decipher_0_iibox_q33),
    .address34(decipher_0_iibox_address34),
    .ce34(decipher_0_iibox_ce34),
    .q34(decipher_0_iibox_q34),
    .address35(decipher_0_iibox_address35),
    .ce35(decipher_0_iibox_ce35),
    .q35(decipher_0_iibox_q35),
    .address36(decipher_0_iibox_address36),
    .ce36(decipher_0_iibox_ce36),
    .q36(decipher_0_iibox_q36),
    .address37(decipher_0_iibox_address37),
    .ce37(decipher_0_iibox_ce37),
    .q37(decipher_0_iibox_q37),
    .address38(decipher_0_iibox_address38),
    .ce38(decipher_0_iibox_ce38),
    .q38(decipher_0_iibox_q38),
    .address39(decipher_0_iibox_address39),
    .ce39(decipher_0_iibox_ce39),
    .q39(decipher_0_iibox_q39),
    .address40(decipher_0_iibox_address40),
    .ce40(decipher_0_iibox_ce40),
    .q40(decipher_0_iibox_q40),
    .address41(decipher_0_iibox_address41),
    .ce41(decipher_0_iibox_ce41),
    .q41(decipher_0_iibox_q41),
    .address42(decipher_0_iibox_address42),
    .ce42(decipher_0_iibox_ce42),
    .q42(decipher_0_iibox_q42),
    .address43(decipher_0_iibox_address43),
    .ce43(decipher_0_iibox_ce43),
    .q43(decipher_0_iibox_q43),
    .address44(decipher_0_iibox_address44),
    .ce44(decipher_0_iibox_ce44),
    .q44(decipher_0_iibox_q44),
    .address45(decipher_0_iibox_address45),
    .ce45(decipher_0_iibox_ce45),
    .q45(decipher_0_iibox_q45),
    .address46(decipher_0_iibox_address46),
    .ce46(decipher_0_iibox_ce46),
    .q46(decipher_0_iibox_q46),
    .address47(decipher_0_iibox_address47),
    .ce47(decipher_0_iibox_ce47),
    .q47(decipher_0_iibox_q47),
    .address48(decipher_0_iibox_address48),
    .ce48(decipher_0_iibox_ce48),
    .q48(decipher_0_iibox_q48),
    .address49(decipher_0_iibox_address49),
    .ce49(decipher_0_iibox_ce49),
    .q49(decipher_0_iibox_q49),
    .address50(decipher_0_iibox_address50),
    .ce50(decipher_0_iibox_ce50),
    .q50(decipher_0_iibox_q50),
    .address51(decipher_0_iibox_address51),
    .ce51(decipher_0_iibox_ce51),
    .q51(decipher_0_iibox_q51),
    .address52(decipher_0_iibox_address52),
    .ce52(decipher_0_iibox_ce52),
    .q52(decipher_0_iibox_q52),
    .address53(decipher_0_iibox_address53),
    .ce53(decipher_0_iibox_ce53),
    .q53(decipher_0_iibox_q53),
    .address54(decipher_0_iibox_address54),
    .ce54(decipher_0_iibox_ce54),
    .q54(decipher_0_iibox_q54),
    .address55(decipher_0_iibox_address55),
    .ce55(decipher_0_iibox_ce55),
    .q55(decipher_0_iibox_q55),
    .address56(decipher_0_iibox_address56),
    .ce56(decipher_0_iibox_ce56),
    .q56(decipher_0_iibox_q56),
    .address57(decipher_0_iibox_address57),
    .ce57(decipher_0_iibox_ce57),
    .q57(decipher_0_iibox_q57),
    .address58(decipher_0_iibox_address58),
    .ce58(decipher_0_iibox_ce58),
    .q58(decipher_0_iibox_q58),
    .address59(decipher_0_iibox_address59),
    .ce59(decipher_0_iibox_ce59),
    .q59(decipher_0_iibox_q59),
    .address60(decipher_0_iibox_address60),
    .ce60(decipher_0_iibox_ce60),
    .q60(decipher_0_iibox_q60),
    .address61(decipher_0_iibox_address61),
    .ce61(decipher_0_iibox_ce61),
    .q61(decipher_0_iibox_q61),
    .address62(decipher_0_iibox_address62),
    .ce62(decipher_0_iibox_ce62),
    .q62(decipher_0_iibox_q62),
    .address63(decipher_0_iibox_address63),
    .ce63(decipher_0_iibox_ce63),
    .q63(decipher_0_iibox_q63),
    .address64(decipher_0_iibox_address64),
    .ce64(decipher_0_iibox_ce64),
    .q64(decipher_0_iibox_q64),
    .address65(decipher_0_iibox_address65),
    .ce65(decipher_0_iibox_ce65),
    .q65(decipher_0_iibox_q65),
    .address66(decipher_0_iibox_address66),
    .ce66(decipher_0_iibox_ce66),
    .q66(decipher_0_iibox_q66),
    .address67(decipher_0_iibox_address67),
    .ce67(decipher_0_iibox_ce67),
    .q67(decipher_0_iibox_q67),
    .address68(decipher_0_iibox_address68),
    .ce68(decipher_0_iibox_ce68),
    .q68(decipher_0_iibox_q68),
    .address69(decipher_0_iibox_address69),
    .ce69(decipher_0_iibox_ce69),
    .q69(decipher_0_iibox_q69),
    .address70(decipher_0_iibox_address70),
    .ce70(decipher_0_iibox_ce70),
    .q70(decipher_0_iibox_q70),
    .address71(decipher_0_iibox_address71),
    .ce71(decipher_0_iibox_ce71),
    .q71(decipher_0_iibox_q71),
    .address72(decipher_0_iibox_address72),
    .ce72(decipher_0_iibox_ce72),
    .q72(decipher_0_iibox_q72),
    .address73(decipher_0_iibox_address73),
    .ce73(decipher_0_iibox_ce73),
    .q73(decipher_0_iibox_q73),
    .address74(decipher_0_iibox_address74),
    .ce74(decipher_0_iibox_ce74),
    .q74(decipher_0_iibox_q74),
    .address75(decipher_0_iibox_address75),
    .ce75(decipher_0_iibox_ce75),
    .q75(decipher_0_iibox_q75),
    .address76(decipher_0_iibox_address76),
    .ce76(decipher_0_iibox_ce76),
    .q76(decipher_0_iibox_q76),
    .address77(decipher_0_iibox_address77),
    .ce77(decipher_0_iibox_ce77),
    .q77(decipher_0_iibox_q77),
    .address78(decipher_0_iibox_address78),
    .ce78(decipher_0_iibox_ce78),
    .q78(decipher_0_iibox_q78),
    .address79(decipher_0_iibox_address79),
    .ce79(decipher_0_iibox_ce79),
    .q79(decipher_0_iibox_q79),
    .address80(decipher_0_iibox_address80),
    .ce80(decipher_0_iibox_ce80),
    .q80(decipher_0_iibox_q80),
    .address81(decipher_0_iibox_address81),
    .ce81(decipher_0_iibox_ce81),
    .q81(decipher_0_iibox_q81),
    .address82(decipher_0_iibox_address82),
    .ce82(decipher_0_iibox_ce82),
    .q82(decipher_0_iibox_q82),
    .address83(decipher_0_iibox_address83),
    .ce83(decipher_0_iibox_ce83),
    .q83(decipher_0_iibox_q83),
    .address84(decipher_0_iibox_address84),
    .ce84(decipher_0_iibox_ce84),
    .q84(decipher_0_iibox_q84),
    .address85(decipher_0_iibox_address85),
    .ce85(decipher_0_iibox_ce85),
    .q85(decipher_0_iibox_q85),
    .address86(decipher_0_iibox_address86),
    .ce86(decipher_0_iibox_ce86),
    .q86(decipher_0_iibox_q86),
    .address87(decipher_0_iibox_address87),
    .ce87(decipher_0_iibox_ce87),
    .q87(decipher_0_iibox_q87),
    .address88(decipher_0_iibox_address88),
    .ce88(decipher_0_iibox_ce88),
    .q88(decipher_0_iibox_q88),
    .address89(decipher_0_iibox_address89),
    .ce89(decipher_0_iibox_ce89),
    .q89(decipher_0_iibox_q89),
    .address90(decipher_0_iibox_address90),
    .ce90(decipher_0_iibox_ce90),
    .q90(decipher_0_iibox_q90),
    .address91(decipher_0_iibox_address91),
    .ce91(decipher_0_iibox_ce91),
    .q91(decipher_0_iibox_q91),
    .address92(decipher_0_iibox_address92),
    .ce92(decipher_0_iibox_ce92),
    .q92(decipher_0_iibox_q92),
    .address93(decipher_0_iibox_address93),
    .ce93(decipher_0_iibox_ce93),
    .q93(decipher_0_iibox_q93),
    .address94(decipher_0_iibox_address94),
    .ce94(decipher_0_iibox_ce94),
    .q94(decipher_0_iibox_q94),
    .address95(decipher_0_iibox_address95),
    .ce95(decipher_0_iibox_ce95),
    .q95(decipher_0_iibox_q95),
    .address96(decipher_0_iibox_address96),
    .ce96(decipher_0_iibox_ce96),
    .q96(decipher_0_iibox_q96),
    .address97(decipher_0_iibox_address97),
    .ce97(decipher_0_iibox_ce97),
    .q97(decipher_0_iibox_q97),
    .address98(decipher_0_iibox_address98),
    .ce98(decipher_0_iibox_ce98),
    .q98(decipher_0_iibox_q98),
    .address99(decipher_0_iibox_address99),
    .ce99(decipher_0_iibox_ce99),
    .q99(decipher_0_iibox_q99),
    .address100(decipher_0_iibox_address100),
    .ce100(decipher_0_iibox_ce100),
    .q100(decipher_0_iibox_q100),
    .address101(decipher_0_iibox_address101),
    .ce101(decipher_0_iibox_ce101),
    .q101(decipher_0_iibox_q101),
    .address102(decipher_0_iibox_address102),
    .ce102(decipher_0_iibox_ce102),
    .q102(decipher_0_iibox_q102),
    .address103(decipher_0_iibox_address103),
    .ce103(decipher_0_iibox_ce103),
    .q103(decipher_0_iibox_q103),
    .address104(decipher_0_iibox_address104),
    .ce104(decipher_0_iibox_ce104),
    .q104(decipher_0_iibox_q104),
    .address105(decipher_0_iibox_address105),
    .ce105(decipher_0_iibox_ce105),
    .q105(decipher_0_iibox_q105),
    .address106(decipher_0_iibox_address106),
    .ce106(decipher_0_iibox_ce106),
    .q106(decipher_0_iibox_q106),
    .address107(decipher_0_iibox_address107),
    .ce107(decipher_0_iibox_ce107),
    .q107(decipher_0_iibox_q107),
    .address108(decipher_0_iibox_address108),
    .ce108(decipher_0_iibox_ce108),
    .q108(decipher_0_iibox_q108),
    .address109(decipher_0_iibox_address109),
    .ce109(decipher_0_iibox_ce109),
    .q109(decipher_0_iibox_q109),
    .address110(decipher_0_iibox_address110),
    .ce110(decipher_0_iibox_ce110),
    .q110(decipher_0_iibox_q110),
    .address111(decipher_0_iibox_address111),
    .ce111(decipher_0_iibox_ce111),
    .q111(decipher_0_iibox_q111),
    .address112(decipher_0_iibox_address112),
    .ce112(decipher_0_iibox_ce112),
    .q112(decipher_0_iibox_q112),
    .address113(decipher_0_iibox_address113),
    .ce113(decipher_0_iibox_ce113),
    .q113(decipher_0_iibox_q113),
    .address114(decipher_0_iibox_address114),
    .ce114(decipher_0_iibox_ce114),
    .q114(decipher_0_iibox_q114),
    .address115(decipher_0_iibox_address115),
    .ce115(decipher_0_iibox_ce115),
    .q115(decipher_0_iibox_q115),
    .address116(decipher_0_iibox_address116),
    .ce116(decipher_0_iibox_ce116),
    .q116(decipher_0_iibox_q116),
    .address117(decipher_0_iibox_address117),
    .ce117(decipher_0_iibox_ce117),
    .q117(decipher_0_iibox_q117),
    .address118(decipher_0_iibox_address118),
    .ce118(decipher_0_iibox_ce118),
    .q118(decipher_0_iibox_q118),
    .address119(decipher_0_iibox_address119),
    .ce119(decipher_0_iibox_ce119),
    .q119(decipher_0_iibox_q119),
    .address120(decipher_0_iibox_address120),
    .ce120(decipher_0_iibox_ce120),
    .q120(decipher_0_iibox_q120),
    .address121(decipher_0_iibox_address121),
    .ce121(decipher_0_iibox_ce121),
    .q121(decipher_0_iibox_q121),
    .address122(decipher_0_iibox_address122),
    .ce122(decipher_0_iibox_ce122),
    .q122(decipher_0_iibox_q122),
    .address123(decipher_0_iibox_address123),
    .ce123(decipher_0_iibox_ce123),
    .q123(decipher_0_iibox_q123),
    .address124(decipher_0_iibox_address124),
    .ce124(decipher_0_iibox_ce124),
    .q124(decipher_0_iibox_q124),
    .address125(decipher_0_iibox_address125),
    .ce125(decipher_0_iibox_ce125),
    .q125(decipher_0_iibox_q125),
    .address126(decipher_0_iibox_address126),
    .ce126(decipher_0_iibox_ce126),
    .q126(decipher_0_iibox_q126),
    .address127(decipher_0_iibox_address127),
    .ce127(decipher_0_iibox_ce127),
    .q127(decipher_0_iibox_q127),
    .address128(decipher_0_iibox_address128),
    .ce128(decipher_0_iibox_ce128),
    .q128(decipher_0_iibox_q128),
    .address129(decipher_0_iibox_address129),
    .ce129(decipher_0_iibox_ce129),
    .q129(decipher_0_iibox_q129),
    .address130(decipher_0_iibox_address130),
    .ce130(decipher_0_iibox_ce130),
    .q130(decipher_0_iibox_q130),
    .address131(decipher_0_iibox_address131),
    .ce131(decipher_0_iibox_ce131),
    .q131(decipher_0_iibox_q131),
    .address132(decipher_0_iibox_address132),
    .ce132(decipher_0_iibox_ce132),
    .q132(decipher_0_iibox_q132),
    .address133(decipher_0_iibox_address133),
    .ce133(decipher_0_iibox_ce133),
    .q133(decipher_0_iibox_q133),
    .address134(decipher_0_iibox_address134),
    .ce134(decipher_0_iibox_ce134),
    .q134(decipher_0_iibox_q134),
    .address135(decipher_0_iibox_address135),
    .ce135(decipher_0_iibox_ce135),
    .q135(decipher_0_iibox_q135),
    .address136(decipher_0_iibox_address136),
    .ce136(decipher_0_iibox_ce136),
    .q136(decipher_0_iibox_q136),
    .address137(decipher_0_iibox_address137),
    .ce137(decipher_0_iibox_ce137),
    .q137(decipher_0_iibox_q137),
    .address138(decipher_0_iibox_address138),
    .ce138(decipher_0_iibox_ce138),
    .q138(decipher_0_iibox_q138),
    .address139(decipher_0_iibox_address139),
    .ce139(decipher_0_iibox_ce139),
    .q139(decipher_0_iibox_q139),
    .address140(decipher_0_iibox_address140),
    .ce140(decipher_0_iibox_ce140),
    .q140(decipher_0_iibox_q140),
    .address141(decipher_0_iibox_address141),
    .ce141(decipher_0_iibox_ce141),
    .q141(decipher_0_iibox_q141),
    .address142(decipher_0_iibox_address142),
    .ce142(decipher_0_iibox_ce142),
    .q142(decipher_0_iibox_q142),
    .address143(decipher_0_iibox_address143),
    .ce143(decipher_0_iibox_ce143),
    .q143(decipher_0_iibox_q143),
    .address144(decipher_0_iibox_address144),
    .ce144(decipher_0_iibox_ce144),
    .q144(decipher_0_iibox_q144),
    .address145(decipher_0_iibox_address145),
    .ce145(decipher_0_iibox_ce145),
    .q145(decipher_0_iibox_q145),
    .address146(decipher_0_iibox_address146),
    .ce146(decipher_0_iibox_ce146),
    .q146(decipher_0_iibox_q146),
    .address147(decipher_0_iibox_address147),
    .ce147(decipher_0_iibox_ce147),
    .q147(decipher_0_iibox_q147),
    .address148(decipher_0_iibox_address148),
    .ce148(decipher_0_iibox_ce148),
    .q148(decipher_0_iibox_q148),
    .address149(decipher_0_iibox_address149),
    .ce149(decipher_0_iibox_ce149),
    .q149(decipher_0_iibox_q149),
    .address150(decipher_0_iibox_address150),
    .ce150(decipher_0_iibox_ce150),
    .q150(decipher_0_iibox_q150),
    .address151(decipher_0_iibox_address151),
    .ce151(decipher_0_iibox_ce151),
    .q151(decipher_0_iibox_q151),
    .address152(decipher_0_iibox_address152),
    .ce152(decipher_0_iibox_ce152),
    .q152(decipher_0_iibox_q152),
    .address153(decipher_0_iibox_address153),
    .ce153(decipher_0_iibox_ce153),
    .q153(decipher_0_iibox_q153),
    .address154(decipher_0_iibox_address154),
    .ce154(decipher_0_iibox_ce154),
    .q154(decipher_0_iibox_q154),
    .address155(decipher_0_iibox_address155),
    .ce155(decipher_0_iibox_ce155),
    .q155(decipher_0_iibox_q155),
    .address156(decipher_0_iibox_address156),
    .ce156(decipher_0_iibox_ce156),
    .q156(decipher_0_iibox_q156),
    .address157(decipher_0_iibox_address157),
    .ce157(decipher_0_iibox_ce157),
    .q157(decipher_0_iibox_q157),
    .address158(decipher_0_iibox_address158),
    .ce158(decipher_0_iibox_ce158),
    .q158(decipher_0_iibox_q158),
    .address159(decipher_0_iibox_address159),
    .ce159(decipher_0_iibox_ce159),
    .q159(decipher_0_iibox_q159)
);

testDec_process_r_decipher_0_i32box_ROM_NP_LUTRAM_1R #(
    .DataWidth( 32 ),
    .AddressRange( 256 ),
    .AddressWidth( 8 ))
decipher_0_i32box_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(decipher_0_i32box_address0),
    .ce0(decipher_0_i32box_ce0),
    .q0(decipher_0_i32box_q0),
    .address1(decipher_0_i32box_address1),
    .ce1(decipher_0_i32box_ce1),
    .q1(decipher_0_i32box_q1),
    .address2(decipher_0_i32box_address2),
    .ce2(decipher_0_i32box_ce2),
    .q2(decipher_0_i32box_q2),
    .address3(decipher_0_i32box_address3),
    .ce3(decipher_0_i32box_ce3),
    .q3(decipher_0_i32box_q3),
    .address4(decipher_0_i32box_address4),
    .ce4(decipher_0_i32box_ce4),
    .q4(decipher_0_i32box_q4),
    .address5(decipher_0_i32box_address5),
    .ce5(decipher_0_i32box_ce5),
    .q5(decipher_0_i32box_q5),
    .address6(decipher_0_i32box_address6),
    .ce6(decipher_0_i32box_ce6),
    .q6(decipher_0_i32box_q6),
    .address7(decipher_0_i32box_address7),
    .ce7(decipher_0_i32box_ce7),
    .q7(decipher_0_i32box_q7),
    .address8(decipher_0_i32box_address8),
    .ce8(decipher_0_i32box_ce8),
    .q8(decipher_0_i32box_q8),
    .address9(decipher_0_i32box_address9),
    .ce9(decipher_0_i32box_ce9),
    .q9(decipher_0_i32box_q9),
    .address10(decipher_0_i32box_address10),
    .ce10(decipher_0_i32box_ce10),
    .q10(decipher_0_i32box_q10),
    .address11(decipher_0_i32box_address11),
    .ce11(decipher_0_i32box_ce11),
    .q11(decipher_0_i32box_q11),
    .address12(decipher_0_i32box_address12),
    .ce12(decipher_0_i32box_ce12),
    .q12(decipher_0_i32box_q12),
    .address13(decipher_0_i32box_address13),
    .ce13(decipher_0_i32box_ce13),
    .q13(decipher_0_i32box_q13),
    .address14(decipher_0_i32box_address14),
    .ce14(decipher_0_i32box_ce14),
    .q14(decipher_0_i32box_q14),
    .address15(decipher_0_i32box_address15),
    .ce15(decipher_0_i32box_ce15),
    .q15(decipher_0_i32box_q15),
    .address16(decipher_0_i32box_address16),
    .ce16(decipher_0_i32box_ce16),
    .q16(decipher_0_i32box_q16),
    .address17(decipher_0_i32box_address17),
    .ce17(decipher_0_i32box_ce17),
    .q17(decipher_0_i32box_q17),
    .address18(decipher_0_i32box_address18),
    .ce18(decipher_0_i32box_ce18),
    .q18(decipher_0_i32box_q18),
    .address19(decipher_0_i32box_address19),
    .ce19(decipher_0_i32box_ce19),
    .q19(decipher_0_i32box_q19),
    .address20(decipher_0_i32box_address20),
    .ce20(decipher_0_i32box_ce20),
    .q20(decipher_0_i32box_q20),
    .address21(decipher_0_i32box_address21),
    .ce21(decipher_0_i32box_ce21),
    .q21(decipher_0_i32box_q21),
    .address22(decipher_0_i32box_address22),
    .ce22(decipher_0_i32box_ce22),
    .q22(decipher_0_i32box_q22),
    .address23(decipher_0_i32box_address23),
    .ce23(decipher_0_i32box_ce23),
    .q23(decipher_0_i32box_q23),
    .address24(decipher_0_i32box_address24),
    .ce24(decipher_0_i32box_ce24),
    .q24(decipher_0_i32box_q24),
    .address25(decipher_0_i32box_address25),
    .ce25(decipher_0_i32box_ce25),
    .q25(decipher_0_i32box_q25),
    .address26(decipher_0_i32box_address26),
    .ce26(decipher_0_i32box_ce26),
    .q26(decipher_0_i32box_q26),
    .address27(decipher_0_i32box_address27),
    .ce27(decipher_0_i32box_ce27),
    .q27(decipher_0_i32box_q27),
    .address28(decipher_0_i32box_address28),
    .ce28(decipher_0_i32box_ce28),
    .q28(decipher_0_i32box_q28),
    .address29(decipher_0_i32box_address29),
    .ce29(decipher_0_i32box_ce29),
    .q29(decipher_0_i32box_q29),
    .address30(decipher_0_i32box_address30),
    .ce30(decipher_0_i32box_ce30),
    .q30(decipher_0_i32box_q30),
    .address31(decipher_0_i32box_address31),
    .ce31(decipher_0_i32box_ce31),
    .q31(decipher_0_i32box_q31),
    .address32(decipher_0_i32box_address32),
    .ce32(decipher_0_i32box_ce32),
    .q32(decipher_0_i32box_q32),
    .address33(decipher_0_i32box_address33),
    .ce33(decipher_0_i32box_ce33),
    .q33(decipher_0_i32box_q33),
    .address34(decipher_0_i32box_address34),
    .ce34(decipher_0_i32box_ce34),
    .q34(decipher_0_i32box_q34),
    .address35(decipher_0_i32box_address35),
    .ce35(decipher_0_i32box_ce35),
    .q35(decipher_0_i32box_q35),
    .address36(decipher_0_i32box_address36),
    .ce36(decipher_0_i32box_ce36),
    .q36(decipher_0_i32box_q36),
    .address37(decipher_0_i32box_address37),
    .ce37(decipher_0_i32box_ce37),
    .q37(decipher_0_i32box_q37),
    .address38(decipher_0_i32box_address38),
    .ce38(decipher_0_i32box_ce38),
    .q38(decipher_0_i32box_q38),
    .address39(decipher_0_i32box_address39),
    .ce39(decipher_0_i32box_ce39),
    .q39(decipher_0_i32box_q39),
    .address40(decipher_0_i32box_address40),
    .ce40(decipher_0_i32box_ce40),
    .q40(decipher_0_i32box_q40),
    .address41(decipher_0_i32box_address41),
    .ce41(decipher_0_i32box_ce41),
    .q41(decipher_0_i32box_q41),
    .address42(decipher_0_i32box_address42),
    .ce42(decipher_0_i32box_ce42),
    .q42(decipher_0_i32box_q42),
    .address43(decipher_0_i32box_address43),
    .ce43(decipher_0_i32box_ce43),
    .q43(decipher_0_i32box_q43),
    .address44(decipher_0_i32box_address44),
    .ce44(decipher_0_i32box_ce44),
    .q44(decipher_0_i32box_q44),
    .address45(decipher_0_i32box_address45),
    .ce45(decipher_0_i32box_ce45),
    .q45(decipher_0_i32box_q45),
    .address46(decipher_0_i32box_address46),
    .ce46(decipher_0_i32box_ce46),
    .q46(decipher_0_i32box_q46),
    .address47(decipher_0_i32box_address47),
    .ce47(decipher_0_i32box_ce47),
    .q47(decipher_0_i32box_q47),
    .address48(decipher_0_i32box_address48),
    .ce48(decipher_0_i32box_ce48),
    .q48(decipher_0_i32box_q48),
    .address49(decipher_0_i32box_address49),
    .ce49(decipher_0_i32box_ce49),
    .q49(decipher_0_i32box_q49),
    .address50(decipher_0_i32box_address50),
    .ce50(decipher_0_i32box_ce50),
    .q50(decipher_0_i32box_q50),
    .address51(decipher_0_i32box_address51),
    .ce51(decipher_0_i32box_ce51),
    .q51(decipher_0_i32box_q51),
    .address52(decipher_0_i32box_address52),
    .ce52(decipher_0_i32box_ce52),
    .q52(decipher_0_i32box_q52),
    .address53(decipher_0_i32box_address53),
    .ce53(decipher_0_i32box_ce53),
    .q53(decipher_0_i32box_q53),
    .address54(decipher_0_i32box_address54),
    .ce54(decipher_0_i32box_ce54),
    .q54(decipher_0_i32box_q54),
    .address55(decipher_0_i32box_address55),
    .ce55(decipher_0_i32box_ce55),
    .q55(decipher_0_i32box_q55),
    .address56(decipher_0_i32box_address56),
    .ce56(decipher_0_i32box_ce56),
    .q56(decipher_0_i32box_q56),
    .address57(decipher_0_i32box_address57),
    .ce57(decipher_0_i32box_ce57),
    .q57(decipher_0_i32box_q57),
    .address58(decipher_0_i32box_address58),
    .ce58(decipher_0_i32box_ce58),
    .q58(decipher_0_i32box_q58),
    .address59(decipher_0_i32box_address59),
    .ce59(decipher_0_i32box_ce59),
    .q59(decipher_0_i32box_q59),
    .address60(decipher_0_i32box_address60),
    .ce60(decipher_0_i32box_ce60),
    .q60(decipher_0_i32box_q60),
    .address61(decipher_0_i32box_address61),
    .ce61(decipher_0_i32box_ce61),
    .q61(decipher_0_i32box_q61),
    .address62(decipher_0_i32box_address62),
    .ce62(decipher_0_i32box_ce62),
    .q62(decipher_0_i32box_q62),
    .address63(decipher_0_i32box_address63),
    .ce63(decipher_0_i32box_ce63),
    .q63(decipher_0_i32box_q63),
    .address64(decipher_0_i32box_address64),
    .ce64(decipher_0_i32box_ce64),
    .q64(decipher_0_i32box_q64),
    .address65(decipher_0_i32box_address65),
    .ce65(decipher_0_i32box_ce65),
    .q65(decipher_0_i32box_q65),
    .address66(decipher_0_i32box_address66),
    .ce66(decipher_0_i32box_ce66),
    .q66(decipher_0_i32box_q66),
    .address67(decipher_0_i32box_address67),
    .ce67(decipher_0_i32box_ce67),
    .q67(decipher_0_i32box_q67),
    .address68(decipher_0_i32box_address68),
    .ce68(decipher_0_i32box_ce68),
    .q68(decipher_0_i32box_q68),
    .address69(decipher_0_i32box_address69),
    .ce69(decipher_0_i32box_ce69),
    .q69(decipher_0_i32box_q69),
    .address70(decipher_0_i32box_address70),
    .ce70(decipher_0_i32box_ce70),
    .q70(decipher_0_i32box_q70),
    .address71(decipher_0_i32box_address71),
    .ce71(decipher_0_i32box_ce71),
    .q71(decipher_0_i32box_q71),
    .address72(decipher_0_i32box_address72),
    .ce72(decipher_0_i32box_ce72),
    .q72(decipher_0_i32box_q72),
    .address73(decipher_0_i32box_address73),
    .ce73(decipher_0_i32box_ce73),
    .q73(decipher_0_i32box_q73),
    .address74(decipher_0_i32box_address74),
    .ce74(decipher_0_i32box_ce74),
    .q74(decipher_0_i32box_q74),
    .address75(decipher_0_i32box_address75),
    .ce75(decipher_0_i32box_ce75),
    .q75(decipher_0_i32box_q75),
    .address76(decipher_0_i32box_address76),
    .ce76(decipher_0_i32box_ce76),
    .q76(decipher_0_i32box_q76),
    .address77(decipher_0_i32box_address77),
    .ce77(decipher_0_i32box_ce77),
    .q77(decipher_0_i32box_q77),
    .address78(decipher_0_i32box_address78),
    .ce78(decipher_0_i32box_ce78),
    .q78(decipher_0_i32box_q78),
    .address79(decipher_0_i32box_address79),
    .ce79(decipher_0_i32box_ce79),
    .q79(decipher_0_i32box_q79),
    .address80(decipher_0_i32box_address80),
    .ce80(decipher_0_i32box_ce80),
    .q80(decipher_0_i32box_q80),
    .address81(decipher_0_i32box_address81),
    .ce81(decipher_0_i32box_ce81),
    .q81(decipher_0_i32box_q81),
    .address82(decipher_0_i32box_address82),
    .ce82(decipher_0_i32box_ce82),
    .q82(decipher_0_i32box_q82),
    .address83(decipher_0_i32box_address83),
    .ce83(decipher_0_i32box_ce83),
    .q83(decipher_0_i32box_q83),
    .address84(decipher_0_i32box_address84),
    .ce84(decipher_0_i32box_ce84),
    .q84(decipher_0_i32box_q84),
    .address85(decipher_0_i32box_address85),
    .ce85(decipher_0_i32box_ce85),
    .q85(decipher_0_i32box_q85),
    .address86(decipher_0_i32box_address86),
    .ce86(decipher_0_i32box_ce86),
    .q86(decipher_0_i32box_q86),
    .address87(decipher_0_i32box_address87),
    .ce87(decipher_0_i32box_ce87),
    .q87(decipher_0_i32box_q87),
    .address88(decipher_0_i32box_address88),
    .ce88(decipher_0_i32box_ce88),
    .q88(decipher_0_i32box_q88),
    .address89(decipher_0_i32box_address89),
    .ce89(decipher_0_i32box_ce89),
    .q89(decipher_0_i32box_q89),
    .address90(decipher_0_i32box_address90),
    .ce90(decipher_0_i32box_ce90),
    .q90(decipher_0_i32box_q90),
    .address91(decipher_0_i32box_address91),
    .ce91(decipher_0_i32box_ce91),
    .q91(decipher_0_i32box_q91),
    .address92(decipher_0_i32box_address92),
    .ce92(decipher_0_i32box_ce92),
    .q92(decipher_0_i32box_q92),
    .address93(decipher_0_i32box_address93),
    .ce93(decipher_0_i32box_ce93),
    .q93(decipher_0_i32box_q93),
    .address94(decipher_0_i32box_address94),
    .ce94(decipher_0_i32box_ce94),
    .q94(decipher_0_i32box_q94),
    .address95(decipher_0_i32box_address95),
    .ce95(decipher_0_i32box_ce95),
    .q95(decipher_0_i32box_q95),
    .address96(decipher_0_i32box_address96),
    .ce96(decipher_0_i32box_ce96),
    .q96(decipher_0_i32box_q96),
    .address97(decipher_0_i32box_address97),
    .ce97(decipher_0_i32box_ce97),
    .q97(decipher_0_i32box_q97),
    .address98(decipher_0_i32box_address98),
    .ce98(decipher_0_i32box_ce98),
    .q98(decipher_0_i32box_q98),
    .address99(decipher_0_i32box_address99),
    .ce99(decipher_0_i32box_ce99),
    .q99(decipher_0_i32box_q99),
    .address100(decipher_0_i32box_address100),
    .ce100(decipher_0_i32box_ce100),
    .q100(decipher_0_i32box_q100),
    .address101(decipher_0_i32box_address101),
    .ce101(decipher_0_i32box_ce101),
    .q101(decipher_0_i32box_q101),
    .address102(decipher_0_i32box_address102),
    .ce102(decipher_0_i32box_ce102),
    .q102(decipher_0_i32box_q102),
    .address103(decipher_0_i32box_address103),
    .ce103(decipher_0_i32box_ce103),
    .q103(decipher_0_i32box_q103),
    .address104(decipher_0_i32box_address104),
    .ce104(decipher_0_i32box_ce104),
    .q104(decipher_0_i32box_q104),
    .address105(decipher_0_i32box_address105),
    .ce105(decipher_0_i32box_ce105),
    .q105(decipher_0_i32box_q105),
    .address106(decipher_0_i32box_address106),
    .ce106(decipher_0_i32box_ce106),
    .q106(decipher_0_i32box_q106),
    .address107(decipher_0_i32box_address107),
    .ce107(decipher_0_i32box_ce107),
    .q107(decipher_0_i32box_q107),
    .address108(decipher_0_i32box_address108),
    .ce108(decipher_0_i32box_ce108),
    .q108(decipher_0_i32box_q108),
    .address109(decipher_0_i32box_address109),
    .ce109(decipher_0_i32box_ce109),
    .q109(decipher_0_i32box_q109),
    .address110(decipher_0_i32box_address110),
    .ce110(decipher_0_i32box_ce110),
    .q110(decipher_0_i32box_q110),
    .address111(decipher_0_i32box_address111),
    .ce111(decipher_0_i32box_ce111),
    .q111(decipher_0_i32box_q111),
    .address112(decipher_0_i32box_address112),
    .ce112(decipher_0_i32box_ce112),
    .q112(decipher_0_i32box_q112),
    .address113(decipher_0_i32box_address113),
    .ce113(decipher_0_i32box_ce113),
    .q113(decipher_0_i32box_q113),
    .address114(decipher_0_i32box_address114),
    .ce114(decipher_0_i32box_ce114),
    .q114(decipher_0_i32box_q114),
    .address115(decipher_0_i32box_address115),
    .ce115(decipher_0_i32box_ce115),
    .q115(decipher_0_i32box_q115),
    .address116(decipher_0_i32box_address116),
    .ce116(decipher_0_i32box_ce116),
    .q116(decipher_0_i32box_q116),
    .address117(decipher_0_i32box_address117),
    .ce117(decipher_0_i32box_ce117),
    .q117(decipher_0_i32box_q117),
    .address118(decipher_0_i32box_address118),
    .ce118(decipher_0_i32box_ce118),
    .q118(decipher_0_i32box_q118),
    .address119(decipher_0_i32box_address119),
    .ce119(decipher_0_i32box_ce119),
    .q119(decipher_0_i32box_q119),
    .address120(decipher_0_i32box_address120),
    .ce120(decipher_0_i32box_ce120),
    .q120(decipher_0_i32box_q120),
    .address121(decipher_0_i32box_address121),
    .ce121(decipher_0_i32box_ce121),
    .q121(decipher_0_i32box_q121),
    .address122(decipher_0_i32box_address122),
    .ce122(decipher_0_i32box_ce122),
    .q122(decipher_0_i32box_q122),
    .address123(decipher_0_i32box_address123),
    .ce123(decipher_0_i32box_ce123),
    .q123(decipher_0_i32box_q123),
    .address124(decipher_0_i32box_address124),
    .ce124(decipher_0_i32box_ce124),
    .q124(decipher_0_i32box_q124),
    .address125(decipher_0_i32box_address125),
    .ce125(decipher_0_i32box_ce125),
    .q125(decipher_0_i32box_q125),
    .address126(decipher_0_i32box_address126),
    .ce126(decipher_0_i32box_ce126),
    .q126(decipher_0_i32box_q126),
    .address127(decipher_0_i32box_address127),
    .ce127(decipher_0_i32box_ce127),
    .q127(decipher_0_i32box_q127),
    .address128(decipher_0_i32box_address128),
    .ce128(decipher_0_i32box_ce128),
    .q128(decipher_0_i32box_q128),
    .address129(decipher_0_i32box_address129),
    .ce129(decipher_0_i32box_ce129),
    .q129(decipher_0_i32box_q129),
    .address130(decipher_0_i32box_address130),
    .ce130(decipher_0_i32box_ce130),
    .q130(decipher_0_i32box_q130),
    .address131(decipher_0_i32box_address131),
    .ce131(decipher_0_i32box_ce131),
    .q131(decipher_0_i32box_q131),
    .address132(decipher_0_i32box_address132),
    .ce132(decipher_0_i32box_ce132),
    .q132(decipher_0_i32box_q132),
    .address133(decipher_0_i32box_address133),
    .ce133(decipher_0_i32box_ce133),
    .q133(decipher_0_i32box_q133),
    .address134(decipher_0_i32box_address134),
    .ce134(decipher_0_i32box_ce134),
    .q134(decipher_0_i32box_q134),
    .address135(decipher_0_i32box_address135),
    .ce135(decipher_0_i32box_ce135),
    .q135(decipher_0_i32box_q135),
    .address136(decipher_0_i32box_address136),
    .ce136(decipher_0_i32box_ce136),
    .q136(decipher_0_i32box_q136),
    .address137(decipher_0_i32box_address137),
    .ce137(decipher_0_i32box_ce137),
    .q137(decipher_0_i32box_q137),
    .address138(decipher_0_i32box_address138),
    .ce138(decipher_0_i32box_ce138),
    .q138(decipher_0_i32box_q138),
    .address139(decipher_0_i32box_address139),
    .ce139(decipher_0_i32box_ce139),
    .q139(decipher_0_i32box_q139),
    .address140(decipher_0_i32box_address140),
    .ce140(decipher_0_i32box_ce140),
    .q140(decipher_0_i32box_q140),
    .address141(decipher_0_i32box_address141),
    .ce141(decipher_0_i32box_ce141),
    .q141(decipher_0_i32box_q141),
    .address142(decipher_0_i32box_address142),
    .ce142(decipher_0_i32box_ce142),
    .q142(decipher_0_i32box_q142),
    .address143(decipher_0_i32box_address143),
    .ce143(decipher_0_i32box_ce143),
    .q143(decipher_0_i32box_q143)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_enable_reg_pp0_iter1 <= ap_start;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter10 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter10 <= ap_enable_reg_pp0_iter9;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter11 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter11 <= ap_enable_reg_pp0_iter10;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter12 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter12 <= ap_enable_reg_pp0_iter11;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter13 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter13 <= ap_enable_reg_pp0_iter12;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter14 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter14 <= ap_enable_reg_pp0_iter13;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter15 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter15 <= ap_enable_reg_pp0_iter14;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter16 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter16 <= ap_enable_reg_pp0_iter15;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter17 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter17 <= ap_enable_reg_pp0_iter16;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter18 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter18 <= ap_enable_reg_pp0_iter17;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter19 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter19 <= ap_enable_reg_pp0_iter18;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter5 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter6 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter7 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter8 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter8 <= ap_enable_reg_pp0_iter7;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter9 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter9 <= ap_enable_reg_pp0_iter8;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        p_read11_reg_14837 <= p_read;
        p_read11_reg_14837_pp0_iter1_reg <= p_read11_reg_14837;
        p_read_10_reg_14832 <= p_read1;
        p_read_10_reg_14832_pp0_iter1_reg <= p_read_10_reg_14832;
        p_read_2_reg_14792 <= p_read9;
        p_read_3_reg_14797 <= p_read8;
        p_read_3_reg_14797_pp0_iter1_reg <= p_read_3_reg_14797;
        p_read_4_reg_14802 <= p_read7;
        p_read_4_reg_14802_pp0_iter1_reg <= p_read_4_reg_14802;
        p_read_5_reg_14807 <= p_read6;
        p_read_5_reg_14807_pp0_iter1_reg <= p_read_5_reg_14807;
        p_read_6_reg_14812 <= p_read5;
        p_read_6_reg_14812_pp0_iter1_reg <= p_read_6_reg_14812;
        p_read_7_reg_14817 <= p_read4;
        p_read_7_reg_14817_pp0_iter1_reg <= p_read_7_reg_14817;
        p_read_8_reg_14822 <= p_read3;
        p_read_8_reg_14822_pp0_iter1_reg <= p_read_8_reg_14822;
        p_read_9_reg_14827 <= p_read2;
        p_read_9_reg_14827_pp0_iter1_reg <= p_read_9_reg_14827;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        p_read11_reg_14837_pp0_iter10_reg <= p_read11_reg_14837_pp0_iter9_reg;
        p_read11_reg_14837_pp0_iter11_reg <= p_read11_reg_14837_pp0_iter10_reg;
        p_read11_reg_14837_pp0_iter12_reg <= p_read11_reg_14837_pp0_iter11_reg;
        p_read11_reg_14837_pp0_iter13_reg <= p_read11_reg_14837_pp0_iter12_reg;
        p_read11_reg_14837_pp0_iter14_reg <= p_read11_reg_14837_pp0_iter13_reg;
        p_read11_reg_14837_pp0_iter15_reg <= p_read11_reg_14837_pp0_iter14_reg;
        p_read11_reg_14837_pp0_iter16_reg <= p_read11_reg_14837_pp0_iter15_reg;
        p_read11_reg_14837_pp0_iter17_reg <= p_read11_reg_14837_pp0_iter16_reg;
        p_read11_reg_14837_pp0_iter18_reg <= p_read11_reg_14837_pp0_iter17_reg;
        p_read11_reg_14837_pp0_iter2_reg <= p_read11_reg_14837_pp0_iter1_reg;
        p_read11_reg_14837_pp0_iter3_reg <= p_read11_reg_14837_pp0_iter2_reg;
        p_read11_reg_14837_pp0_iter4_reg <= p_read11_reg_14837_pp0_iter3_reg;
        p_read11_reg_14837_pp0_iter5_reg <= p_read11_reg_14837_pp0_iter4_reg;
        p_read11_reg_14837_pp0_iter6_reg <= p_read11_reg_14837_pp0_iter5_reg;
        p_read11_reg_14837_pp0_iter7_reg <= p_read11_reg_14837_pp0_iter6_reg;
        p_read11_reg_14837_pp0_iter8_reg <= p_read11_reg_14837_pp0_iter7_reg;
        p_read11_reg_14837_pp0_iter9_reg <= p_read11_reg_14837_pp0_iter8_reg;
        p_read_10_reg_14832_pp0_iter10_reg <= p_read_10_reg_14832_pp0_iter9_reg;
        p_read_10_reg_14832_pp0_iter11_reg <= p_read_10_reg_14832_pp0_iter10_reg;
        p_read_10_reg_14832_pp0_iter12_reg <= p_read_10_reg_14832_pp0_iter11_reg;
        p_read_10_reg_14832_pp0_iter13_reg <= p_read_10_reg_14832_pp0_iter12_reg;
        p_read_10_reg_14832_pp0_iter14_reg <= p_read_10_reg_14832_pp0_iter13_reg;
        p_read_10_reg_14832_pp0_iter15_reg <= p_read_10_reg_14832_pp0_iter14_reg;
        p_read_10_reg_14832_pp0_iter16_reg <= p_read_10_reg_14832_pp0_iter15_reg;
        p_read_10_reg_14832_pp0_iter2_reg <= p_read_10_reg_14832_pp0_iter1_reg;
        p_read_10_reg_14832_pp0_iter3_reg <= p_read_10_reg_14832_pp0_iter2_reg;
        p_read_10_reg_14832_pp0_iter4_reg <= p_read_10_reg_14832_pp0_iter3_reg;
        p_read_10_reg_14832_pp0_iter5_reg <= p_read_10_reg_14832_pp0_iter4_reg;
        p_read_10_reg_14832_pp0_iter6_reg <= p_read_10_reg_14832_pp0_iter5_reg;
        p_read_10_reg_14832_pp0_iter7_reg <= p_read_10_reg_14832_pp0_iter6_reg;
        p_read_10_reg_14832_pp0_iter8_reg <= p_read_10_reg_14832_pp0_iter7_reg;
        p_read_10_reg_14832_pp0_iter9_reg <= p_read_10_reg_14832_pp0_iter8_reg;
        p_read_3_reg_14797_pp0_iter2_reg <= p_read_3_reg_14797_pp0_iter1_reg;
        p_read_4_reg_14802_pp0_iter2_reg <= p_read_4_reg_14802_pp0_iter1_reg;
        p_read_4_reg_14802_pp0_iter3_reg <= p_read_4_reg_14802_pp0_iter2_reg;
        p_read_4_reg_14802_pp0_iter4_reg <= p_read_4_reg_14802_pp0_iter3_reg;
        p_read_5_reg_14807_pp0_iter2_reg <= p_read_5_reg_14807_pp0_iter1_reg;
        p_read_5_reg_14807_pp0_iter3_reg <= p_read_5_reg_14807_pp0_iter2_reg;
        p_read_5_reg_14807_pp0_iter4_reg <= p_read_5_reg_14807_pp0_iter3_reg;
        p_read_5_reg_14807_pp0_iter5_reg <= p_read_5_reg_14807_pp0_iter4_reg;
        p_read_5_reg_14807_pp0_iter6_reg <= p_read_5_reg_14807_pp0_iter5_reg;
        p_read_6_reg_14812_pp0_iter2_reg <= p_read_6_reg_14812_pp0_iter1_reg;
        p_read_6_reg_14812_pp0_iter3_reg <= p_read_6_reg_14812_pp0_iter2_reg;
        p_read_6_reg_14812_pp0_iter4_reg <= p_read_6_reg_14812_pp0_iter3_reg;
        p_read_6_reg_14812_pp0_iter5_reg <= p_read_6_reg_14812_pp0_iter4_reg;
        p_read_6_reg_14812_pp0_iter6_reg <= p_read_6_reg_14812_pp0_iter5_reg;
        p_read_6_reg_14812_pp0_iter7_reg <= p_read_6_reg_14812_pp0_iter6_reg;
        p_read_6_reg_14812_pp0_iter8_reg <= p_read_6_reg_14812_pp0_iter7_reg;
        p_read_7_reg_14817_pp0_iter10_reg <= p_read_7_reg_14817_pp0_iter9_reg;
        p_read_7_reg_14817_pp0_iter2_reg <= p_read_7_reg_14817_pp0_iter1_reg;
        p_read_7_reg_14817_pp0_iter3_reg <= p_read_7_reg_14817_pp0_iter2_reg;
        p_read_7_reg_14817_pp0_iter4_reg <= p_read_7_reg_14817_pp0_iter3_reg;
        p_read_7_reg_14817_pp0_iter5_reg <= p_read_7_reg_14817_pp0_iter4_reg;
        p_read_7_reg_14817_pp0_iter6_reg <= p_read_7_reg_14817_pp0_iter5_reg;
        p_read_7_reg_14817_pp0_iter7_reg <= p_read_7_reg_14817_pp0_iter6_reg;
        p_read_7_reg_14817_pp0_iter8_reg <= p_read_7_reg_14817_pp0_iter7_reg;
        p_read_7_reg_14817_pp0_iter9_reg <= p_read_7_reg_14817_pp0_iter8_reg;
        p_read_8_reg_14822_pp0_iter10_reg <= p_read_8_reg_14822_pp0_iter9_reg;
        p_read_8_reg_14822_pp0_iter11_reg <= p_read_8_reg_14822_pp0_iter10_reg;
        p_read_8_reg_14822_pp0_iter12_reg <= p_read_8_reg_14822_pp0_iter11_reg;
        p_read_8_reg_14822_pp0_iter2_reg <= p_read_8_reg_14822_pp0_iter1_reg;
        p_read_8_reg_14822_pp0_iter3_reg <= p_read_8_reg_14822_pp0_iter2_reg;
        p_read_8_reg_14822_pp0_iter4_reg <= p_read_8_reg_14822_pp0_iter3_reg;
        p_read_8_reg_14822_pp0_iter5_reg <= p_read_8_reg_14822_pp0_iter4_reg;
        p_read_8_reg_14822_pp0_iter6_reg <= p_read_8_reg_14822_pp0_iter5_reg;
        p_read_8_reg_14822_pp0_iter7_reg <= p_read_8_reg_14822_pp0_iter6_reg;
        p_read_8_reg_14822_pp0_iter8_reg <= p_read_8_reg_14822_pp0_iter7_reg;
        p_read_8_reg_14822_pp0_iter9_reg <= p_read_8_reg_14822_pp0_iter8_reg;
        p_read_9_reg_14827_pp0_iter10_reg <= p_read_9_reg_14827_pp0_iter9_reg;
        p_read_9_reg_14827_pp0_iter11_reg <= p_read_9_reg_14827_pp0_iter10_reg;
        p_read_9_reg_14827_pp0_iter12_reg <= p_read_9_reg_14827_pp0_iter11_reg;
        p_read_9_reg_14827_pp0_iter13_reg <= p_read_9_reg_14827_pp0_iter12_reg;
        p_read_9_reg_14827_pp0_iter14_reg <= p_read_9_reg_14827_pp0_iter13_reg;
        p_read_9_reg_14827_pp0_iter2_reg <= p_read_9_reg_14827_pp0_iter1_reg;
        p_read_9_reg_14827_pp0_iter3_reg <= p_read_9_reg_14827_pp0_iter2_reg;
        p_read_9_reg_14827_pp0_iter4_reg <= p_read_9_reg_14827_pp0_iter3_reg;
        p_read_9_reg_14827_pp0_iter5_reg <= p_read_9_reg_14827_pp0_iter4_reg;
        p_read_9_reg_14827_pp0_iter6_reg <= p_read_9_reg_14827_pp0_iter5_reg;
        p_read_9_reg_14827_pp0_iter7_reg <= p_read_9_reg_14827_pp0_iter6_reg;
        p_read_9_reg_14827_pp0_iter8_reg <= p_read_9_reg_14827_pp0_iter7_reg;
        p_read_9_reg_14827_pp0_iter9_reg <= p_read_9_reg_14827_pp0_iter8_reg;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_idle_pp0 == 1'b1) & (ap_start == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter19 == 1'b0) & (ap_enable_reg_pp0_iter18 == 1'b0) & (ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b0) & (ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0_0to18 = 1'b1;
    end else begin
        ap_idle_pp0_0to18 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((ap_idle_pp0_0to18 == 1'b1) & (ap_start == 1'b0))) begin
        ap_reset_idle_pp0 = 1'b1;
    end else begin
        ap_reset_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce0 = 1'b1;
    end else begin
        decipher_0_i32box_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce1 = 1'b1;
    end else begin
        decipher_0_i32box_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce10 = 1'b1;
    end else begin
        decipher_0_i32box_ce10 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce100 = 1'b1;
    end else begin
        decipher_0_i32box_ce100 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce101 = 1'b1;
    end else begin
        decipher_0_i32box_ce101 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce102 = 1'b1;
    end else begin
        decipher_0_i32box_ce102 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce103 = 1'b1;
    end else begin
        decipher_0_i32box_ce103 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce104 = 1'b1;
    end else begin
        decipher_0_i32box_ce104 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce105 = 1'b1;
    end else begin
        decipher_0_i32box_ce105 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce106 = 1'b1;
    end else begin
        decipher_0_i32box_ce106 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce107 = 1'b1;
    end else begin
        decipher_0_i32box_ce107 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce108 = 1'b1;
    end else begin
        decipher_0_i32box_ce108 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce109 = 1'b1;
    end else begin
        decipher_0_i32box_ce109 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce11 = 1'b1;
    end else begin
        decipher_0_i32box_ce11 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce110 = 1'b1;
    end else begin
        decipher_0_i32box_ce110 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce111 = 1'b1;
    end else begin
        decipher_0_i32box_ce111 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce112 = 1'b1;
    end else begin
        decipher_0_i32box_ce112 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce113 = 1'b1;
    end else begin
        decipher_0_i32box_ce113 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce114 = 1'b1;
    end else begin
        decipher_0_i32box_ce114 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce115 = 1'b1;
    end else begin
        decipher_0_i32box_ce115 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce116 = 1'b1;
    end else begin
        decipher_0_i32box_ce116 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce117 = 1'b1;
    end else begin
        decipher_0_i32box_ce117 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce118 = 1'b1;
    end else begin
        decipher_0_i32box_ce118 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce119 = 1'b1;
    end else begin
        decipher_0_i32box_ce119 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce12 = 1'b1;
    end else begin
        decipher_0_i32box_ce12 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce120 = 1'b1;
    end else begin
        decipher_0_i32box_ce120 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce121 = 1'b1;
    end else begin
        decipher_0_i32box_ce121 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce122 = 1'b1;
    end else begin
        decipher_0_i32box_ce122 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce123 = 1'b1;
    end else begin
        decipher_0_i32box_ce123 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce124 = 1'b1;
    end else begin
        decipher_0_i32box_ce124 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce125 = 1'b1;
    end else begin
        decipher_0_i32box_ce125 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce126 = 1'b1;
    end else begin
        decipher_0_i32box_ce126 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce127 = 1'b1;
    end else begin
        decipher_0_i32box_ce127 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce128 = 1'b1;
    end else begin
        decipher_0_i32box_ce128 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce129 = 1'b1;
    end else begin
        decipher_0_i32box_ce129 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce13 = 1'b1;
    end else begin
        decipher_0_i32box_ce13 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce130 = 1'b1;
    end else begin
        decipher_0_i32box_ce130 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce131 = 1'b1;
    end else begin
        decipher_0_i32box_ce131 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce132 = 1'b1;
    end else begin
        decipher_0_i32box_ce132 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce133 = 1'b1;
    end else begin
        decipher_0_i32box_ce133 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce134 = 1'b1;
    end else begin
        decipher_0_i32box_ce134 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce135 = 1'b1;
    end else begin
        decipher_0_i32box_ce135 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce136 = 1'b1;
    end else begin
        decipher_0_i32box_ce136 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce137 = 1'b1;
    end else begin
        decipher_0_i32box_ce137 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce138 = 1'b1;
    end else begin
        decipher_0_i32box_ce138 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce139 = 1'b1;
    end else begin
        decipher_0_i32box_ce139 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce14 = 1'b1;
    end else begin
        decipher_0_i32box_ce14 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce140 = 1'b1;
    end else begin
        decipher_0_i32box_ce140 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce141 = 1'b1;
    end else begin
        decipher_0_i32box_ce141 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce142 = 1'b1;
    end else begin
        decipher_0_i32box_ce142 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce143 = 1'b1;
    end else begin
        decipher_0_i32box_ce143 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce15 = 1'b1;
    end else begin
        decipher_0_i32box_ce15 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce16 = 1'b1;
    end else begin
        decipher_0_i32box_ce16 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce17 = 1'b1;
    end else begin
        decipher_0_i32box_ce17 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce18 = 1'b1;
    end else begin
        decipher_0_i32box_ce18 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce19 = 1'b1;
    end else begin
        decipher_0_i32box_ce19 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce2 = 1'b1;
    end else begin
        decipher_0_i32box_ce2 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce20 = 1'b1;
    end else begin
        decipher_0_i32box_ce20 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce21 = 1'b1;
    end else begin
        decipher_0_i32box_ce21 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce22 = 1'b1;
    end else begin
        decipher_0_i32box_ce22 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce23 = 1'b1;
    end else begin
        decipher_0_i32box_ce23 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce24 = 1'b1;
    end else begin
        decipher_0_i32box_ce24 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce25 = 1'b1;
    end else begin
        decipher_0_i32box_ce25 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce26 = 1'b1;
    end else begin
        decipher_0_i32box_ce26 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce27 = 1'b1;
    end else begin
        decipher_0_i32box_ce27 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce28 = 1'b1;
    end else begin
        decipher_0_i32box_ce28 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce29 = 1'b1;
    end else begin
        decipher_0_i32box_ce29 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce3 = 1'b1;
    end else begin
        decipher_0_i32box_ce3 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce30 = 1'b1;
    end else begin
        decipher_0_i32box_ce30 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce31 = 1'b1;
    end else begin
        decipher_0_i32box_ce31 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce32 = 1'b1;
    end else begin
        decipher_0_i32box_ce32 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce33 = 1'b1;
    end else begin
        decipher_0_i32box_ce33 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce34 = 1'b1;
    end else begin
        decipher_0_i32box_ce34 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce35 = 1'b1;
    end else begin
        decipher_0_i32box_ce35 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce36 = 1'b1;
    end else begin
        decipher_0_i32box_ce36 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce37 = 1'b1;
    end else begin
        decipher_0_i32box_ce37 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce38 = 1'b1;
    end else begin
        decipher_0_i32box_ce38 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce39 = 1'b1;
    end else begin
        decipher_0_i32box_ce39 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce4 = 1'b1;
    end else begin
        decipher_0_i32box_ce4 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce40 = 1'b1;
    end else begin
        decipher_0_i32box_ce40 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce41 = 1'b1;
    end else begin
        decipher_0_i32box_ce41 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce42 = 1'b1;
    end else begin
        decipher_0_i32box_ce42 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce43 = 1'b1;
    end else begin
        decipher_0_i32box_ce43 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce44 = 1'b1;
    end else begin
        decipher_0_i32box_ce44 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce45 = 1'b1;
    end else begin
        decipher_0_i32box_ce45 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce46 = 1'b1;
    end else begin
        decipher_0_i32box_ce46 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce47 = 1'b1;
    end else begin
        decipher_0_i32box_ce47 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce48 = 1'b1;
    end else begin
        decipher_0_i32box_ce48 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce49 = 1'b1;
    end else begin
        decipher_0_i32box_ce49 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce5 = 1'b1;
    end else begin
        decipher_0_i32box_ce5 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce50 = 1'b1;
    end else begin
        decipher_0_i32box_ce50 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce51 = 1'b1;
    end else begin
        decipher_0_i32box_ce51 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce52 = 1'b1;
    end else begin
        decipher_0_i32box_ce52 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce53 = 1'b1;
    end else begin
        decipher_0_i32box_ce53 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce54 = 1'b1;
    end else begin
        decipher_0_i32box_ce54 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce55 = 1'b1;
    end else begin
        decipher_0_i32box_ce55 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce56 = 1'b1;
    end else begin
        decipher_0_i32box_ce56 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce57 = 1'b1;
    end else begin
        decipher_0_i32box_ce57 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce58 = 1'b1;
    end else begin
        decipher_0_i32box_ce58 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce59 = 1'b1;
    end else begin
        decipher_0_i32box_ce59 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce6 = 1'b1;
    end else begin
        decipher_0_i32box_ce6 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce60 = 1'b1;
    end else begin
        decipher_0_i32box_ce60 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce61 = 1'b1;
    end else begin
        decipher_0_i32box_ce61 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce62 = 1'b1;
    end else begin
        decipher_0_i32box_ce62 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce63 = 1'b1;
    end else begin
        decipher_0_i32box_ce63 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce64 = 1'b1;
    end else begin
        decipher_0_i32box_ce64 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce65 = 1'b1;
    end else begin
        decipher_0_i32box_ce65 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce66 = 1'b1;
    end else begin
        decipher_0_i32box_ce66 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce67 = 1'b1;
    end else begin
        decipher_0_i32box_ce67 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce68 = 1'b1;
    end else begin
        decipher_0_i32box_ce68 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce69 = 1'b1;
    end else begin
        decipher_0_i32box_ce69 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce7 = 1'b1;
    end else begin
        decipher_0_i32box_ce7 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce70 = 1'b1;
    end else begin
        decipher_0_i32box_ce70 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce71 = 1'b1;
    end else begin
        decipher_0_i32box_ce71 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce72 = 1'b1;
    end else begin
        decipher_0_i32box_ce72 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce73 = 1'b1;
    end else begin
        decipher_0_i32box_ce73 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce74 = 1'b1;
    end else begin
        decipher_0_i32box_ce74 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce75 = 1'b1;
    end else begin
        decipher_0_i32box_ce75 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce76 = 1'b1;
    end else begin
        decipher_0_i32box_ce76 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce77 = 1'b1;
    end else begin
        decipher_0_i32box_ce77 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce78 = 1'b1;
    end else begin
        decipher_0_i32box_ce78 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce79 = 1'b1;
    end else begin
        decipher_0_i32box_ce79 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce8 = 1'b1;
    end else begin
        decipher_0_i32box_ce8 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce80 = 1'b1;
    end else begin
        decipher_0_i32box_ce80 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce81 = 1'b1;
    end else begin
        decipher_0_i32box_ce81 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce82 = 1'b1;
    end else begin
        decipher_0_i32box_ce82 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce83 = 1'b1;
    end else begin
        decipher_0_i32box_ce83 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce84 = 1'b1;
    end else begin
        decipher_0_i32box_ce84 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce85 = 1'b1;
    end else begin
        decipher_0_i32box_ce85 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce86 = 1'b1;
    end else begin
        decipher_0_i32box_ce86 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce87 = 1'b1;
    end else begin
        decipher_0_i32box_ce87 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce88 = 1'b1;
    end else begin
        decipher_0_i32box_ce88 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce89 = 1'b1;
    end else begin
        decipher_0_i32box_ce89 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce9 = 1'b1;
    end else begin
        decipher_0_i32box_ce9 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce90 = 1'b1;
    end else begin
        decipher_0_i32box_ce90 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce91 = 1'b1;
    end else begin
        decipher_0_i32box_ce91 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce92 = 1'b1;
    end else begin
        decipher_0_i32box_ce92 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce93 = 1'b1;
    end else begin
        decipher_0_i32box_ce93 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce94 = 1'b1;
    end else begin
        decipher_0_i32box_ce94 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce95 = 1'b1;
    end else begin
        decipher_0_i32box_ce95 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce96 = 1'b1;
    end else begin
        decipher_0_i32box_ce96 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce97 = 1'b1;
    end else begin
        decipher_0_i32box_ce97 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce98 = 1'b1;
    end else begin
        decipher_0_i32box_ce98 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_i32box_ce99 = 1'b1;
    end else begin
        decipher_0_i32box_ce99 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce0 = 1'b1;
    end else begin
        decipher_0_iibox_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce1 = 1'b1;
    end else begin
        decipher_0_iibox_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce10 = 1'b1;
    end else begin
        decipher_0_iibox_ce10 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce100 = 1'b1;
    end else begin
        decipher_0_iibox_ce100 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce101 = 1'b1;
    end else begin
        decipher_0_iibox_ce101 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce102 = 1'b1;
    end else begin
        decipher_0_iibox_ce102 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce103 = 1'b1;
    end else begin
        decipher_0_iibox_ce103 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce104 = 1'b1;
    end else begin
        decipher_0_iibox_ce104 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce105 = 1'b1;
    end else begin
        decipher_0_iibox_ce105 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce106 = 1'b1;
    end else begin
        decipher_0_iibox_ce106 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce107 = 1'b1;
    end else begin
        decipher_0_iibox_ce107 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce108 = 1'b1;
    end else begin
        decipher_0_iibox_ce108 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce109 = 1'b1;
    end else begin
        decipher_0_iibox_ce109 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce11 = 1'b1;
    end else begin
        decipher_0_iibox_ce11 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce110 = 1'b1;
    end else begin
        decipher_0_iibox_ce110 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce111 = 1'b1;
    end else begin
        decipher_0_iibox_ce111 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce112 = 1'b1;
    end else begin
        decipher_0_iibox_ce112 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce113 = 1'b1;
    end else begin
        decipher_0_iibox_ce113 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce114 = 1'b1;
    end else begin
        decipher_0_iibox_ce114 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce115 = 1'b1;
    end else begin
        decipher_0_iibox_ce115 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce116 = 1'b1;
    end else begin
        decipher_0_iibox_ce116 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce117 = 1'b1;
    end else begin
        decipher_0_iibox_ce117 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce118 = 1'b1;
    end else begin
        decipher_0_iibox_ce118 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce119 = 1'b1;
    end else begin
        decipher_0_iibox_ce119 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce12 = 1'b1;
    end else begin
        decipher_0_iibox_ce12 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce120 = 1'b1;
    end else begin
        decipher_0_iibox_ce120 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce121 = 1'b1;
    end else begin
        decipher_0_iibox_ce121 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce122 = 1'b1;
    end else begin
        decipher_0_iibox_ce122 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce123 = 1'b1;
    end else begin
        decipher_0_iibox_ce123 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce124 = 1'b1;
    end else begin
        decipher_0_iibox_ce124 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce125 = 1'b1;
    end else begin
        decipher_0_iibox_ce125 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce126 = 1'b1;
    end else begin
        decipher_0_iibox_ce126 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce127 = 1'b1;
    end else begin
        decipher_0_iibox_ce127 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce128 = 1'b1;
    end else begin
        decipher_0_iibox_ce128 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce129 = 1'b1;
    end else begin
        decipher_0_iibox_ce129 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce13 = 1'b1;
    end else begin
        decipher_0_iibox_ce13 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce130 = 1'b1;
    end else begin
        decipher_0_iibox_ce130 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce131 = 1'b1;
    end else begin
        decipher_0_iibox_ce131 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce132 = 1'b1;
    end else begin
        decipher_0_iibox_ce132 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce133 = 1'b1;
    end else begin
        decipher_0_iibox_ce133 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce134 = 1'b1;
    end else begin
        decipher_0_iibox_ce134 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce135 = 1'b1;
    end else begin
        decipher_0_iibox_ce135 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce136 = 1'b1;
    end else begin
        decipher_0_iibox_ce136 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce137 = 1'b1;
    end else begin
        decipher_0_iibox_ce137 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce138 = 1'b1;
    end else begin
        decipher_0_iibox_ce138 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce139 = 1'b1;
    end else begin
        decipher_0_iibox_ce139 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce14 = 1'b1;
    end else begin
        decipher_0_iibox_ce14 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce140 = 1'b1;
    end else begin
        decipher_0_iibox_ce140 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce141 = 1'b1;
    end else begin
        decipher_0_iibox_ce141 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce142 = 1'b1;
    end else begin
        decipher_0_iibox_ce142 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce143 = 1'b1;
    end else begin
        decipher_0_iibox_ce143 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce144 = 1'b1;
    end else begin
        decipher_0_iibox_ce144 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce145 = 1'b1;
    end else begin
        decipher_0_iibox_ce145 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce146 = 1'b1;
    end else begin
        decipher_0_iibox_ce146 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce147 = 1'b1;
    end else begin
        decipher_0_iibox_ce147 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce148 = 1'b1;
    end else begin
        decipher_0_iibox_ce148 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce149 = 1'b1;
    end else begin
        decipher_0_iibox_ce149 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce15 = 1'b1;
    end else begin
        decipher_0_iibox_ce15 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce150 = 1'b1;
    end else begin
        decipher_0_iibox_ce150 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce151 = 1'b1;
    end else begin
        decipher_0_iibox_ce151 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce152 = 1'b1;
    end else begin
        decipher_0_iibox_ce152 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce153 = 1'b1;
    end else begin
        decipher_0_iibox_ce153 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce154 = 1'b1;
    end else begin
        decipher_0_iibox_ce154 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce155 = 1'b1;
    end else begin
        decipher_0_iibox_ce155 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce156 = 1'b1;
    end else begin
        decipher_0_iibox_ce156 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce157 = 1'b1;
    end else begin
        decipher_0_iibox_ce157 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce158 = 1'b1;
    end else begin
        decipher_0_iibox_ce158 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce159 = 1'b1;
    end else begin
        decipher_0_iibox_ce159 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce16 = 1'b1;
    end else begin
        decipher_0_iibox_ce16 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce17 = 1'b1;
    end else begin
        decipher_0_iibox_ce17 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce18 = 1'b1;
    end else begin
        decipher_0_iibox_ce18 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce19 = 1'b1;
    end else begin
        decipher_0_iibox_ce19 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce2 = 1'b1;
    end else begin
        decipher_0_iibox_ce2 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce20 = 1'b1;
    end else begin
        decipher_0_iibox_ce20 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce21 = 1'b1;
    end else begin
        decipher_0_iibox_ce21 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce22 = 1'b1;
    end else begin
        decipher_0_iibox_ce22 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce23 = 1'b1;
    end else begin
        decipher_0_iibox_ce23 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce24 = 1'b1;
    end else begin
        decipher_0_iibox_ce24 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce25 = 1'b1;
    end else begin
        decipher_0_iibox_ce25 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce26 = 1'b1;
    end else begin
        decipher_0_iibox_ce26 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce27 = 1'b1;
    end else begin
        decipher_0_iibox_ce27 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce28 = 1'b1;
    end else begin
        decipher_0_iibox_ce28 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce29 = 1'b1;
    end else begin
        decipher_0_iibox_ce29 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce3 = 1'b1;
    end else begin
        decipher_0_iibox_ce3 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce30 = 1'b1;
    end else begin
        decipher_0_iibox_ce30 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce31 = 1'b1;
    end else begin
        decipher_0_iibox_ce31 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce32 = 1'b1;
    end else begin
        decipher_0_iibox_ce32 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce33 = 1'b1;
    end else begin
        decipher_0_iibox_ce33 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce34 = 1'b1;
    end else begin
        decipher_0_iibox_ce34 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce35 = 1'b1;
    end else begin
        decipher_0_iibox_ce35 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce36 = 1'b1;
    end else begin
        decipher_0_iibox_ce36 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce37 = 1'b1;
    end else begin
        decipher_0_iibox_ce37 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce38 = 1'b1;
    end else begin
        decipher_0_iibox_ce38 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce39 = 1'b1;
    end else begin
        decipher_0_iibox_ce39 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce4 = 1'b1;
    end else begin
        decipher_0_iibox_ce4 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce40 = 1'b1;
    end else begin
        decipher_0_iibox_ce40 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce41 = 1'b1;
    end else begin
        decipher_0_iibox_ce41 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce42 = 1'b1;
    end else begin
        decipher_0_iibox_ce42 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce43 = 1'b1;
    end else begin
        decipher_0_iibox_ce43 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce44 = 1'b1;
    end else begin
        decipher_0_iibox_ce44 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce45 = 1'b1;
    end else begin
        decipher_0_iibox_ce45 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce46 = 1'b1;
    end else begin
        decipher_0_iibox_ce46 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce47 = 1'b1;
    end else begin
        decipher_0_iibox_ce47 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce48 = 1'b1;
    end else begin
        decipher_0_iibox_ce48 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce49 = 1'b1;
    end else begin
        decipher_0_iibox_ce49 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce5 = 1'b1;
    end else begin
        decipher_0_iibox_ce5 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce50 = 1'b1;
    end else begin
        decipher_0_iibox_ce50 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce51 = 1'b1;
    end else begin
        decipher_0_iibox_ce51 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce52 = 1'b1;
    end else begin
        decipher_0_iibox_ce52 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce53 = 1'b1;
    end else begin
        decipher_0_iibox_ce53 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce54 = 1'b1;
    end else begin
        decipher_0_iibox_ce54 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce55 = 1'b1;
    end else begin
        decipher_0_iibox_ce55 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce56 = 1'b1;
    end else begin
        decipher_0_iibox_ce56 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce57 = 1'b1;
    end else begin
        decipher_0_iibox_ce57 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce58 = 1'b1;
    end else begin
        decipher_0_iibox_ce58 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce59 = 1'b1;
    end else begin
        decipher_0_iibox_ce59 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce6 = 1'b1;
    end else begin
        decipher_0_iibox_ce6 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce60 = 1'b1;
    end else begin
        decipher_0_iibox_ce60 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce61 = 1'b1;
    end else begin
        decipher_0_iibox_ce61 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce62 = 1'b1;
    end else begin
        decipher_0_iibox_ce62 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce63 = 1'b1;
    end else begin
        decipher_0_iibox_ce63 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce64 = 1'b1;
    end else begin
        decipher_0_iibox_ce64 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce65 = 1'b1;
    end else begin
        decipher_0_iibox_ce65 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce66 = 1'b1;
    end else begin
        decipher_0_iibox_ce66 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce67 = 1'b1;
    end else begin
        decipher_0_iibox_ce67 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce68 = 1'b1;
    end else begin
        decipher_0_iibox_ce68 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce69 = 1'b1;
    end else begin
        decipher_0_iibox_ce69 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce7 = 1'b1;
    end else begin
        decipher_0_iibox_ce7 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce70 = 1'b1;
    end else begin
        decipher_0_iibox_ce70 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce71 = 1'b1;
    end else begin
        decipher_0_iibox_ce71 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce72 = 1'b1;
    end else begin
        decipher_0_iibox_ce72 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce73 = 1'b1;
    end else begin
        decipher_0_iibox_ce73 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce74 = 1'b1;
    end else begin
        decipher_0_iibox_ce74 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce75 = 1'b1;
    end else begin
        decipher_0_iibox_ce75 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce76 = 1'b1;
    end else begin
        decipher_0_iibox_ce76 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce77 = 1'b1;
    end else begin
        decipher_0_iibox_ce77 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce78 = 1'b1;
    end else begin
        decipher_0_iibox_ce78 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce79 = 1'b1;
    end else begin
        decipher_0_iibox_ce79 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce8 = 1'b1;
    end else begin
        decipher_0_iibox_ce8 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce80 = 1'b1;
    end else begin
        decipher_0_iibox_ce80 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce81 = 1'b1;
    end else begin
        decipher_0_iibox_ce81 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce82 = 1'b1;
    end else begin
        decipher_0_iibox_ce82 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce83 = 1'b1;
    end else begin
        decipher_0_iibox_ce83 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce84 = 1'b1;
    end else begin
        decipher_0_iibox_ce84 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce85 = 1'b1;
    end else begin
        decipher_0_iibox_ce85 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce86 = 1'b1;
    end else begin
        decipher_0_iibox_ce86 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce87 = 1'b1;
    end else begin
        decipher_0_iibox_ce87 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce88 = 1'b1;
    end else begin
        decipher_0_iibox_ce88 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce89 = 1'b1;
    end else begin
        decipher_0_iibox_ce89 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce9 = 1'b1;
    end else begin
        decipher_0_iibox_ce9 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce90 = 1'b1;
    end else begin
        decipher_0_iibox_ce90 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce91 = 1'b1;
    end else begin
        decipher_0_iibox_ce91 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce92 = 1'b1;
    end else begin
        decipher_0_iibox_ce92 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce93 = 1'b1;
    end else begin
        decipher_0_iibox_ce93 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce94 = 1'b1;
    end else begin
        decipher_0_iibox_ce94 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce95 = 1'b1;
    end else begin
        decipher_0_iibox_ce95 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce96 = 1'b1;
    end else begin
        decipher_0_iibox_ce96 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce97 = 1'b1;
    end else begin
        decipher_0_iibox_ce97 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce98 = 1'b1;
    end else begin
        decipher_0_iibox_ce98 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        decipher_0_iibox_ce99 = 1'b1;
    end else begin
        decipher_0_iibox_ce99 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_state10_pp0_stage0_iter9 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage0_iter10 = ~(1'b1 == 1'b1);

assign ap_block_state12_pp0_stage0_iter11 = ~(1'b1 == 1'b1);

assign ap_block_state13_pp0_stage0_iter12 = ~(1'b1 == 1'b1);

assign ap_block_state14_pp0_stage0_iter13 = ~(1'b1 == 1'b1);

assign ap_block_state15_pp0_stage0_iter14 = ~(1'b1 == 1'b1);

assign ap_block_state16_pp0_stage0_iter15 = ~(1'b1 == 1'b1);

assign ap_block_state17_pp0_stage0_iter16 = ~(1'b1 == 1'b1);

assign ap_block_state18_pp0_stage0_iter17 = ~(1'b1 == 1'b1);

assign ap_block_state19_pp0_stage0_iter18 = ~(1'b1 == 1'b1);

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state20_pp0_stage0_iter19 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter8 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_enable_reg_pp0_iter0 = ap_start;

assign ap_return = (p_read11_reg_14837_pp0_iter18_reg ^ p_Result_10_fu_14751_p17);

assign decipher_0_i32box_address0 = zext_ln708_290_fu_13834_p1;

assign decipher_0_i32box_address1 = zext_ln708_289_fu_13819_p1;

assign decipher_0_i32box_address10 = zext_ln708_280_fu_13684_p1;

assign decipher_0_i32box_address100 = zext_ln708_94_fu_6652_p1;

assign decipher_0_i32box_address101 = zext_ln708_93_fu_6637_p1;

assign decipher_0_i32box_address102 = zext_ln708_92_fu_6622_p1;

assign decipher_0_i32box_address103 = zext_ln708_91_fu_6607_p1;

assign decipher_0_i32box_address104 = zext_ln708_90_fu_6592_p1;

assign decipher_0_i32box_address105 = zext_ln708_89_fu_6577_p1;

assign decipher_0_i32box_address106 = zext_ln708_88_fu_6562_p1;

assign decipher_0_i32box_address107 = zext_ln708_87_fu_6547_p1;

assign decipher_0_i32box_address108 = zext_ln708_86_fu_6532_p1;

assign decipher_0_i32box_address109 = zext_ln708_85_fu_6517_p1;

assign decipher_0_i32box_address11 = zext_ln708_279_fu_13669_p1;

assign decipher_0_i32box_address110 = zext_ln708_84_fu_6502_p1;

assign decipher_0_i32box_address111 = zext_ln708_83_fu_6487_p1;

assign decipher_0_i32box_address112 = zext_ln708_66_fu_5525_p1;

assign decipher_0_i32box_address113 = zext_ln708_65_fu_5510_p1;

assign decipher_0_i32box_address114 = zext_ln708_64_fu_5495_p1;

assign decipher_0_i32box_address115 = zext_ln708_63_fu_5480_p1;

assign decipher_0_i32box_address116 = zext_ln708_62_fu_5465_p1;

assign decipher_0_i32box_address117 = zext_ln708_61_fu_5450_p1;

assign decipher_0_i32box_address118 = zext_ln708_60_fu_5435_p1;

assign decipher_0_i32box_address119 = zext_ln708_59_fu_5420_p1;

assign decipher_0_i32box_address12 = zext_ln708_278_fu_13654_p1;

assign decipher_0_i32box_address120 = zext_ln708_58_fu_5405_p1;

assign decipher_0_i32box_address121 = zext_ln708_57_fu_5390_p1;

assign decipher_0_i32box_address122 = zext_ln708_56_fu_5375_p1;

assign decipher_0_i32box_address123 = zext_ln708_55_fu_5360_p1;

assign decipher_0_i32box_address124 = zext_ln708_54_fu_5345_p1;

assign decipher_0_i32box_address125 = zext_ln708_53_fu_5330_p1;

assign decipher_0_i32box_address126 = zext_ln708_52_fu_5315_p1;

assign decipher_0_i32box_address127 = zext_ln708_51_fu_5300_p1;

assign decipher_0_i32box_address128 = zext_ln708_34_fu_4338_p1;

assign decipher_0_i32box_address129 = zext_ln708_33_fu_4323_p1;

assign decipher_0_i32box_address13 = zext_ln708_277_fu_13639_p1;

assign decipher_0_i32box_address130 = zext_ln708_32_fu_4308_p1;

assign decipher_0_i32box_address131 = zext_ln708_31_fu_4293_p1;

assign decipher_0_i32box_address132 = zext_ln708_30_fu_4278_p1;

assign decipher_0_i32box_address133 = zext_ln708_29_fu_4263_p1;

assign decipher_0_i32box_address134 = zext_ln708_28_fu_4248_p1;

assign decipher_0_i32box_address135 = zext_ln708_27_fu_4233_p1;

assign decipher_0_i32box_address136 = zext_ln708_26_fu_4218_p1;

assign decipher_0_i32box_address137 = zext_ln708_25_fu_4203_p1;

assign decipher_0_i32box_address138 = zext_ln708_24_fu_4188_p1;

assign decipher_0_i32box_address139 = zext_ln708_23_fu_4173_p1;

assign decipher_0_i32box_address14 = zext_ln708_276_fu_13624_p1;

assign decipher_0_i32box_address140 = zext_ln708_22_fu_4158_p1;

assign decipher_0_i32box_address141 = zext_ln708_21_fu_4143_p1;

assign decipher_0_i32box_address142 = zext_ln708_20_fu_4128_p1;

assign decipher_0_i32box_address143 = zext_ln708_19_fu_4113_p1;

assign decipher_0_i32box_address15 = zext_ln708_275_fu_13609_p1;

assign decipher_0_i32box_address16 = zext_ln708_258_fu_12647_p1;

assign decipher_0_i32box_address17 = zext_ln708_257_fu_12632_p1;

assign decipher_0_i32box_address18 = zext_ln708_256_fu_12617_p1;

assign decipher_0_i32box_address19 = zext_ln708_255_fu_12602_p1;

assign decipher_0_i32box_address2 = zext_ln708_288_fu_13804_p1;

assign decipher_0_i32box_address20 = zext_ln708_254_fu_12587_p1;

assign decipher_0_i32box_address21 = zext_ln708_253_fu_12572_p1;

assign decipher_0_i32box_address22 = zext_ln708_252_fu_12557_p1;

assign decipher_0_i32box_address23 = zext_ln708_251_fu_12542_p1;

assign decipher_0_i32box_address24 = zext_ln708_250_fu_12527_p1;

assign decipher_0_i32box_address25 = zext_ln708_249_fu_12512_p1;

assign decipher_0_i32box_address26 = zext_ln708_248_fu_12497_p1;

assign decipher_0_i32box_address27 = zext_ln708_247_fu_12482_p1;

assign decipher_0_i32box_address28 = zext_ln708_246_fu_12467_p1;

assign decipher_0_i32box_address29 = zext_ln708_245_fu_12452_p1;

assign decipher_0_i32box_address3 = zext_ln708_287_fu_13789_p1;

assign decipher_0_i32box_address30 = zext_ln708_244_fu_12437_p1;

assign decipher_0_i32box_address31 = zext_ln708_243_fu_12422_p1;

assign decipher_0_i32box_address32 = zext_ln708_226_fu_11460_p1;

assign decipher_0_i32box_address33 = zext_ln708_225_fu_11445_p1;

assign decipher_0_i32box_address34 = zext_ln708_224_fu_11430_p1;

assign decipher_0_i32box_address35 = zext_ln708_223_fu_11415_p1;

assign decipher_0_i32box_address36 = zext_ln708_222_fu_11400_p1;

assign decipher_0_i32box_address37 = zext_ln708_221_fu_11385_p1;

assign decipher_0_i32box_address38 = zext_ln708_220_fu_11370_p1;

assign decipher_0_i32box_address39 = zext_ln708_219_fu_11355_p1;

assign decipher_0_i32box_address4 = zext_ln708_286_fu_13774_p1;

assign decipher_0_i32box_address40 = zext_ln708_218_fu_11340_p1;

assign decipher_0_i32box_address41 = zext_ln708_217_fu_11325_p1;

assign decipher_0_i32box_address42 = zext_ln708_216_fu_11310_p1;

assign decipher_0_i32box_address43 = zext_ln708_215_fu_11295_p1;

assign decipher_0_i32box_address44 = zext_ln708_214_fu_11280_p1;

assign decipher_0_i32box_address45 = zext_ln708_213_fu_11265_p1;

assign decipher_0_i32box_address46 = zext_ln708_212_fu_11250_p1;

assign decipher_0_i32box_address47 = zext_ln708_211_fu_11235_p1;

assign decipher_0_i32box_address48 = zext_ln708_194_fu_10273_p1;

assign decipher_0_i32box_address49 = zext_ln708_193_fu_10258_p1;

assign decipher_0_i32box_address5 = zext_ln708_285_fu_13759_p1;

assign decipher_0_i32box_address50 = zext_ln708_192_fu_10243_p1;

assign decipher_0_i32box_address51 = zext_ln708_191_fu_10228_p1;

assign decipher_0_i32box_address52 = zext_ln708_190_fu_10213_p1;

assign decipher_0_i32box_address53 = zext_ln708_189_fu_10198_p1;

assign decipher_0_i32box_address54 = zext_ln708_188_fu_10183_p1;

assign decipher_0_i32box_address55 = zext_ln708_187_fu_10168_p1;

assign decipher_0_i32box_address56 = zext_ln708_186_fu_10153_p1;

assign decipher_0_i32box_address57 = zext_ln708_185_fu_10138_p1;

assign decipher_0_i32box_address58 = zext_ln708_184_fu_10123_p1;

assign decipher_0_i32box_address59 = zext_ln708_183_fu_10108_p1;

assign decipher_0_i32box_address6 = zext_ln708_284_fu_13744_p1;

assign decipher_0_i32box_address60 = zext_ln708_182_fu_10093_p1;

assign decipher_0_i32box_address61 = zext_ln708_181_fu_10078_p1;

assign decipher_0_i32box_address62 = zext_ln708_180_fu_10063_p1;

assign decipher_0_i32box_address63 = zext_ln708_179_fu_10048_p1;

assign decipher_0_i32box_address64 = zext_ln708_162_fu_9086_p1;

assign decipher_0_i32box_address65 = zext_ln708_161_fu_9071_p1;

assign decipher_0_i32box_address66 = zext_ln708_160_fu_9056_p1;

assign decipher_0_i32box_address67 = zext_ln708_159_fu_9041_p1;

assign decipher_0_i32box_address68 = zext_ln708_158_fu_9026_p1;

assign decipher_0_i32box_address69 = zext_ln708_157_fu_9011_p1;

assign decipher_0_i32box_address7 = zext_ln708_283_fu_13729_p1;

assign decipher_0_i32box_address70 = zext_ln708_156_fu_8996_p1;

assign decipher_0_i32box_address71 = zext_ln708_155_fu_8981_p1;

assign decipher_0_i32box_address72 = zext_ln708_154_fu_8966_p1;

assign decipher_0_i32box_address73 = zext_ln708_153_fu_8951_p1;

assign decipher_0_i32box_address74 = zext_ln708_152_fu_8936_p1;

assign decipher_0_i32box_address75 = zext_ln708_151_fu_8921_p1;

assign decipher_0_i32box_address76 = zext_ln708_150_fu_8906_p1;

assign decipher_0_i32box_address77 = zext_ln708_149_fu_8891_p1;

assign decipher_0_i32box_address78 = zext_ln708_148_fu_8876_p1;

assign decipher_0_i32box_address79 = zext_ln708_147_fu_8861_p1;

assign decipher_0_i32box_address8 = zext_ln708_282_fu_13714_p1;

assign decipher_0_i32box_address80 = zext_ln708_130_fu_7899_p1;

assign decipher_0_i32box_address81 = zext_ln708_129_fu_7884_p1;

assign decipher_0_i32box_address82 = zext_ln708_128_fu_7869_p1;

assign decipher_0_i32box_address83 = zext_ln708_127_fu_7854_p1;

assign decipher_0_i32box_address84 = zext_ln708_126_fu_7839_p1;

assign decipher_0_i32box_address85 = zext_ln708_125_fu_7824_p1;

assign decipher_0_i32box_address86 = zext_ln708_124_fu_7809_p1;

assign decipher_0_i32box_address87 = zext_ln708_123_fu_7794_p1;

assign decipher_0_i32box_address88 = zext_ln708_122_fu_7779_p1;

assign decipher_0_i32box_address89 = zext_ln708_121_fu_7764_p1;

assign decipher_0_i32box_address9 = zext_ln708_281_fu_13699_p1;

assign decipher_0_i32box_address90 = zext_ln708_120_fu_7749_p1;

assign decipher_0_i32box_address91 = zext_ln708_119_fu_7734_p1;

assign decipher_0_i32box_address92 = zext_ln708_118_fu_7719_p1;

assign decipher_0_i32box_address93 = zext_ln708_117_fu_7704_p1;

assign decipher_0_i32box_address94 = zext_ln708_116_fu_7689_p1;

assign decipher_0_i32box_address95 = zext_ln708_115_fu_7674_p1;

assign decipher_0_i32box_address96 = zext_ln708_98_fu_6712_p1;

assign decipher_0_i32box_address97 = zext_ln708_97_fu_6697_p1;

assign decipher_0_i32box_address98 = zext_ln708_96_fu_6682_p1;

assign decipher_0_i32box_address99 = zext_ln708_95_fu_6667_p1;

assign decipher_0_iibox_address0 = zext_ln708_306_fu_14746_p1;

assign decipher_0_iibox_address1 = zext_ln708_305_fu_14741_p1;

assign decipher_0_iibox_address10 = zext_ln708_296_fu_14696_p1;

assign decipher_0_iibox_address100 = zext_ln708_110_fu_7604_p1;

assign decipher_0_iibox_address101 = zext_ln708_109_fu_7599_p1;

assign decipher_0_iibox_address102 = zext_ln708_108_fu_7594_p1;

assign decipher_0_iibox_address103 = zext_ln708_107_fu_7589_p1;

assign decipher_0_iibox_address104 = zext_ln708_106_fu_7584_p1;

assign decipher_0_iibox_address105 = zext_ln708_105_fu_7579_p1;

assign decipher_0_iibox_address106 = zext_ln708_104_fu_7574_p1;

assign decipher_0_iibox_address107 = zext_ln708_103_fu_7569_p1;

assign decipher_0_iibox_address108 = zext_ln708_102_fu_7564_p1;

assign decipher_0_iibox_address109 = zext_ln708_101_fu_7559_p1;

assign decipher_0_iibox_address11 = zext_ln708_295_fu_14691_p1;

assign decipher_0_iibox_address110 = zext_ln708_100_fu_7554_p1;

assign decipher_0_iibox_address111 = zext_ln708_99_fu_7549_p1;

assign decipher_0_iibox_address112 = zext_ln708_82_fu_6437_p1;

assign decipher_0_iibox_address113 = zext_ln708_81_fu_6432_p1;

assign decipher_0_iibox_address114 = zext_ln708_80_fu_6427_p1;

assign decipher_0_iibox_address115 = zext_ln708_79_fu_6422_p1;

assign decipher_0_iibox_address116 = zext_ln708_78_fu_6417_p1;

assign decipher_0_iibox_address117 = zext_ln708_77_fu_6412_p1;

assign decipher_0_iibox_address118 = zext_ln708_76_fu_6407_p1;

assign decipher_0_iibox_address119 = zext_ln708_75_fu_6402_p1;

assign decipher_0_iibox_address12 = zext_ln708_294_fu_14686_p1;

assign decipher_0_iibox_address120 = zext_ln708_74_fu_6397_p1;

assign decipher_0_iibox_address121 = zext_ln708_73_fu_6392_p1;

assign decipher_0_iibox_address122 = zext_ln708_72_fu_6387_p1;

assign decipher_0_iibox_address123 = zext_ln708_71_fu_6382_p1;

assign decipher_0_iibox_address124 = zext_ln708_70_fu_6377_p1;

assign decipher_0_iibox_address125 = zext_ln708_69_fu_6372_p1;

assign decipher_0_iibox_address126 = zext_ln708_68_fu_6367_p1;

assign decipher_0_iibox_address127 = zext_ln708_67_fu_6362_p1;

assign decipher_0_iibox_address128 = zext_ln708_50_fu_5250_p1;

assign decipher_0_iibox_address129 = zext_ln708_49_fu_5245_p1;

assign decipher_0_iibox_address13 = zext_ln708_293_fu_14681_p1;

assign decipher_0_iibox_address130 = zext_ln708_48_fu_5240_p1;

assign decipher_0_iibox_address131 = zext_ln708_47_fu_5235_p1;

assign decipher_0_iibox_address132 = zext_ln708_46_fu_5230_p1;

assign decipher_0_iibox_address133 = zext_ln708_45_fu_5225_p1;

assign decipher_0_iibox_address134 = zext_ln708_44_fu_5220_p1;

assign decipher_0_iibox_address135 = zext_ln708_43_fu_5215_p1;

assign decipher_0_iibox_address136 = zext_ln708_42_fu_5210_p1;

assign decipher_0_iibox_address137 = zext_ln708_41_fu_5205_p1;

assign decipher_0_iibox_address138 = zext_ln708_40_fu_5200_p1;

assign decipher_0_iibox_address139 = zext_ln708_39_fu_5195_p1;

assign decipher_0_iibox_address14 = zext_ln708_292_fu_14676_p1;

assign decipher_0_iibox_address140 = zext_ln708_38_fu_5190_p1;

assign decipher_0_iibox_address141 = zext_ln708_37_fu_5185_p1;

assign decipher_0_iibox_address142 = zext_ln708_36_fu_5180_p1;

assign decipher_0_iibox_address143 = zext_ln708_35_fu_5175_p1;

assign decipher_0_iibox_address144 = zext_ln708_18_fu_4063_p1;

assign decipher_0_iibox_address145 = zext_ln708_17_fu_4048_p1;

assign decipher_0_iibox_address146 = zext_ln708_16_fu_4033_p1;

assign decipher_0_iibox_address147 = zext_ln708_15_fu_4018_p1;

assign decipher_0_iibox_address148 = zext_ln708_14_fu_4003_p1;

assign decipher_0_iibox_address149 = zext_ln708_13_fu_3988_p1;

assign decipher_0_iibox_address15 = zext_ln708_291_fu_14671_p1;

assign decipher_0_iibox_address150 = zext_ln708_12_fu_3973_p1;

assign decipher_0_iibox_address151 = zext_ln708_11_fu_3958_p1;

assign decipher_0_iibox_address152 = zext_ln708_10_fu_3943_p1;

assign decipher_0_iibox_address153 = zext_ln708_9_fu_3928_p1;

assign decipher_0_iibox_address154 = zext_ln708_8_fu_3913_p1;

assign decipher_0_iibox_address155 = zext_ln708_7_fu_3898_p1;

assign decipher_0_iibox_address156 = zext_ln708_6_fu_3883_p1;

assign decipher_0_iibox_address157 = zext_ln708_5_fu_3868_p1;

assign decipher_0_iibox_address158 = zext_ln708_4_fu_3853_p1;

assign decipher_0_iibox_address159 = zext_ln708_fu_3838_p1;

assign decipher_0_iibox_address16 = zext_ln708_274_fu_13559_p1;

assign decipher_0_iibox_address17 = zext_ln708_273_fu_13554_p1;

assign decipher_0_iibox_address18 = zext_ln708_272_fu_13549_p1;

assign decipher_0_iibox_address19 = zext_ln708_271_fu_13544_p1;

assign decipher_0_iibox_address2 = zext_ln708_304_fu_14736_p1;

assign decipher_0_iibox_address20 = zext_ln708_270_fu_13539_p1;

assign decipher_0_iibox_address21 = zext_ln708_269_fu_13534_p1;

assign decipher_0_iibox_address22 = zext_ln708_268_fu_13529_p1;

assign decipher_0_iibox_address23 = zext_ln708_267_fu_13524_p1;

assign decipher_0_iibox_address24 = zext_ln708_266_fu_13519_p1;

assign decipher_0_iibox_address25 = zext_ln708_265_fu_13514_p1;

assign decipher_0_iibox_address26 = zext_ln708_264_fu_13509_p1;

assign decipher_0_iibox_address27 = zext_ln708_263_fu_13504_p1;

assign decipher_0_iibox_address28 = zext_ln708_262_fu_13499_p1;

assign decipher_0_iibox_address29 = zext_ln708_261_fu_13494_p1;

assign decipher_0_iibox_address3 = zext_ln708_303_fu_14731_p1;

assign decipher_0_iibox_address30 = zext_ln708_260_fu_13489_p1;

assign decipher_0_iibox_address31 = zext_ln708_259_fu_13484_p1;

assign decipher_0_iibox_address32 = zext_ln708_242_fu_12372_p1;

assign decipher_0_iibox_address33 = zext_ln708_241_fu_12367_p1;

assign decipher_0_iibox_address34 = zext_ln708_240_fu_12362_p1;

assign decipher_0_iibox_address35 = zext_ln708_239_fu_12357_p1;

assign decipher_0_iibox_address36 = zext_ln708_238_fu_12352_p1;

assign decipher_0_iibox_address37 = zext_ln708_237_fu_12347_p1;

assign decipher_0_iibox_address38 = zext_ln708_236_fu_12342_p1;

assign decipher_0_iibox_address39 = zext_ln708_235_fu_12337_p1;

assign decipher_0_iibox_address4 = zext_ln708_302_fu_14726_p1;

assign decipher_0_iibox_address40 = zext_ln708_234_fu_12332_p1;

assign decipher_0_iibox_address41 = zext_ln708_233_fu_12327_p1;

assign decipher_0_iibox_address42 = zext_ln708_232_fu_12322_p1;

assign decipher_0_iibox_address43 = zext_ln708_231_fu_12317_p1;

assign decipher_0_iibox_address44 = zext_ln708_230_fu_12312_p1;

assign decipher_0_iibox_address45 = zext_ln708_229_fu_12307_p1;

assign decipher_0_iibox_address46 = zext_ln708_228_fu_12302_p1;

assign decipher_0_iibox_address47 = zext_ln708_227_fu_12297_p1;

assign decipher_0_iibox_address48 = zext_ln708_210_fu_11185_p1;

assign decipher_0_iibox_address49 = zext_ln708_209_fu_11180_p1;

assign decipher_0_iibox_address5 = zext_ln708_301_fu_14721_p1;

assign decipher_0_iibox_address50 = zext_ln708_208_fu_11175_p1;

assign decipher_0_iibox_address51 = zext_ln708_207_fu_11170_p1;

assign decipher_0_iibox_address52 = zext_ln708_206_fu_11165_p1;

assign decipher_0_iibox_address53 = zext_ln708_205_fu_11160_p1;

assign decipher_0_iibox_address54 = zext_ln708_204_fu_11155_p1;

assign decipher_0_iibox_address55 = zext_ln708_203_fu_11150_p1;

assign decipher_0_iibox_address56 = zext_ln708_202_fu_11145_p1;

assign decipher_0_iibox_address57 = zext_ln708_201_fu_11140_p1;

assign decipher_0_iibox_address58 = zext_ln708_200_fu_11135_p1;

assign decipher_0_iibox_address59 = zext_ln708_199_fu_11130_p1;

assign decipher_0_iibox_address6 = zext_ln708_300_fu_14716_p1;

assign decipher_0_iibox_address60 = zext_ln708_198_fu_11125_p1;

assign decipher_0_iibox_address61 = zext_ln708_197_fu_11120_p1;

assign decipher_0_iibox_address62 = zext_ln708_196_fu_11115_p1;

assign decipher_0_iibox_address63 = zext_ln708_195_fu_11110_p1;

assign decipher_0_iibox_address64 = zext_ln708_178_fu_9998_p1;

assign decipher_0_iibox_address65 = zext_ln708_177_fu_9993_p1;

assign decipher_0_iibox_address66 = zext_ln708_176_fu_9988_p1;

assign decipher_0_iibox_address67 = zext_ln708_175_fu_9983_p1;

assign decipher_0_iibox_address68 = zext_ln708_174_fu_9978_p1;

assign decipher_0_iibox_address69 = zext_ln708_173_fu_9973_p1;

assign decipher_0_iibox_address7 = zext_ln708_299_fu_14711_p1;

assign decipher_0_iibox_address70 = zext_ln708_172_fu_9968_p1;

assign decipher_0_iibox_address71 = zext_ln708_171_fu_9963_p1;

assign decipher_0_iibox_address72 = zext_ln708_170_fu_9958_p1;

assign decipher_0_iibox_address73 = zext_ln708_169_fu_9953_p1;

assign decipher_0_iibox_address74 = zext_ln708_168_fu_9948_p1;

assign decipher_0_iibox_address75 = zext_ln708_167_fu_9943_p1;

assign decipher_0_iibox_address76 = zext_ln708_166_fu_9938_p1;

assign decipher_0_iibox_address77 = zext_ln708_165_fu_9933_p1;

assign decipher_0_iibox_address78 = zext_ln708_164_fu_9928_p1;

assign decipher_0_iibox_address79 = zext_ln708_163_fu_9923_p1;

assign decipher_0_iibox_address8 = zext_ln708_298_fu_14706_p1;

assign decipher_0_iibox_address80 = zext_ln708_146_fu_8811_p1;

assign decipher_0_iibox_address81 = zext_ln708_145_fu_8806_p1;

assign decipher_0_iibox_address82 = zext_ln708_144_fu_8801_p1;

assign decipher_0_iibox_address83 = zext_ln708_143_fu_8796_p1;

assign decipher_0_iibox_address84 = zext_ln708_142_fu_8791_p1;

assign decipher_0_iibox_address85 = zext_ln708_141_fu_8786_p1;

assign decipher_0_iibox_address86 = zext_ln708_140_fu_8781_p1;

assign decipher_0_iibox_address87 = zext_ln708_139_fu_8776_p1;

assign decipher_0_iibox_address88 = zext_ln708_138_fu_8771_p1;

assign decipher_0_iibox_address89 = zext_ln708_137_fu_8766_p1;

assign decipher_0_iibox_address9 = zext_ln708_297_fu_14701_p1;

assign decipher_0_iibox_address90 = zext_ln708_136_fu_8761_p1;

assign decipher_0_iibox_address91 = zext_ln708_135_fu_8756_p1;

assign decipher_0_iibox_address92 = zext_ln708_134_fu_8751_p1;

assign decipher_0_iibox_address93 = zext_ln708_133_fu_8746_p1;

assign decipher_0_iibox_address94 = zext_ln708_132_fu_8741_p1;

assign decipher_0_iibox_address95 = zext_ln708_131_fu_8736_p1;

assign decipher_0_iibox_address96 = zext_ln708_114_fu_7624_p1;

assign decipher_0_iibox_address97 = zext_ln708_113_fu_7619_p1;

assign decipher_0_iibox_address98 = zext_ln708_112_fu_7614_p1;

assign decipher_0_iibox_address99 = zext_ln708_111_fu_7609_p1;

assign p_Result_10_fu_14751_p17 = {{{{{{{{{{{{{{{{decipher_0_iibox_q0}, {decipher_0_iibox_q1}}, {decipher_0_iibox_q2}}, {decipher_0_iibox_q3}}, {decipher_0_iibox_q4}}, {decipher_0_iibox_q5}}, {decipher_0_iibox_q6}}, {decipher_0_iibox_q7}}, {decipher_0_iibox_q8}}, {decipher_0_iibox_q9}}, {decipher_0_iibox_q10}}, {decipher_0_iibox_q11}}, {decipher_0_iibox_q12}}, {decipher_0_iibox_q13}}, {decipher_0_iibox_q14}}, {decipher_0_iibox_q15}};

assign p_Result_2_fu_5255_p17 = {{{{{{{{{{{{{{{{decipher_0_iibox_q128}, {decipher_0_iibox_q129}}, {decipher_0_iibox_q130}}, {decipher_0_iibox_q131}}, {decipher_0_iibox_q132}}, {decipher_0_iibox_q133}}, {decipher_0_iibox_q134}}, {decipher_0_iibox_q135}}, {decipher_0_iibox_q136}}, {decipher_0_iibox_q137}}, {decipher_0_iibox_q138}}, {decipher_0_iibox_q139}}, {decipher_0_iibox_q140}}, {decipher_0_iibox_q141}}, {decipher_0_iibox_q142}}, {decipher_0_iibox_q143}};

assign p_Result_3_fu_6442_p17 = {{{{{{{{{{{{{{{{decipher_0_iibox_q112}, {decipher_0_iibox_q113}}, {decipher_0_iibox_q114}}, {decipher_0_iibox_q115}}, {decipher_0_iibox_q116}}, {decipher_0_iibox_q117}}, {decipher_0_iibox_q118}}, {decipher_0_iibox_q119}}, {decipher_0_iibox_q120}}, {decipher_0_iibox_q121}}, {decipher_0_iibox_q122}}, {decipher_0_iibox_q123}}, {decipher_0_iibox_q124}}, {decipher_0_iibox_q125}}, {decipher_0_iibox_q126}}, {decipher_0_iibox_q127}};

assign p_Result_4_fu_7629_p17 = {{{{{{{{{{{{{{{{decipher_0_iibox_q96}, {decipher_0_iibox_q97}}, {decipher_0_iibox_q98}}, {decipher_0_iibox_q99}}, {decipher_0_iibox_q100}}, {decipher_0_iibox_q101}}, {decipher_0_iibox_q102}}, {decipher_0_iibox_q103}}, {decipher_0_iibox_q104}}, {decipher_0_iibox_q105}}, {decipher_0_iibox_q106}}, {decipher_0_iibox_q107}}, {decipher_0_iibox_q108}}, {decipher_0_iibox_q109}}, {decipher_0_iibox_q110}}, {decipher_0_iibox_q111}};

assign p_Result_5_fu_8816_p17 = {{{{{{{{{{{{{{{{decipher_0_iibox_q80}, {decipher_0_iibox_q81}}, {decipher_0_iibox_q82}}, {decipher_0_iibox_q83}}, {decipher_0_iibox_q84}}, {decipher_0_iibox_q85}}, {decipher_0_iibox_q86}}, {decipher_0_iibox_q87}}, {decipher_0_iibox_q88}}, {decipher_0_iibox_q89}}, {decipher_0_iibox_q90}}, {decipher_0_iibox_q91}}, {decipher_0_iibox_q92}}, {decipher_0_iibox_q93}}, {decipher_0_iibox_q94}}, {decipher_0_iibox_q95}};

assign p_Result_6_fu_10003_p17 = {{{{{{{{{{{{{{{{decipher_0_iibox_q64}, {decipher_0_iibox_q65}}, {decipher_0_iibox_q66}}, {decipher_0_iibox_q67}}, {decipher_0_iibox_q68}}, {decipher_0_iibox_q69}}, {decipher_0_iibox_q70}}, {decipher_0_iibox_q71}}, {decipher_0_iibox_q72}}, {decipher_0_iibox_q73}}, {decipher_0_iibox_q74}}, {decipher_0_iibox_q75}}, {decipher_0_iibox_q76}}, {decipher_0_iibox_q77}}, {decipher_0_iibox_q78}}, {decipher_0_iibox_q79}};

assign p_Result_7_fu_11190_p17 = {{{{{{{{{{{{{{{{decipher_0_iibox_q48}, {decipher_0_iibox_q49}}, {decipher_0_iibox_q50}}, {decipher_0_iibox_q51}}, {decipher_0_iibox_q52}}, {decipher_0_iibox_q53}}, {decipher_0_iibox_q54}}, {decipher_0_iibox_q55}}, {decipher_0_iibox_q56}}, {decipher_0_iibox_q57}}, {decipher_0_iibox_q58}}, {decipher_0_iibox_q59}}, {decipher_0_iibox_q60}}, {decipher_0_iibox_q61}}, {decipher_0_iibox_q62}}, {decipher_0_iibox_q63}};

assign p_Result_8_fu_12377_p17 = {{{{{{{{{{{{{{{{decipher_0_iibox_q32}, {decipher_0_iibox_q33}}, {decipher_0_iibox_q34}}, {decipher_0_iibox_q35}}, {decipher_0_iibox_q36}}, {decipher_0_iibox_q37}}, {decipher_0_iibox_q38}}, {decipher_0_iibox_q39}}, {decipher_0_iibox_q40}}, {decipher_0_iibox_q41}}, {decipher_0_iibox_q42}}, {decipher_0_iibox_q43}}, {decipher_0_iibox_q44}}, {decipher_0_iibox_q45}}, {decipher_0_iibox_q46}}, {decipher_0_iibox_q47}};

assign p_Result_9_fu_13564_p17 = {{{{{{{{{{{{{{{{decipher_0_iibox_q16}, {decipher_0_iibox_q17}}, {decipher_0_iibox_q18}}, {decipher_0_iibox_q19}}, {decipher_0_iibox_q20}}, {decipher_0_iibox_q21}}, {decipher_0_iibox_q22}}, {decipher_0_iibox_q23}}, {decipher_0_iibox_q24}}, {decipher_0_iibox_q25}}, {decipher_0_iibox_q26}}, {decipher_0_iibox_q27}}, {decipher_0_iibox_q28}}, {decipher_0_iibox_q29}}, {decipher_0_iibox_q30}}, {decipher_0_iibox_q31}};

assign p_Result_s_fu_4068_p17 = {{{{{{{{{{{{{{{{decipher_0_iibox_q144}, {decipher_0_iibox_q145}}, {decipher_0_iibox_q146}}, {decipher_0_iibox_q147}}, {decipher_0_iibox_q148}}, {decipher_0_iibox_q149}}, {decipher_0_iibox_q150}}, {decipher_0_iibox_q151}}, {decipher_0_iibox_q152}}, {decipher_0_iibox_q153}}, {decipher_0_iibox_q154}}, {decipher_0_iibox_q155}}, {decipher_0_iibox_q156}}, {decipher_0_iibox_q157}}, {decipher_0_iibox_q158}}, {decipher_0_iibox_q159}};

assign ret_V_fu_3828_p2 = (p_read10 ^ ciphertext);

assign state_V_20_fu_4104_p2 = (p_read_2_reg_14792 ^ p_Result_s_fu_4068_p17);

assign state_V_21_fu_5291_p2 = (p_read_3_reg_14797_pp0_iter2_reg ^ p_Result_2_fu_5255_p17);

assign state_V_22_fu_6478_p2 = (p_read_4_reg_14802_pp0_iter4_reg ^ p_Result_3_fu_6442_p17);

assign state_V_23_fu_7665_p2 = (p_read_5_reg_14807_pp0_iter6_reg ^ p_Result_4_fu_7629_p17);

assign state_V_24_fu_8852_p2 = (p_read_6_reg_14812_pp0_iter8_reg ^ p_Result_5_fu_8816_p17);

assign state_V_25_fu_10039_p2 = (p_read_7_reg_14817_pp0_iter10_reg ^ p_Result_6_fu_10003_p17);

assign state_V_26_fu_12413_p2 = (p_read_9_reg_14827_pp0_iter14_reg ^ p_Result_8_fu_12377_p17);

assign state_V_27_fu_13600_p2 = (p_read_10_reg_14832_pp0_iter16_reg ^ p_Result_9_fu_13564_p17);

assign state_V_fu_11226_p2 = (p_read_8_reg_14822_pp0_iter12_reg ^ p_Result_7_fu_11190_p17);

assign tmp_100_fu_5724_p4 = {{decipher_0_i32box_q122[31:24]}};

assign tmp_101_fu_5380_p4 = {{state_V_21_fu_5291_p2[55:48]}};

assign tmp_102_fu_5738_p4 = {{decipher_0_i32box_q121[15:8]}};

assign tmp_103_fu_5748_p4 = {{decipher_0_i32box_q121[23:16]}};

assign tmp_104_fu_5758_p4 = {{decipher_0_i32box_q121[31:24]}};

assign tmp_105_fu_5395_p4 = {{state_V_21_fu_5291_p2[63:56]}};

assign tmp_106_fu_5772_p4 = {{decipher_0_i32box_q120[15:8]}};

assign tmp_107_fu_5782_p4 = {{decipher_0_i32box_q120[23:16]}};

assign tmp_108_fu_5792_p4 = {{decipher_0_i32box_q120[31:24]}};

assign tmp_109_fu_5410_p4 = {{state_V_21_fu_5291_p2[71:64]}};

assign tmp_10_fu_3993_p4 = {{ret_V_fu_3828_p2[127:120]}};

assign tmp_110_fu_5806_p4 = {{decipher_0_i32box_q119[15:8]}};

assign tmp_111_fu_5816_p4 = {{decipher_0_i32box_q119[23:16]}};

assign tmp_112_fu_5826_p4 = {{decipher_0_i32box_q119[31:24]}};

assign tmp_113_fu_5425_p4 = {{state_V_21_fu_5291_p2[79:72]}};

assign tmp_114_fu_5840_p4 = {{decipher_0_i32box_q118[15:8]}};

assign tmp_115_fu_5850_p4 = {{decipher_0_i32box_q118[23:16]}};

assign tmp_116_fu_5860_p4 = {{decipher_0_i32box_q118[31:24]}};

assign tmp_117_fu_5440_p4 = {{state_V_21_fu_5291_p2[87:80]}};

assign tmp_118_fu_5874_p4 = {{decipher_0_i32box_q117[15:8]}};

assign tmp_119_fu_5884_p4 = {{decipher_0_i32box_q117[23:16]}};

assign tmp_11_fu_4008_p4 = {{ret_V_fu_3828_p2[103:96]}};

assign tmp_120_fu_5894_p4 = {{decipher_0_i32box_q117[31:24]}};

assign tmp_121_fu_5455_p4 = {{state_V_21_fu_5291_p2[95:88]}};

assign tmp_122_fu_5908_p4 = {{decipher_0_i32box_q116[15:8]}};

assign tmp_123_fu_5918_p4 = {{decipher_0_i32box_q116[23:16]}};

assign tmp_124_fu_5928_p4 = {{decipher_0_i32box_q116[31:24]}};

assign tmp_125_fu_5470_p4 = {{state_V_21_fu_5291_p2[103:96]}};

assign tmp_126_fu_5942_p4 = {{decipher_0_i32box_q115[15:8]}};

assign tmp_127_fu_5952_p4 = {{decipher_0_i32box_q115[23:16]}};

assign tmp_128_fu_5962_p4 = {{decipher_0_i32box_q115[31:24]}};

assign tmp_129_fu_5485_p4 = {{state_V_21_fu_5291_p2[111:104]}};

assign tmp_12_fu_4023_p4 = {{ret_V_fu_3828_p2[79:72]}};

assign tmp_130_fu_5976_p4 = {{decipher_0_i32box_q114[15:8]}};

assign tmp_131_fu_5986_p4 = {{decipher_0_i32box_q114[23:16]}};

assign tmp_132_fu_5996_p4 = {{decipher_0_i32box_q114[31:24]}};

assign tmp_133_fu_5500_p4 = {{state_V_21_fu_5291_p2[119:112]}};

assign tmp_134_fu_6010_p4 = {{decipher_0_i32box_q113[15:8]}};

assign tmp_135_fu_6020_p4 = {{decipher_0_i32box_q113[23:16]}};

assign tmp_136_fu_6030_p4 = {{decipher_0_i32box_q113[31:24]}};

assign tmp_137_fu_5515_p4 = {{state_V_21_fu_5291_p2[127:120]}};

assign tmp_138_fu_6044_p4 = {{decipher_0_i32box_q112[15:8]}};

assign tmp_139_fu_6054_p4 = {{decipher_0_i32box_q112[23:16]}};

assign tmp_13_fu_4038_p4 = {{ret_V_fu_3828_p2[55:48]}};

assign tmp_140_fu_6064_p4 = {{decipher_0_i32box_q112[31:24]}};

assign tmp_141_fu_6721_p4 = {{decipher_0_i32box_q111[15:8]}};

assign tmp_142_fu_6731_p4 = {{decipher_0_i32box_q111[23:16]}};

assign tmp_143_fu_6741_p4 = {{decipher_0_i32box_q111[31:24]}};

assign tmp_144_fu_6492_p4 = {{state_V_22_fu_6478_p2[15:8]}};

assign tmp_145_fu_6755_p4 = {{decipher_0_i32box_q110[15:8]}};

assign tmp_146_fu_6765_p4 = {{decipher_0_i32box_q110[23:16]}};

assign tmp_147_fu_6775_p4 = {{decipher_0_i32box_q110[31:24]}};

assign tmp_148_fu_6507_p4 = {{state_V_22_fu_6478_p2[23:16]}};

assign tmp_149_fu_6789_p4 = {{decipher_0_i32box_q109[15:8]}};

assign tmp_14_fu_4053_p4 = {{ret_V_fu_3828_p2[31:24]}};

assign tmp_150_fu_6799_p4 = {{decipher_0_i32box_q109[23:16]}};

assign tmp_151_fu_6809_p4 = {{decipher_0_i32box_q109[31:24]}};

assign tmp_152_fu_6522_p4 = {{state_V_22_fu_6478_p2[31:24]}};

assign tmp_153_fu_6823_p4 = {{decipher_0_i32box_q108[15:8]}};

assign tmp_154_fu_6833_p4 = {{decipher_0_i32box_q108[23:16]}};

assign tmp_155_fu_6843_p4 = {{decipher_0_i32box_q108[31:24]}};

assign tmp_156_fu_6537_p4 = {{state_V_22_fu_6478_p2[39:32]}};

assign tmp_157_fu_6857_p4 = {{decipher_0_i32box_q107[15:8]}};

assign tmp_158_fu_6867_p4 = {{decipher_0_i32box_q107[23:16]}};

assign tmp_159_fu_6877_p4 = {{decipher_0_i32box_q107[31:24]}};

assign tmp_15_fu_4347_p4 = {{decipher_0_i32box_q143[15:8]}};

assign tmp_160_fu_6552_p4 = {{state_V_22_fu_6478_p2[47:40]}};

assign tmp_161_fu_6891_p4 = {{decipher_0_i32box_q106[15:8]}};

assign tmp_162_fu_6901_p4 = {{decipher_0_i32box_q106[23:16]}};

assign tmp_163_fu_6911_p4 = {{decipher_0_i32box_q106[31:24]}};

assign tmp_164_fu_6567_p4 = {{state_V_22_fu_6478_p2[55:48]}};

assign tmp_165_fu_6925_p4 = {{decipher_0_i32box_q105[15:8]}};

assign tmp_166_fu_6935_p4 = {{decipher_0_i32box_q105[23:16]}};

assign tmp_167_fu_6945_p4 = {{decipher_0_i32box_q105[31:24]}};

assign tmp_168_fu_6582_p4 = {{state_V_22_fu_6478_p2[63:56]}};

assign tmp_169_fu_6959_p4 = {{decipher_0_i32box_q104[15:8]}};

assign tmp_16_fu_4357_p4 = {{decipher_0_i32box_q143[23:16]}};

assign tmp_170_fu_6969_p4 = {{decipher_0_i32box_q104[23:16]}};

assign tmp_171_fu_6979_p4 = {{decipher_0_i32box_q104[31:24]}};

assign tmp_172_fu_6597_p4 = {{state_V_22_fu_6478_p2[71:64]}};

assign tmp_173_fu_6993_p4 = {{decipher_0_i32box_q103[15:8]}};

assign tmp_174_fu_7003_p4 = {{decipher_0_i32box_q103[23:16]}};

assign tmp_175_fu_7013_p4 = {{decipher_0_i32box_q103[31:24]}};

assign tmp_176_fu_6612_p4 = {{state_V_22_fu_6478_p2[79:72]}};

assign tmp_177_fu_7027_p4 = {{decipher_0_i32box_q102[15:8]}};

assign tmp_178_fu_7037_p4 = {{decipher_0_i32box_q102[23:16]}};

assign tmp_179_fu_7047_p4 = {{decipher_0_i32box_q102[31:24]}};

assign tmp_17_fu_4367_p4 = {{decipher_0_i32box_q143[31:24]}};

assign tmp_180_fu_6627_p4 = {{state_V_22_fu_6478_p2[87:80]}};

assign tmp_181_fu_7061_p4 = {{decipher_0_i32box_q101[15:8]}};

assign tmp_182_fu_7071_p4 = {{decipher_0_i32box_q101[23:16]}};

assign tmp_183_fu_7081_p4 = {{decipher_0_i32box_q101[31:24]}};

assign tmp_184_fu_6642_p4 = {{state_V_22_fu_6478_p2[95:88]}};

assign tmp_185_fu_7095_p4 = {{decipher_0_i32box_q100[15:8]}};

assign tmp_186_fu_7105_p4 = {{decipher_0_i32box_q100[23:16]}};

assign tmp_187_fu_7115_p4 = {{decipher_0_i32box_q100[31:24]}};

assign tmp_188_fu_6657_p4 = {{state_V_22_fu_6478_p2[103:96]}};

assign tmp_189_fu_7129_p4 = {{decipher_0_i32box_q99[15:8]}};

assign tmp_18_fu_4118_p4 = {{state_V_20_fu_4104_p2[15:8]}};

assign tmp_190_fu_7139_p4 = {{decipher_0_i32box_q99[23:16]}};

assign tmp_191_fu_7149_p4 = {{decipher_0_i32box_q99[31:24]}};

assign tmp_192_fu_6672_p4 = {{state_V_22_fu_6478_p2[111:104]}};

assign tmp_193_fu_7163_p4 = {{decipher_0_i32box_q98[15:8]}};

assign tmp_194_fu_7173_p4 = {{decipher_0_i32box_q98[23:16]}};

assign tmp_195_fu_7183_p4 = {{decipher_0_i32box_q98[31:24]}};

assign tmp_196_fu_6687_p4 = {{state_V_22_fu_6478_p2[119:112]}};

assign tmp_197_fu_7197_p4 = {{decipher_0_i32box_q97[15:8]}};

assign tmp_198_fu_7207_p4 = {{decipher_0_i32box_q97[23:16]}};

assign tmp_199_fu_7217_p4 = {{decipher_0_i32box_q97[31:24]}};

assign tmp_19_fu_4381_p4 = {{decipher_0_i32box_q142[15:8]}};

assign tmp_1_V_1_fu_6320_p2 = (xor_ln1545_92_fu_6314_p2 ^ xor_ln1545_91_fu_6308_p2);

assign tmp_1_V_2_fu_7507_p2 = (xor_ln1545_140_fu_7501_p2 ^ xor_ln1545_139_fu_7495_p2);

assign tmp_1_V_3_fu_8694_p2 = (xor_ln1545_188_fu_8688_p2 ^ xor_ln1545_187_fu_8682_p2);

assign tmp_1_V_4_fu_9881_p2 = (xor_ln1545_236_fu_9875_p2 ^ xor_ln1545_235_fu_9869_p2);

assign tmp_1_V_5_fu_11068_p2 = (xor_ln1545_284_fu_11062_p2 ^ xor_ln1545_283_fu_11056_p2);

assign tmp_1_V_6_fu_12255_p2 = (xor_ln1545_332_fu_12249_p2 ^ xor_ln1545_331_fu_12243_p2);

assign tmp_1_V_7_fu_13442_p2 = (xor_ln1545_380_fu_13436_p2 ^ xor_ln1545_379_fu_13430_p2);

assign tmp_1_V_8_fu_14629_p2 = (xor_ln1545_428_fu_14623_p2 ^ xor_ln1545_427_fu_14617_p2);

assign tmp_1_V_fu_5133_p2 = (xor_ln1545_44_fu_5127_p2 ^ xor_ln1545_43_fu_5121_p2);

assign tmp_1_fu_3843_p4 = {{ret_V_fu_3828_p2[111:104]}};

assign tmp_200_fu_6702_p4 = {{state_V_22_fu_6478_p2[127:120]}};

assign tmp_201_fu_7231_p4 = {{decipher_0_i32box_q96[15:8]}};

assign tmp_202_fu_7241_p4 = {{decipher_0_i32box_q96[23:16]}};

assign tmp_203_fu_7251_p4 = {{decipher_0_i32box_q96[31:24]}};

assign tmp_204_fu_7908_p4 = {{decipher_0_i32box_q95[15:8]}};

assign tmp_205_fu_7918_p4 = {{decipher_0_i32box_q95[23:16]}};

assign tmp_206_fu_7928_p4 = {{decipher_0_i32box_q95[31:24]}};

assign tmp_207_fu_7679_p4 = {{state_V_23_fu_7665_p2[15:8]}};

assign tmp_208_fu_7942_p4 = {{decipher_0_i32box_q94[15:8]}};

assign tmp_209_fu_7952_p4 = {{decipher_0_i32box_q94[23:16]}};

assign tmp_20_fu_4391_p4 = {{decipher_0_i32box_q142[23:16]}};

assign tmp_210_fu_7962_p4 = {{decipher_0_i32box_q94[31:24]}};

assign tmp_211_fu_7694_p4 = {{state_V_23_fu_7665_p2[23:16]}};

assign tmp_212_fu_7976_p4 = {{decipher_0_i32box_q93[15:8]}};

assign tmp_213_fu_7986_p4 = {{decipher_0_i32box_q93[23:16]}};

assign tmp_214_fu_7996_p4 = {{decipher_0_i32box_q93[31:24]}};

assign tmp_215_fu_7709_p4 = {{state_V_23_fu_7665_p2[31:24]}};

assign tmp_216_fu_8010_p4 = {{decipher_0_i32box_q92[15:8]}};

assign tmp_217_fu_8020_p4 = {{decipher_0_i32box_q92[23:16]}};

assign tmp_218_fu_8030_p4 = {{decipher_0_i32box_q92[31:24]}};

assign tmp_219_fu_7724_p4 = {{state_V_23_fu_7665_p2[39:32]}};

assign tmp_21_fu_4401_p4 = {{decipher_0_i32box_q142[31:24]}};

assign tmp_220_fu_8044_p4 = {{decipher_0_i32box_q91[15:8]}};

assign tmp_221_fu_8054_p4 = {{decipher_0_i32box_q91[23:16]}};

assign tmp_222_fu_8064_p4 = {{decipher_0_i32box_q91[31:24]}};

assign tmp_223_fu_7739_p4 = {{state_V_23_fu_7665_p2[47:40]}};

assign tmp_224_fu_8078_p4 = {{decipher_0_i32box_q90[15:8]}};

assign tmp_225_fu_8088_p4 = {{decipher_0_i32box_q90[23:16]}};

assign tmp_226_fu_8098_p4 = {{decipher_0_i32box_q90[31:24]}};

assign tmp_227_fu_7754_p4 = {{state_V_23_fu_7665_p2[55:48]}};

assign tmp_228_fu_8112_p4 = {{decipher_0_i32box_q89[15:8]}};

assign tmp_229_fu_8122_p4 = {{decipher_0_i32box_q89[23:16]}};

assign tmp_22_fu_4133_p4 = {{state_V_20_fu_4104_p2[23:16]}};

assign tmp_230_fu_8132_p4 = {{decipher_0_i32box_q89[31:24]}};

assign tmp_231_fu_7769_p4 = {{state_V_23_fu_7665_p2[63:56]}};

assign tmp_232_fu_8146_p4 = {{decipher_0_i32box_q88[15:8]}};

assign tmp_233_fu_8156_p4 = {{decipher_0_i32box_q88[23:16]}};

assign tmp_234_fu_8166_p4 = {{decipher_0_i32box_q88[31:24]}};

assign tmp_235_fu_7784_p4 = {{state_V_23_fu_7665_p2[71:64]}};

assign tmp_236_fu_8180_p4 = {{decipher_0_i32box_q87[15:8]}};

assign tmp_237_fu_8190_p4 = {{decipher_0_i32box_q87[23:16]}};

assign tmp_238_fu_8200_p4 = {{decipher_0_i32box_q87[31:24]}};

assign tmp_239_fu_7799_p4 = {{state_V_23_fu_7665_p2[79:72]}};

assign tmp_23_fu_4415_p4 = {{decipher_0_i32box_q141[15:8]}};

assign tmp_240_fu_8214_p4 = {{decipher_0_i32box_q86[15:8]}};

assign tmp_241_fu_8224_p4 = {{decipher_0_i32box_q86[23:16]}};

assign tmp_242_fu_8234_p4 = {{decipher_0_i32box_q86[31:24]}};

assign tmp_243_fu_7814_p4 = {{state_V_23_fu_7665_p2[87:80]}};

assign tmp_244_fu_8248_p4 = {{decipher_0_i32box_q85[15:8]}};

assign tmp_245_fu_8258_p4 = {{decipher_0_i32box_q85[23:16]}};

assign tmp_246_fu_8268_p4 = {{decipher_0_i32box_q85[31:24]}};

assign tmp_247_fu_7829_p4 = {{state_V_23_fu_7665_p2[95:88]}};

assign tmp_248_fu_8282_p4 = {{decipher_0_i32box_q84[15:8]}};

assign tmp_249_fu_8292_p4 = {{decipher_0_i32box_q84[23:16]}};

assign tmp_24_fu_4425_p4 = {{decipher_0_i32box_q141[23:16]}};

assign tmp_250_fu_8302_p4 = {{decipher_0_i32box_q84[31:24]}};

assign tmp_251_fu_7844_p4 = {{state_V_23_fu_7665_p2[103:96]}};

assign tmp_252_fu_8316_p4 = {{decipher_0_i32box_q83[15:8]}};

assign tmp_253_fu_8326_p4 = {{decipher_0_i32box_q83[23:16]}};

assign tmp_254_fu_8336_p4 = {{decipher_0_i32box_q83[31:24]}};

assign tmp_255_fu_7859_p4 = {{state_V_23_fu_7665_p2[111:104]}};

assign tmp_256_fu_8350_p4 = {{decipher_0_i32box_q82[15:8]}};

assign tmp_257_fu_8360_p4 = {{decipher_0_i32box_q82[23:16]}};

assign tmp_258_fu_8370_p4 = {{decipher_0_i32box_q82[31:24]}};

assign tmp_259_fu_7874_p4 = {{state_V_23_fu_7665_p2[119:112]}};

assign tmp_25_fu_4435_p4 = {{decipher_0_i32box_q141[31:24]}};

assign tmp_260_fu_8384_p4 = {{decipher_0_i32box_q81[15:8]}};

assign tmp_261_fu_8394_p4 = {{decipher_0_i32box_q81[23:16]}};

assign tmp_262_fu_8404_p4 = {{decipher_0_i32box_q81[31:24]}};

assign tmp_263_fu_7889_p4 = {{state_V_23_fu_7665_p2[127:120]}};

assign tmp_264_fu_8418_p4 = {{decipher_0_i32box_q80[15:8]}};

assign tmp_265_fu_8428_p4 = {{decipher_0_i32box_q80[23:16]}};

assign tmp_266_fu_8438_p4 = {{decipher_0_i32box_q80[31:24]}};

assign tmp_267_fu_9095_p4 = {{decipher_0_i32box_q79[15:8]}};

assign tmp_268_fu_9105_p4 = {{decipher_0_i32box_q79[23:16]}};

assign tmp_269_fu_9115_p4 = {{decipher_0_i32box_q79[31:24]}};

assign tmp_26_fu_4148_p4 = {{state_V_20_fu_4104_p2[31:24]}};

assign tmp_270_fu_8866_p4 = {{state_V_24_fu_8852_p2[15:8]}};

assign tmp_271_fu_9129_p4 = {{decipher_0_i32box_q78[15:8]}};

assign tmp_272_fu_9139_p4 = {{decipher_0_i32box_q78[23:16]}};

assign tmp_273_fu_9149_p4 = {{decipher_0_i32box_q78[31:24]}};

assign tmp_274_fu_8881_p4 = {{state_V_24_fu_8852_p2[23:16]}};

assign tmp_275_fu_9163_p4 = {{decipher_0_i32box_q77[15:8]}};

assign tmp_276_fu_9173_p4 = {{decipher_0_i32box_q77[23:16]}};

assign tmp_277_fu_9183_p4 = {{decipher_0_i32box_q77[31:24]}};

assign tmp_278_fu_8896_p4 = {{state_V_24_fu_8852_p2[31:24]}};

assign tmp_279_fu_9197_p4 = {{decipher_0_i32box_q76[15:8]}};

assign tmp_27_fu_4449_p4 = {{decipher_0_i32box_q140[15:8]}};

assign tmp_280_fu_9207_p4 = {{decipher_0_i32box_q76[23:16]}};

assign tmp_281_fu_9217_p4 = {{decipher_0_i32box_q76[31:24]}};

assign tmp_282_fu_8911_p4 = {{state_V_24_fu_8852_p2[39:32]}};

assign tmp_283_fu_9231_p4 = {{decipher_0_i32box_q75[15:8]}};

assign tmp_284_fu_9241_p4 = {{decipher_0_i32box_q75[23:16]}};

assign tmp_285_fu_9251_p4 = {{decipher_0_i32box_q75[31:24]}};

assign tmp_286_fu_8926_p4 = {{state_V_24_fu_8852_p2[47:40]}};

assign tmp_287_fu_9265_p4 = {{decipher_0_i32box_q74[15:8]}};

assign tmp_288_fu_9275_p4 = {{decipher_0_i32box_q74[23:16]}};

assign tmp_289_fu_9285_p4 = {{decipher_0_i32box_q74[31:24]}};

assign tmp_28_fu_4459_p4 = {{decipher_0_i32box_q140[23:16]}};

assign tmp_290_fu_8941_p4 = {{state_V_24_fu_8852_p2[55:48]}};

assign tmp_291_fu_9299_p4 = {{decipher_0_i32box_q73[15:8]}};

assign tmp_292_fu_9309_p4 = {{decipher_0_i32box_q73[23:16]}};

assign tmp_293_fu_9319_p4 = {{decipher_0_i32box_q73[31:24]}};

assign tmp_294_fu_8956_p4 = {{state_V_24_fu_8852_p2[63:56]}};

assign tmp_295_fu_9333_p4 = {{decipher_0_i32box_q72[15:8]}};

assign tmp_296_fu_9343_p4 = {{decipher_0_i32box_q72[23:16]}};

assign tmp_297_fu_9353_p4 = {{decipher_0_i32box_q72[31:24]}};

assign tmp_298_fu_8971_p4 = {{state_V_24_fu_8852_p2[71:64]}};

assign tmp_299_fu_9367_p4 = {{decipher_0_i32box_q71[15:8]}};

assign tmp_29_fu_4469_p4 = {{decipher_0_i32box_q140[31:24]}};

assign tmp_2_1_V_1_fu_6266_p2 = (xor_ln1545_83_fu_6260_p2 ^ xor_ln1545_82_fu_6254_p2);

assign tmp_2_1_V_2_fu_7453_p2 = (xor_ln1545_131_fu_7447_p2 ^ xor_ln1545_130_fu_7441_p2);

assign tmp_2_1_V_3_fu_8640_p2 = (xor_ln1545_179_fu_8634_p2 ^ xor_ln1545_178_fu_8628_p2);

assign tmp_2_1_V_4_fu_9827_p2 = (xor_ln1545_227_fu_9821_p2 ^ xor_ln1545_226_fu_9815_p2);

assign tmp_2_1_V_5_fu_11014_p2 = (xor_ln1545_275_fu_11008_p2 ^ xor_ln1545_274_fu_11002_p2);

assign tmp_2_1_V_6_fu_12201_p2 = (xor_ln1545_323_fu_12195_p2 ^ xor_ln1545_322_fu_12189_p2);

assign tmp_2_1_V_7_fu_13388_p2 = (xor_ln1545_371_fu_13382_p2 ^ xor_ln1545_370_fu_13376_p2);

assign tmp_2_1_V_8_fu_14575_p2 = (xor_ln1545_419_fu_14569_p2 ^ xor_ln1545_418_fu_14563_p2);

assign tmp_2_1_V_fu_5079_p2 = (xor_ln1545_35_fu_5073_p2 ^ xor_ln1545_34_fu_5067_p2);

assign tmp_2_2_V_1_fu_6338_p2 = (xor_ln1545_95_fu_6332_p2 ^ xor_ln1545_94_fu_6326_p2);

assign tmp_2_2_V_2_fu_7525_p2 = (xor_ln1545_143_fu_7519_p2 ^ xor_ln1545_142_fu_7513_p2);

assign tmp_2_2_V_3_fu_8712_p2 = (xor_ln1545_191_fu_8706_p2 ^ xor_ln1545_190_fu_8700_p2);

assign tmp_2_2_V_4_fu_9899_p2 = (xor_ln1545_239_fu_9893_p2 ^ xor_ln1545_238_fu_9887_p2);

assign tmp_2_2_V_5_fu_11086_p2 = (xor_ln1545_287_fu_11080_p2 ^ xor_ln1545_286_fu_11074_p2);

assign tmp_2_2_V_6_fu_12273_p2 = (xor_ln1545_335_fu_12267_p2 ^ xor_ln1545_334_fu_12261_p2);

assign tmp_2_2_V_7_fu_13460_p2 = (xor_ln1545_383_fu_13454_p2 ^ xor_ln1545_382_fu_13448_p2);

assign tmp_2_2_V_8_fu_14647_p2 = (xor_ln1545_431_fu_14641_p2 ^ xor_ln1545_430_fu_14635_p2);

assign tmp_2_2_V_fu_5151_p2 = (xor_ln1545_47_fu_5145_p2 ^ xor_ln1545_46_fu_5139_p2);

assign tmp_2_fu_3858_p4 = {{ret_V_fu_3828_p2[87:80]}};

assign tmp_300_fu_9377_p4 = {{decipher_0_i32box_q71[23:16]}};

assign tmp_301_fu_9387_p4 = {{decipher_0_i32box_q71[31:24]}};

assign tmp_302_fu_8986_p4 = {{state_V_24_fu_8852_p2[79:72]}};

assign tmp_303_fu_9401_p4 = {{decipher_0_i32box_q70[15:8]}};

assign tmp_304_fu_9411_p4 = {{decipher_0_i32box_q70[23:16]}};

assign tmp_305_fu_9421_p4 = {{decipher_0_i32box_q70[31:24]}};

assign tmp_306_fu_9001_p4 = {{state_V_24_fu_8852_p2[87:80]}};

assign tmp_307_fu_9435_p4 = {{decipher_0_i32box_q69[15:8]}};

assign tmp_308_fu_9445_p4 = {{decipher_0_i32box_q69[23:16]}};

assign tmp_309_fu_9455_p4 = {{decipher_0_i32box_q69[31:24]}};

assign tmp_30_fu_4163_p4 = {{state_V_20_fu_4104_p2[39:32]}};

assign tmp_310_fu_9016_p4 = {{state_V_24_fu_8852_p2[95:88]}};

assign tmp_311_fu_9469_p4 = {{decipher_0_i32box_q68[15:8]}};

assign tmp_312_fu_9479_p4 = {{decipher_0_i32box_q68[23:16]}};

assign tmp_313_fu_9489_p4 = {{decipher_0_i32box_q68[31:24]}};

assign tmp_314_fu_9031_p4 = {{state_V_24_fu_8852_p2[103:96]}};

assign tmp_315_fu_9503_p4 = {{decipher_0_i32box_q67[15:8]}};

assign tmp_316_fu_9513_p4 = {{decipher_0_i32box_q67[23:16]}};

assign tmp_317_fu_9523_p4 = {{decipher_0_i32box_q67[31:24]}};

assign tmp_318_fu_9046_p4 = {{state_V_24_fu_8852_p2[111:104]}};

assign tmp_319_fu_9537_p4 = {{decipher_0_i32box_q66[15:8]}};

assign tmp_31_fu_4483_p4 = {{decipher_0_i32box_q139[15:8]}};

assign tmp_320_fu_9547_p4 = {{decipher_0_i32box_q66[23:16]}};

assign tmp_321_fu_9557_p4 = {{decipher_0_i32box_q66[31:24]}};

assign tmp_322_fu_9061_p4 = {{state_V_24_fu_8852_p2[119:112]}};

assign tmp_323_fu_9571_p4 = {{decipher_0_i32box_q65[15:8]}};

assign tmp_324_fu_9581_p4 = {{decipher_0_i32box_q65[23:16]}};

assign tmp_325_fu_9591_p4 = {{decipher_0_i32box_q65[31:24]}};

assign tmp_326_fu_9076_p4 = {{state_V_24_fu_8852_p2[127:120]}};

assign tmp_327_fu_9605_p4 = {{decipher_0_i32box_q64[15:8]}};

assign tmp_328_fu_9615_p4 = {{decipher_0_i32box_q64[23:16]}};

assign tmp_329_fu_9625_p4 = {{decipher_0_i32box_q64[31:24]}};

assign tmp_32_fu_4493_p4 = {{decipher_0_i32box_q139[23:16]}};

assign tmp_330_fu_10282_p4 = {{decipher_0_i32box_q63[15:8]}};

assign tmp_331_fu_10292_p4 = {{decipher_0_i32box_q63[23:16]}};

assign tmp_332_fu_10302_p4 = {{decipher_0_i32box_q63[31:24]}};

assign tmp_333_fu_10053_p4 = {{state_V_25_fu_10039_p2[15:8]}};

assign tmp_334_fu_10316_p4 = {{decipher_0_i32box_q62[15:8]}};

assign tmp_335_fu_10326_p4 = {{decipher_0_i32box_q62[23:16]}};

assign tmp_336_fu_10336_p4 = {{decipher_0_i32box_q62[31:24]}};

assign tmp_337_fu_10068_p4 = {{state_V_25_fu_10039_p2[23:16]}};

assign tmp_338_fu_10350_p4 = {{decipher_0_i32box_q61[15:8]}};

assign tmp_339_fu_10360_p4 = {{decipher_0_i32box_q61[23:16]}};

assign tmp_33_fu_4503_p4 = {{decipher_0_i32box_q139[31:24]}};

assign tmp_340_fu_10370_p4 = {{decipher_0_i32box_q61[31:24]}};

assign tmp_341_fu_10083_p4 = {{state_V_25_fu_10039_p2[31:24]}};

assign tmp_342_fu_10384_p4 = {{decipher_0_i32box_q60[15:8]}};

assign tmp_343_fu_10394_p4 = {{decipher_0_i32box_q60[23:16]}};

assign tmp_344_fu_10404_p4 = {{decipher_0_i32box_q60[31:24]}};

assign tmp_345_fu_10098_p4 = {{state_V_25_fu_10039_p2[39:32]}};

assign tmp_346_fu_10418_p4 = {{decipher_0_i32box_q59[15:8]}};

assign tmp_347_fu_10428_p4 = {{decipher_0_i32box_q59[23:16]}};

assign tmp_348_fu_10438_p4 = {{decipher_0_i32box_q59[31:24]}};

assign tmp_349_fu_10113_p4 = {{state_V_25_fu_10039_p2[47:40]}};

assign tmp_34_fu_4178_p4 = {{state_V_20_fu_4104_p2[47:40]}};

assign tmp_350_fu_10452_p4 = {{decipher_0_i32box_q58[15:8]}};

assign tmp_351_fu_10462_p4 = {{decipher_0_i32box_q58[23:16]}};

assign tmp_352_fu_10472_p4 = {{decipher_0_i32box_q58[31:24]}};

assign tmp_353_fu_10128_p4 = {{state_V_25_fu_10039_p2[55:48]}};

assign tmp_354_fu_10486_p4 = {{decipher_0_i32box_q57[15:8]}};

assign tmp_355_fu_10496_p4 = {{decipher_0_i32box_q57[23:16]}};

assign tmp_356_fu_10506_p4 = {{decipher_0_i32box_q57[31:24]}};

assign tmp_357_fu_10143_p4 = {{state_V_25_fu_10039_p2[63:56]}};

assign tmp_358_fu_10520_p4 = {{decipher_0_i32box_q56[15:8]}};

assign tmp_359_fu_10530_p4 = {{decipher_0_i32box_q56[23:16]}};

assign tmp_35_fu_4517_p4 = {{decipher_0_i32box_q138[15:8]}};

assign tmp_360_fu_10540_p4 = {{decipher_0_i32box_q56[31:24]}};

assign tmp_361_fu_10158_p4 = {{state_V_25_fu_10039_p2[71:64]}};

assign tmp_362_fu_10554_p4 = {{decipher_0_i32box_q55[15:8]}};

assign tmp_363_fu_10564_p4 = {{decipher_0_i32box_q55[23:16]}};

assign tmp_364_fu_10574_p4 = {{decipher_0_i32box_q55[31:24]}};

assign tmp_365_fu_10173_p4 = {{state_V_25_fu_10039_p2[79:72]}};

assign tmp_366_fu_10588_p4 = {{decipher_0_i32box_q54[15:8]}};

assign tmp_367_fu_10598_p4 = {{decipher_0_i32box_q54[23:16]}};

assign tmp_368_fu_10608_p4 = {{decipher_0_i32box_q54[31:24]}};

assign tmp_369_fu_10188_p4 = {{state_V_25_fu_10039_p2[87:80]}};

assign tmp_36_fu_4527_p4 = {{decipher_0_i32box_q138[23:16]}};

assign tmp_370_fu_10622_p4 = {{decipher_0_i32box_q53[15:8]}};

assign tmp_371_fu_10632_p4 = {{decipher_0_i32box_q53[23:16]}};

assign tmp_372_fu_10642_p4 = {{decipher_0_i32box_q53[31:24]}};

assign tmp_373_fu_10203_p4 = {{state_V_25_fu_10039_p2[95:88]}};

assign tmp_374_fu_10656_p4 = {{decipher_0_i32box_q52[15:8]}};

assign tmp_375_fu_10666_p4 = {{decipher_0_i32box_q52[23:16]}};

assign tmp_376_fu_10676_p4 = {{decipher_0_i32box_q52[31:24]}};

assign tmp_377_fu_10218_p4 = {{state_V_25_fu_10039_p2[103:96]}};

assign tmp_378_fu_10690_p4 = {{decipher_0_i32box_q51[15:8]}};

assign tmp_379_fu_10700_p4 = {{decipher_0_i32box_q51[23:16]}};

assign tmp_37_fu_4537_p4 = {{decipher_0_i32box_q138[31:24]}};

assign tmp_380_fu_10710_p4 = {{decipher_0_i32box_q51[31:24]}};

assign tmp_381_fu_10233_p4 = {{state_V_25_fu_10039_p2[111:104]}};

assign tmp_382_fu_10724_p4 = {{decipher_0_i32box_q50[15:8]}};

assign tmp_383_fu_10734_p4 = {{decipher_0_i32box_q50[23:16]}};

assign tmp_384_fu_10744_p4 = {{decipher_0_i32box_q50[31:24]}};

assign tmp_385_fu_10248_p4 = {{state_V_25_fu_10039_p2[119:112]}};

assign tmp_386_fu_10758_p4 = {{decipher_0_i32box_q49[15:8]}};

assign tmp_387_fu_10768_p4 = {{decipher_0_i32box_q49[23:16]}};

assign tmp_388_fu_10778_p4 = {{decipher_0_i32box_q49[31:24]}};

assign tmp_389_fu_10263_p4 = {{state_V_25_fu_10039_p2[127:120]}};

assign tmp_38_fu_4193_p4 = {{state_V_20_fu_4104_p2[55:48]}};

assign tmp_390_fu_10792_p4 = {{decipher_0_i32box_q48[15:8]}};

assign tmp_391_fu_10802_p4 = {{decipher_0_i32box_q48[23:16]}};

assign tmp_392_fu_10812_p4 = {{decipher_0_i32box_q48[31:24]}};

assign tmp_393_fu_11469_p4 = {{decipher_0_i32box_q47[15:8]}};

assign tmp_394_fu_11479_p4 = {{decipher_0_i32box_q47[23:16]}};

assign tmp_395_fu_11489_p4 = {{decipher_0_i32box_q47[31:24]}};

assign tmp_396_fu_11240_p4 = {{state_V_fu_11226_p2[15:8]}};

assign tmp_397_fu_11503_p4 = {{decipher_0_i32box_q46[15:8]}};

assign tmp_398_fu_11513_p4 = {{decipher_0_i32box_q46[23:16]}};

assign tmp_399_fu_11523_p4 = {{decipher_0_i32box_q46[31:24]}};

assign tmp_39_fu_4551_p4 = {{decipher_0_i32box_q137[15:8]}};

assign tmp_3_V_1_fu_6140_p2 = (xor_ln1545_62_fu_6134_p2 ^ xor_ln1545_61_fu_6128_p2);

assign tmp_3_V_2_fu_7327_p2 = (xor_ln1545_110_fu_7321_p2 ^ xor_ln1545_109_fu_7315_p2);

assign tmp_3_V_3_fu_8514_p2 = (xor_ln1545_158_fu_8508_p2 ^ xor_ln1545_157_fu_8502_p2);

assign tmp_3_V_4_fu_9701_p2 = (xor_ln1545_206_fu_9695_p2 ^ xor_ln1545_205_fu_9689_p2);

assign tmp_3_V_5_fu_10888_p2 = (xor_ln1545_254_fu_10882_p2 ^ xor_ln1545_253_fu_10876_p2);

assign tmp_3_V_6_fu_12075_p2 = (xor_ln1545_302_fu_12069_p2 ^ xor_ln1545_301_fu_12063_p2);

assign tmp_3_V_7_fu_13262_p2 = (xor_ln1545_350_fu_13256_p2 ^ xor_ln1545_349_fu_13250_p2);

assign tmp_3_V_8_fu_14449_p2 = (xor_ln1545_398_fu_14443_p2 ^ xor_ln1545_397_fu_14437_p2);

assign tmp_3_V_fu_4953_p2 = (xor_ln1545_14_fu_4947_p2 ^ xor_ln1545_13_fu_4941_p2);

assign tmp_3_fu_3873_p4 = {{ret_V_fu_3828_p2[63:56]}};

assign tmp_400_fu_11255_p4 = {{state_V_fu_11226_p2[23:16]}};

assign tmp_401_fu_11537_p4 = {{decipher_0_i32box_q45[15:8]}};

assign tmp_402_fu_11547_p4 = {{decipher_0_i32box_q45[23:16]}};

assign tmp_403_fu_11557_p4 = {{decipher_0_i32box_q45[31:24]}};

assign tmp_404_fu_11270_p4 = {{state_V_fu_11226_p2[31:24]}};

assign tmp_405_fu_11571_p4 = {{decipher_0_i32box_q44[15:8]}};

assign tmp_406_fu_11581_p4 = {{decipher_0_i32box_q44[23:16]}};

assign tmp_407_fu_11591_p4 = {{decipher_0_i32box_q44[31:24]}};

assign tmp_408_fu_11285_p4 = {{state_V_fu_11226_p2[39:32]}};

assign tmp_409_fu_11605_p4 = {{decipher_0_i32box_q43[15:8]}};

assign tmp_40_fu_4561_p4 = {{decipher_0_i32box_q137[23:16]}};

assign tmp_410_fu_11615_p4 = {{decipher_0_i32box_q43[23:16]}};

assign tmp_411_fu_11625_p4 = {{decipher_0_i32box_q43[31:24]}};

assign tmp_412_fu_11300_p4 = {{state_V_fu_11226_p2[47:40]}};

assign tmp_413_fu_11639_p4 = {{decipher_0_i32box_q42[15:8]}};

assign tmp_414_fu_11649_p4 = {{decipher_0_i32box_q42[23:16]}};

assign tmp_415_fu_11659_p4 = {{decipher_0_i32box_q42[31:24]}};

assign tmp_416_fu_11315_p4 = {{state_V_fu_11226_p2[55:48]}};

assign tmp_417_fu_11673_p4 = {{decipher_0_i32box_q41[15:8]}};

assign tmp_418_fu_11683_p4 = {{decipher_0_i32box_q41[23:16]}};

assign tmp_419_fu_11693_p4 = {{decipher_0_i32box_q41[31:24]}};

assign tmp_41_fu_4571_p4 = {{decipher_0_i32box_q137[31:24]}};

assign tmp_420_fu_11330_p4 = {{state_V_fu_11226_p2[63:56]}};

assign tmp_421_fu_11707_p4 = {{decipher_0_i32box_q40[15:8]}};

assign tmp_422_fu_11717_p4 = {{decipher_0_i32box_q40[23:16]}};

assign tmp_423_fu_11727_p4 = {{decipher_0_i32box_q40[31:24]}};

assign tmp_424_fu_11345_p4 = {{state_V_fu_11226_p2[71:64]}};

assign tmp_425_fu_11741_p4 = {{decipher_0_i32box_q39[15:8]}};

assign tmp_426_fu_11751_p4 = {{decipher_0_i32box_q39[23:16]}};

assign tmp_427_fu_11761_p4 = {{decipher_0_i32box_q39[31:24]}};

assign tmp_428_fu_11360_p4 = {{state_V_fu_11226_p2[79:72]}};

assign tmp_429_fu_11775_p4 = {{decipher_0_i32box_q38[15:8]}};

assign tmp_42_fu_4208_p4 = {{state_V_20_fu_4104_p2[63:56]}};

assign tmp_430_fu_11785_p4 = {{decipher_0_i32box_q38[23:16]}};

assign tmp_431_fu_11795_p4 = {{decipher_0_i32box_q38[31:24]}};

assign tmp_432_fu_11375_p4 = {{state_V_fu_11226_p2[87:80]}};

assign tmp_433_fu_11809_p4 = {{decipher_0_i32box_q37[15:8]}};

assign tmp_434_fu_11819_p4 = {{decipher_0_i32box_q37[23:16]}};

assign tmp_435_fu_11829_p4 = {{decipher_0_i32box_q37[31:24]}};

assign tmp_436_fu_11390_p4 = {{state_V_fu_11226_p2[95:88]}};

assign tmp_437_fu_11843_p4 = {{decipher_0_i32box_q36[15:8]}};

assign tmp_438_fu_11853_p4 = {{decipher_0_i32box_q36[23:16]}};

assign tmp_439_fu_11863_p4 = {{decipher_0_i32box_q36[31:24]}};

assign tmp_43_fu_4585_p4 = {{decipher_0_i32box_q136[15:8]}};

assign tmp_440_fu_11405_p4 = {{state_V_fu_11226_p2[103:96]}};

assign tmp_441_fu_11877_p4 = {{decipher_0_i32box_q35[15:8]}};

assign tmp_442_fu_11887_p4 = {{decipher_0_i32box_q35[23:16]}};

assign tmp_443_fu_11897_p4 = {{decipher_0_i32box_q35[31:24]}};

assign tmp_444_fu_11420_p4 = {{state_V_fu_11226_p2[111:104]}};

assign tmp_445_fu_11911_p4 = {{decipher_0_i32box_q34[15:8]}};

assign tmp_446_fu_11921_p4 = {{decipher_0_i32box_q34[23:16]}};

assign tmp_447_fu_11931_p4 = {{decipher_0_i32box_q34[31:24]}};

assign tmp_448_fu_11435_p4 = {{state_V_fu_11226_p2[119:112]}};

assign tmp_449_fu_11945_p4 = {{decipher_0_i32box_q33[15:8]}};

assign tmp_44_fu_4595_p4 = {{decipher_0_i32box_q136[23:16]}};

assign tmp_450_fu_11955_p4 = {{decipher_0_i32box_q33[23:16]}};

assign tmp_451_fu_11965_p4 = {{decipher_0_i32box_q33[31:24]}};

assign tmp_452_fu_11450_p4 = {{state_V_fu_11226_p2[127:120]}};

assign tmp_453_fu_11979_p4 = {{decipher_0_i32box_q32[15:8]}};

assign tmp_454_fu_11989_p4 = {{decipher_0_i32box_q32[23:16]}};

assign tmp_455_fu_11999_p4 = {{decipher_0_i32box_q32[31:24]}};

assign tmp_456_fu_12656_p4 = {{decipher_0_i32box_q31[15:8]}};

assign tmp_457_fu_12666_p4 = {{decipher_0_i32box_q31[23:16]}};

assign tmp_458_fu_12676_p4 = {{decipher_0_i32box_q31[31:24]}};

assign tmp_459_fu_12427_p4 = {{state_V_26_fu_12413_p2[15:8]}};

assign tmp_45_fu_4605_p4 = {{decipher_0_i32box_q136[31:24]}};

assign tmp_460_fu_12690_p4 = {{decipher_0_i32box_q30[15:8]}};

assign tmp_461_fu_12700_p4 = {{decipher_0_i32box_q30[23:16]}};

assign tmp_462_fu_12710_p4 = {{decipher_0_i32box_q30[31:24]}};

assign tmp_463_fu_12442_p4 = {{state_V_26_fu_12413_p2[23:16]}};

assign tmp_464_fu_12724_p4 = {{decipher_0_i32box_q29[15:8]}};

assign tmp_465_fu_12734_p4 = {{decipher_0_i32box_q29[23:16]}};

assign tmp_466_fu_12744_p4 = {{decipher_0_i32box_q29[31:24]}};

assign tmp_467_fu_12457_p4 = {{state_V_26_fu_12413_p2[31:24]}};

assign tmp_468_fu_12758_p4 = {{decipher_0_i32box_q28[15:8]}};

assign tmp_469_fu_12768_p4 = {{decipher_0_i32box_q28[23:16]}};

assign tmp_46_fu_4223_p4 = {{state_V_20_fu_4104_p2[71:64]}};

assign tmp_470_fu_12778_p4 = {{decipher_0_i32box_q28[31:24]}};

assign tmp_471_fu_12472_p4 = {{state_V_26_fu_12413_p2[39:32]}};

assign tmp_472_fu_12792_p4 = {{decipher_0_i32box_q27[15:8]}};

assign tmp_473_fu_12802_p4 = {{decipher_0_i32box_q27[23:16]}};

assign tmp_474_fu_12812_p4 = {{decipher_0_i32box_q27[31:24]}};

assign tmp_475_fu_12487_p4 = {{state_V_26_fu_12413_p2[47:40]}};

assign tmp_476_fu_12826_p4 = {{decipher_0_i32box_q26[15:8]}};

assign tmp_477_fu_12836_p4 = {{decipher_0_i32box_q26[23:16]}};

assign tmp_478_fu_12846_p4 = {{decipher_0_i32box_q26[31:24]}};

assign tmp_479_fu_12502_p4 = {{state_V_26_fu_12413_p2[55:48]}};

assign tmp_47_fu_4619_p4 = {{decipher_0_i32box_q135[15:8]}};

assign tmp_480_fu_12860_p4 = {{decipher_0_i32box_q25[15:8]}};

assign tmp_481_fu_12870_p4 = {{decipher_0_i32box_q25[23:16]}};

assign tmp_482_fu_12880_p4 = {{decipher_0_i32box_q25[31:24]}};

assign tmp_483_fu_12517_p4 = {{state_V_26_fu_12413_p2[63:56]}};

assign tmp_484_fu_12894_p4 = {{decipher_0_i32box_q24[15:8]}};

assign tmp_485_fu_12904_p4 = {{decipher_0_i32box_q24[23:16]}};

assign tmp_486_fu_12914_p4 = {{decipher_0_i32box_q24[31:24]}};

assign tmp_487_fu_12532_p4 = {{state_V_26_fu_12413_p2[71:64]}};

assign tmp_488_fu_12928_p4 = {{decipher_0_i32box_q23[15:8]}};

assign tmp_489_fu_12938_p4 = {{decipher_0_i32box_q23[23:16]}};

assign tmp_48_fu_4629_p4 = {{decipher_0_i32box_q135[23:16]}};

assign tmp_490_fu_12948_p4 = {{decipher_0_i32box_q23[31:24]}};

assign tmp_491_fu_12547_p4 = {{state_V_26_fu_12413_p2[79:72]}};

assign tmp_492_fu_12962_p4 = {{decipher_0_i32box_q22[15:8]}};

assign tmp_493_fu_12972_p4 = {{decipher_0_i32box_q22[23:16]}};

assign tmp_494_fu_12982_p4 = {{decipher_0_i32box_q22[31:24]}};

assign tmp_495_fu_12562_p4 = {{state_V_26_fu_12413_p2[87:80]}};

assign tmp_496_fu_12996_p4 = {{decipher_0_i32box_q21[15:8]}};

assign tmp_497_fu_13006_p4 = {{decipher_0_i32box_q21[23:16]}};

assign tmp_498_fu_13016_p4 = {{decipher_0_i32box_q21[31:24]}};

assign tmp_499_fu_12577_p4 = {{state_V_26_fu_12413_p2[95:88]}};

assign tmp_49_fu_4639_p4 = {{decipher_0_i32box_q135[31:24]}};

assign tmp_4_fu_3948_p4 = {{ret_V_fu_3828_p2[71:64]}};

assign tmp_500_fu_13030_p4 = {{decipher_0_i32box_q20[15:8]}};

assign tmp_501_fu_13040_p4 = {{decipher_0_i32box_q20[23:16]}};

assign tmp_502_fu_13050_p4 = {{decipher_0_i32box_q20[31:24]}};

assign tmp_503_fu_12592_p4 = {{state_V_26_fu_12413_p2[103:96]}};

assign tmp_504_fu_13064_p4 = {{decipher_0_i32box_q19[15:8]}};

assign tmp_505_fu_13074_p4 = {{decipher_0_i32box_q19[23:16]}};

assign tmp_506_fu_13084_p4 = {{decipher_0_i32box_q19[31:24]}};

assign tmp_507_fu_12607_p4 = {{state_V_26_fu_12413_p2[111:104]}};

assign tmp_508_fu_13098_p4 = {{decipher_0_i32box_q18[15:8]}};

assign tmp_509_fu_13108_p4 = {{decipher_0_i32box_q18[23:16]}};

assign tmp_50_fu_4238_p4 = {{state_V_20_fu_4104_p2[79:72]}};

assign tmp_510_fu_13118_p4 = {{decipher_0_i32box_q18[31:24]}};

assign tmp_511_fu_12622_p4 = {{state_V_26_fu_12413_p2[119:112]}};

assign tmp_512_fu_13132_p4 = {{decipher_0_i32box_q17[15:8]}};

assign tmp_513_fu_13142_p4 = {{decipher_0_i32box_q17[23:16]}};

assign tmp_514_fu_13152_p4 = {{decipher_0_i32box_q17[31:24]}};

assign tmp_515_fu_12637_p4 = {{state_V_26_fu_12413_p2[127:120]}};

assign tmp_516_fu_13166_p4 = {{decipher_0_i32box_q16[15:8]}};

assign tmp_517_fu_13176_p4 = {{decipher_0_i32box_q16[23:16]}};

assign tmp_518_fu_13186_p4 = {{decipher_0_i32box_q16[31:24]}};

assign tmp_519_fu_13843_p4 = {{decipher_0_i32box_q15[15:8]}};

assign tmp_51_fu_4653_p4 = {{decipher_0_i32box_q134[15:8]}};

assign tmp_520_fu_13853_p4 = {{decipher_0_i32box_q15[23:16]}};

assign tmp_521_fu_13863_p4 = {{decipher_0_i32box_q15[31:24]}};

assign tmp_522_fu_13614_p4 = {{state_V_27_fu_13600_p2[15:8]}};

assign tmp_523_fu_13877_p4 = {{decipher_0_i32box_q14[15:8]}};

assign tmp_524_fu_13887_p4 = {{decipher_0_i32box_q14[23:16]}};

assign tmp_525_fu_13897_p4 = {{decipher_0_i32box_q14[31:24]}};

assign tmp_526_fu_13629_p4 = {{state_V_27_fu_13600_p2[23:16]}};

assign tmp_527_fu_13911_p4 = {{decipher_0_i32box_q13[15:8]}};

assign tmp_528_fu_13921_p4 = {{decipher_0_i32box_q13[23:16]}};

assign tmp_529_fu_13931_p4 = {{decipher_0_i32box_q13[31:24]}};

assign tmp_52_fu_4663_p4 = {{decipher_0_i32box_q134[23:16]}};

assign tmp_530_fu_13644_p4 = {{state_V_27_fu_13600_p2[31:24]}};

assign tmp_531_fu_13945_p4 = {{decipher_0_i32box_q12[15:8]}};

assign tmp_532_fu_13955_p4 = {{decipher_0_i32box_q12[23:16]}};

assign tmp_533_fu_13965_p4 = {{decipher_0_i32box_q12[31:24]}};

assign tmp_534_fu_13659_p4 = {{state_V_27_fu_13600_p2[39:32]}};

assign tmp_535_fu_13979_p4 = {{decipher_0_i32box_q11[15:8]}};

assign tmp_536_fu_13989_p4 = {{decipher_0_i32box_q11[23:16]}};

assign tmp_537_fu_13999_p4 = {{decipher_0_i32box_q11[31:24]}};

assign tmp_538_fu_13674_p4 = {{state_V_27_fu_13600_p2[47:40]}};

assign tmp_539_fu_14013_p4 = {{decipher_0_i32box_q10[15:8]}};

assign tmp_53_fu_4673_p4 = {{decipher_0_i32box_q134[31:24]}};

assign tmp_540_fu_14023_p4 = {{decipher_0_i32box_q10[23:16]}};

assign tmp_541_fu_14033_p4 = {{decipher_0_i32box_q10[31:24]}};

assign tmp_542_fu_13689_p4 = {{state_V_27_fu_13600_p2[55:48]}};

assign tmp_543_fu_14047_p4 = {{decipher_0_i32box_q9[15:8]}};

assign tmp_544_fu_14057_p4 = {{decipher_0_i32box_q9[23:16]}};

assign tmp_545_fu_14067_p4 = {{decipher_0_i32box_q9[31:24]}};

assign tmp_546_fu_13704_p4 = {{state_V_27_fu_13600_p2[63:56]}};

assign tmp_547_fu_14081_p4 = {{decipher_0_i32box_q8[15:8]}};

assign tmp_548_fu_14091_p4 = {{decipher_0_i32box_q8[23:16]}};

assign tmp_549_fu_14101_p4 = {{decipher_0_i32box_q8[31:24]}};

assign tmp_54_fu_4253_p4 = {{state_V_20_fu_4104_p2[87:80]}};

assign tmp_550_fu_13719_p4 = {{state_V_27_fu_13600_p2[71:64]}};

assign tmp_551_fu_14115_p4 = {{decipher_0_i32box_q7[15:8]}};

assign tmp_552_fu_14125_p4 = {{decipher_0_i32box_q7[23:16]}};

assign tmp_553_fu_14135_p4 = {{decipher_0_i32box_q7[31:24]}};

assign tmp_554_fu_13734_p4 = {{state_V_27_fu_13600_p2[79:72]}};

assign tmp_555_fu_14149_p4 = {{decipher_0_i32box_q6[15:8]}};

assign tmp_556_fu_14159_p4 = {{decipher_0_i32box_q6[23:16]}};

assign tmp_557_fu_14169_p4 = {{decipher_0_i32box_q6[31:24]}};

assign tmp_558_fu_13749_p4 = {{state_V_27_fu_13600_p2[87:80]}};

assign tmp_559_fu_14183_p4 = {{decipher_0_i32box_q5[15:8]}};

assign tmp_55_fu_4687_p4 = {{decipher_0_i32box_q133[15:8]}};

assign tmp_560_fu_14193_p4 = {{decipher_0_i32box_q5[23:16]}};

assign tmp_561_fu_14203_p4 = {{decipher_0_i32box_q5[31:24]}};

assign tmp_562_fu_13764_p4 = {{state_V_27_fu_13600_p2[95:88]}};

assign tmp_563_fu_14217_p4 = {{decipher_0_i32box_q4[15:8]}};

assign tmp_564_fu_14227_p4 = {{decipher_0_i32box_q4[23:16]}};

assign tmp_565_fu_14237_p4 = {{decipher_0_i32box_q4[31:24]}};

assign tmp_566_fu_13779_p4 = {{state_V_27_fu_13600_p2[103:96]}};

assign tmp_567_fu_14251_p4 = {{decipher_0_i32box_q3[15:8]}};

assign tmp_568_fu_14261_p4 = {{decipher_0_i32box_q3[23:16]}};

assign tmp_569_fu_14271_p4 = {{decipher_0_i32box_q3[31:24]}};

assign tmp_56_fu_4697_p4 = {{decipher_0_i32box_q133[23:16]}};

assign tmp_570_fu_13794_p4 = {{state_V_27_fu_13600_p2[111:104]}};

assign tmp_571_fu_14285_p4 = {{decipher_0_i32box_q2[15:8]}};

assign tmp_572_fu_14295_p4 = {{decipher_0_i32box_q2[23:16]}};

assign tmp_573_fu_14305_p4 = {{decipher_0_i32box_q2[31:24]}};

assign tmp_574_fu_13809_p4 = {{state_V_27_fu_13600_p2[119:112]}};

assign tmp_575_fu_14319_p4 = {{decipher_0_i32box_q1[15:8]}};

assign tmp_576_fu_14329_p4 = {{decipher_0_i32box_q1[23:16]}};

assign tmp_577_fu_14339_p4 = {{decipher_0_i32box_q1[31:24]}};

assign tmp_578_fu_13824_p4 = {{state_V_27_fu_13600_p2[127:120]}};

assign tmp_579_fu_14353_p4 = {{decipher_0_i32box_q0[15:8]}};

assign tmp_57_fu_4707_p4 = {{decipher_0_i32box_q133[31:24]}};

assign tmp_580_fu_14363_p4 = {{decipher_0_i32box_q0[23:16]}};

assign tmp_581_fu_14373_p4 = {{decipher_0_i32box_q0[31:24]}};

assign tmp_58_fu_4268_p4 = {{state_V_20_fu_4104_p2[95:88]}};

assign tmp_59_fu_4721_p4 = {{decipher_0_i32box_q132[15:8]}};

assign tmp_5_fu_3903_p4 = {{ret_V_fu_3828_p2[15:8]}};

assign tmp_60_fu_4731_p4 = {{decipher_0_i32box_q132[23:16]}};

assign tmp_61_fu_4741_p4 = {{decipher_0_i32box_q132[31:24]}};

assign tmp_62_fu_4283_p4 = {{state_V_20_fu_4104_p2[103:96]}};

assign tmp_63_fu_4755_p4 = {{decipher_0_i32box_q131[15:8]}};

assign tmp_64_fu_4765_p4 = {{decipher_0_i32box_q131[23:16]}};

assign tmp_65_fu_4775_p4 = {{decipher_0_i32box_q131[31:24]}};

assign tmp_66_fu_4298_p4 = {{state_V_20_fu_4104_p2[111:104]}};

assign tmp_67_fu_4789_p4 = {{decipher_0_i32box_q130[15:8]}};

assign tmp_68_fu_4799_p4 = {{decipher_0_i32box_q130[23:16]}};

assign tmp_69_fu_4809_p4 = {{decipher_0_i32box_q130[31:24]}};

assign tmp_6_fu_3918_p4 = {{ret_V_fu_3828_p2[119:112]}};

assign tmp_70_fu_4313_p4 = {{state_V_20_fu_4104_p2[119:112]}};

assign tmp_71_fu_4823_p4 = {{decipher_0_i32box_q129[15:8]}};

assign tmp_72_fu_4833_p4 = {{decipher_0_i32box_q129[23:16]}};

assign tmp_73_fu_4843_p4 = {{decipher_0_i32box_q129[31:24]}};

assign tmp_74_fu_4328_p4 = {{state_V_20_fu_4104_p2[127:120]}};

assign tmp_75_fu_4857_p4 = {{decipher_0_i32box_q128[15:8]}};

assign tmp_76_fu_4867_p4 = {{decipher_0_i32box_q128[23:16]}};

assign tmp_77_fu_4877_p4 = {{decipher_0_i32box_q128[31:24]}};

assign tmp_78_fu_5534_p4 = {{decipher_0_i32box_q127[15:8]}};

assign tmp_79_fu_5544_p4 = {{decipher_0_i32box_q127[23:16]}};

assign tmp_7_fu_3933_p4 = {{ret_V_fu_3828_p2[95:88]}};

assign tmp_80_fu_5554_p4 = {{decipher_0_i32box_q127[31:24]}};

assign tmp_81_fu_5305_p4 = {{state_V_21_fu_5291_p2[15:8]}};

assign tmp_82_fu_5568_p4 = {{decipher_0_i32box_q126[15:8]}};

assign tmp_83_fu_5578_p4 = {{decipher_0_i32box_q126[23:16]}};

assign tmp_84_fu_5588_p4 = {{decipher_0_i32box_q126[31:24]}};

assign tmp_85_fu_5320_p4 = {{state_V_21_fu_5291_p2[23:16]}};

assign tmp_86_fu_5602_p4 = {{decipher_0_i32box_q125[15:8]}};

assign tmp_87_fu_5612_p4 = {{decipher_0_i32box_q125[23:16]}};

assign tmp_88_fu_5622_p4 = {{decipher_0_i32box_q125[31:24]}};

assign tmp_89_fu_5335_p4 = {{state_V_21_fu_5291_p2[31:24]}};

assign tmp_8_fu_3978_p4 = {{ret_V_fu_3828_p2[23:16]}};

assign tmp_90_fu_5636_p4 = {{decipher_0_i32box_q124[15:8]}};

assign tmp_91_fu_5646_p4 = {{decipher_0_i32box_q124[23:16]}};

assign tmp_92_fu_5656_p4 = {{decipher_0_i32box_q124[31:24]}};

assign tmp_93_fu_5350_p4 = {{state_V_21_fu_5291_p2[39:32]}};

assign tmp_94_fu_5670_p4 = {{decipher_0_i32box_q123[15:8]}};

assign tmp_95_fu_5680_p4 = {{decipher_0_i32box_q123[23:16]}};

assign tmp_96_fu_5690_p4 = {{decipher_0_i32box_q123[31:24]}};

assign tmp_97_fu_5365_p4 = {{state_V_21_fu_5291_p2[47:40]}};

assign tmp_98_fu_5704_p4 = {{decipher_0_i32box_q122[15:8]}};

assign tmp_99_fu_5714_p4 = {{decipher_0_i32box_q122[23:16]}};

assign tmp_9_fu_3963_p4 = {{ret_V_fu_3828_p2[47:40]}};

assign tmp_s_fu_3888_p4 = {{ret_V_fu_3828_p2[39:32]}};

assign trunc_ln674_100_fu_11601_p1 = decipher_0_i32box_q43[7:0];

assign trunc_ln674_101_fu_11635_p1 = decipher_0_i32box_q42[7:0];

assign trunc_ln674_102_fu_11669_p1 = decipher_0_i32box_q41[7:0];

assign trunc_ln674_103_fu_11703_p1 = decipher_0_i32box_q40[7:0];

assign trunc_ln674_104_fu_11737_p1 = decipher_0_i32box_q39[7:0];

assign trunc_ln674_105_fu_11771_p1 = decipher_0_i32box_q38[7:0];

assign trunc_ln674_106_fu_11805_p1 = decipher_0_i32box_q37[7:0];

assign trunc_ln674_107_fu_11839_p1 = decipher_0_i32box_q36[7:0];

assign trunc_ln674_108_fu_11873_p1 = decipher_0_i32box_q35[7:0];

assign trunc_ln674_109_fu_11907_p1 = decipher_0_i32box_q34[7:0];

assign trunc_ln674_10_fu_4683_p1 = decipher_0_i32box_q133[7:0];

assign trunc_ln674_110_fu_11941_p1 = decipher_0_i32box_q33[7:0];

assign trunc_ln674_111_fu_11975_p1 = decipher_0_i32box_q32[7:0];

assign trunc_ln674_112_fu_12652_p1 = decipher_0_i32box_q31[7:0];

assign trunc_ln674_113_fu_12686_p1 = decipher_0_i32box_q30[7:0];

assign trunc_ln674_114_fu_12720_p1 = decipher_0_i32box_q29[7:0];

assign trunc_ln674_115_fu_12754_p1 = decipher_0_i32box_q28[7:0];

assign trunc_ln674_116_fu_12788_p1 = decipher_0_i32box_q27[7:0];

assign trunc_ln674_117_fu_12822_p1 = decipher_0_i32box_q26[7:0];

assign trunc_ln674_118_fu_12856_p1 = decipher_0_i32box_q25[7:0];

assign trunc_ln674_119_fu_12890_p1 = decipher_0_i32box_q24[7:0];

assign trunc_ln674_11_fu_4717_p1 = decipher_0_i32box_q132[7:0];

assign trunc_ln674_120_fu_12924_p1 = decipher_0_i32box_q23[7:0];

assign trunc_ln674_121_fu_12958_p1 = decipher_0_i32box_q22[7:0];

assign trunc_ln674_122_fu_12992_p1 = decipher_0_i32box_q21[7:0];

assign trunc_ln674_123_fu_13026_p1 = decipher_0_i32box_q20[7:0];

assign trunc_ln674_124_fu_13060_p1 = decipher_0_i32box_q19[7:0];

assign trunc_ln674_125_fu_13094_p1 = decipher_0_i32box_q18[7:0];

assign trunc_ln674_126_fu_13128_p1 = decipher_0_i32box_q17[7:0];

assign trunc_ln674_127_fu_13162_p1 = decipher_0_i32box_q16[7:0];

assign trunc_ln674_128_fu_13839_p1 = decipher_0_i32box_q15[7:0];

assign trunc_ln674_129_fu_13873_p1 = decipher_0_i32box_q14[7:0];

assign trunc_ln674_12_fu_4751_p1 = decipher_0_i32box_q131[7:0];

assign trunc_ln674_130_fu_13907_p1 = decipher_0_i32box_q13[7:0];

assign trunc_ln674_131_fu_13941_p1 = decipher_0_i32box_q12[7:0];

assign trunc_ln674_132_fu_13975_p1 = decipher_0_i32box_q11[7:0];

assign trunc_ln674_133_fu_14009_p1 = decipher_0_i32box_q10[7:0];

assign trunc_ln674_134_fu_14043_p1 = decipher_0_i32box_q9[7:0];

assign trunc_ln674_135_fu_14077_p1 = decipher_0_i32box_q8[7:0];

assign trunc_ln674_136_fu_14111_p1 = decipher_0_i32box_q7[7:0];

assign trunc_ln674_137_fu_14145_p1 = decipher_0_i32box_q6[7:0];

assign trunc_ln674_138_fu_14179_p1 = decipher_0_i32box_q5[7:0];

assign trunc_ln674_139_fu_14213_p1 = decipher_0_i32box_q4[7:0];

assign trunc_ln674_13_fu_4785_p1 = decipher_0_i32box_q130[7:0];

assign trunc_ln674_140_fu_14247_p1 = decipher_0_i32box_q3[7:0];

assign trunc_ln674_141_fu_14281_p1 = decipher_0_i32box_q2[7:0];

assign trunc_ln674_142_fu_14315_p1 = decipher_0_i32box_q1[7:0];

assign trunc_ln674_143_fu_14349_p1 = decipher_0_i32box_q0[7:0];

assign trunc_ln674_14_fu_4819_p1 = decipher_0_i32box_q129[7:0];

assign trunc_ln674_15_fu_4853_p1 = decipher_0_i32box_q128[7:0];

assign trunc_ln674_16_fu_5530_p1 = decipher_0_i32box_q127[7:0];

assign trunc_ln674_17_fu_5564_p1 = decipher_0_i32box_q126[7:0];

assign trunc_ln674_18_fu_5598_p1 = decipher_0_i32box_q125[7:0];

assign trunc_ln674_19_fu_5632_p1 = decipher_0_i32box_q124[7:0];

assign trunc_ln674_1_fu_4377_p1 = decipher_0_i32box_q142[7:0];

assign trunc_ln674_20_fu_5666_p1 = decipher_0_i32box_q123[7:0];

assign trunc_ln674_21_fu_5700_p1 = decipher_0_i32box_q122[7:0];

assign trunc_ln674_22_fu_5734_p1 = decipher_0_i32box_q121[7:0];

assign trunc_ln674_23_fu_5768_p1 = decipher_0_i32box_q120[7:0];

assign trunc_ln674_24_fu_5802_p1 = decipher_0_i32box_q119[7:0];

assign trunc_ln674_25_fu_5836_p1 = decipher_0_i32box_q118[7:0];

assign trunc_ln674_26_fu_5870_p1 = decipher_0_i32box_q117[7:0];

assign trunc_ln674_27_fu_5904_p1 = decipher_0_i32box_q116[7:0];

assign trunc_ln674_28_fu_5938_p1 = decipher_0_i32box_q115[7:0];

assign trunc_ln674_29_fu_5972_p1 = decipher_0_i32box_q114[7:0];

assign trunc_ln674_2_fu_4411_p1 = decipher_0_i32box_q141[7:0];

assign trunc_ln674_30_fu_6006_p1 = decipher_0_i32box_q113[7:0];

assign trunc_ln674_31_fu_6040_p1 = decipher_0_i32box_q112[7:0];

assign trunc_ln674_32_fu_6717_p1 = decipher_0_i32box_q111[7:0];

assign trunc_ln674_33_fu_6751_p1 = decipher_0_i32box_q110[7:0];

assign trunc_ln674_34_fu_6785_p1 = decipher_0_i32box_q109[7:0];

assign trunc_ln674_35_fu_6819_p1 = decipher_0_i32box_q108[7:0];

assign trunc_ln674_36_fu_6853_p1 = decipher_0_i32box_q107[7:0];

assign trunc_ln674_37_fu_6887_p1 = decipher_0_i32box_q106[7:0];

assign trunc_ln674_38_fu_6921_p1 = decipher_0_i32box_q105[7:0];

assign trunc_ln674_39_fu_6955_p1 = decipher_0_i32box_q104[7:0];

assign trunc_ln674_3_fu_4445_p1 = decipher_0_i32box_q140[7:0];

assign trunc_ln674_40_fu_6989_p1 = decipher_0_i32box_q103[7:0];

assign trunc_ln674_41_fu_7023_p1 = decipher_0_i32box_q102[7:0];

assign trunc_ln674_42_fu_7057_p1 = decipher_0_i32box_q101[7:0];

assign trunc_ln674_43_fu_7091_p1 = decipher_0_i32box_q100[7:0];

assign trunc_ln674_44_fu_7125_p1 = decipher_0_i32box_q99[7:0];

assign trunc_ln674_45_fu_7159_p1 = decipher_0_i32box_q98[7:0];

assign trunc_ln674_46_fu_7193_p1 = decipher_0_i32box_q97[7:0];

assign trunc_ln674_47_fu_7227_p1 = decipher_0_i32box_q96[7:0];

assign trunc_ln674_48_fu_7904_p1 = decipher_0_i32box_q95[7:0];

assign trunc_ln674_49_fu_7938_p1 = decipher_0_i32box_q94[7:0];

assign trunc_ln674_4_fu_4479_p1 = decipher_0_i32box_q139[7:0];

assign trunc_ln674_50_fu_7972_p1 = decipher_0_i32box_q93[7:0];

assign trunc_ln674_51_fu_8006_p1 = decipher_0_i32box_q92[7:0];

assign trunc_ln674_52_fu_8040_p1 = decipher_0_i32box_q91[7:0];

assign trunc_ln674_53_fu_8074_p1 = decipher_0_i32box_q90[7:0];

assign trunc_ln674_54_fu_8108_p1 = decipher_0_i32box_q89[7:0];

assign trunc_ln674_55_fu_8142_p1 = decipher_0_i32box_q88[7:0];

assign trunc_ln674_56_fu_8176_p1 = decipher_0_i32box_q87[7:0];

assign trunc_ln674_57_fu_8210_p1 = decipher_0_i32box_q86[7:0];

assign trunc_ln674_58_fu_8244_p1 = decipher_0_i32box_q85[7:0];

assign trunc_ln674_59_fu_8278_p1 = decipher_0_i32box_q84[7:0];

assign trunc_ln674_5_fu_4513_p1 = decipher_0_i32box_q138[7:0];

assign trunc_ln674_60_fu_8312_p1 = decipher_0_i32box_q83[7:0];

assign trunc_ln674_61_fu_8346_p1 = decipher_0_i32box_q82[7:0];

assign trunc_ln674_62_fu_8380_p1 = decipher_0_i32box_q81[7:0];

assign trunc_ln674_63_fu_8414_p1 = decipher_0_i32box_q80[7:0];

assign trunc_ln674_64_fu_9091_p1 = decipher_0_i32box_q79[7:0];

assign trunc_ln674_65_fu_9125_p1 = decipher_0_i32box_q78[7:0];

assign trunc_ln674_66_fu_9159_p1 = decipher_0_i32box_q77[7:0];

assign trunc_ln674_67_fu_9193_p1 = decipher_0_i32box_q76[7:0];

assign trunc_ln674_68_fu_9227_p1 = decipher_0_i32box_q75[7:0];

assign trunc_ln674_69_fu_9261_p1 = decipher_0_i32box_q74[7:0];

assign trunc_ln674_6_fu_4547_p1 = decipher_0_i32box_q137[7:0];

assign trunc_ln674_70_fu_9295_p1 = decipher_0_i32box_q73[7:0];

assign trunc_ln674_71_fu_9329_p1 = decipher_0_i32box_q72[7:0];

assign trunc_ln674_72_fu_9363_p1 = decipher_0_i32box_q71[7:0];

assign trunc_ln674_73_fu_9397_p1 = decipher_0_i32box_q70[7:0];

assign trunc_ln674_74_fu_9431_p1 = decipher_0_i32box_q69[7:0];

assign trunc_ln674_75_fu_9465_p1 = decipher_0_i32box_q68[7:0];

assign trunc_ln674_76_fu_9499_p1 = decipher_0_i32box_q67[7:0];

assign trunc_ln674_77_fu_9533_p1 = decipher_0_i32box_q66[7:0];

assign trunc_ln674_78_fu_9567_p1 = decipher_0_i32box_q65[7:0];

assign trunc_ln674_79_fu_9601_p1 = decipher_0_i32box_q64[7:0];

assign trunc_ln674_7_fu_4581_p1 = decipher_0_i32box_q136[7:0];

assign trunc_ln674_80_fu_10278_p1 = decipher_0_i32box_q63[7:0];

assign trunc_ln674_81_fu_10312_p1 = decipher_0_i32box_q62[7:0];

assign trunc_ln674_82_fu_10346_p1 = decipher_0_i32box_q61[7:0];

assign trunc_ln674_83_fu_10380_p1 = decipher_0_i32box_q60[7:0];

assign trunc_ln674_84_fu_10414_p1 = decipher_0_i32box_q59[7:0];

assign trunc_ln674_85_fu_10448_p1 = decipher_0_i32box_q58[7:0];

assign trunc_ln674_86_fu_10482_p1 = decipher_0_i32box_q57[7:0];

assign trunc_ln674_87_fu_10516_p1 = decipher_0_i32box_q56[7:0];

assign trunc_ln674_88_fu_10550_p1 = decipher_0_i32box_q55[7:0];

assign trunc_ln674_89_fu_10584_p1 = decipher_0_i32box_q54[7:0];

assign trunc_ln674_8_fu_4615_p1 = decipher_0_i32box_q135[7:0];

assign trunc_ln674_90_fu_10618_p1 = decipher_0_i32box_q53[7:0];

assign trunc_ln674_91_fu_10652_p1 = decipher_0_i32box_q52[7:0];

assign trunc_ln674_92_fu_10686_p1 = decipher_0_i32box_q51[7:0];

assign trunc_ln674_93_fu_10720_p1 = decipher_0_i32box_q50[7:0];

assign trunc_ln674_94_fu_10754_p1 = decipher_0_i32box_q49[7:0];

assign trunc_ln674_95_fu_10788_p1 = decipher_0_i32box_q48[7:0];

assign trunc_ln674_96_fu_11465_p1 = decipher_0_i32box_q47[7:0];

assign trunc_ln674_97_fu_11499_p1 = decipher_0_i32box_q46[7:0];

assign trunc_ln674_98_fu_11533_p1 = decipher_0_i32box_q45[7:0];

assign trunc_ln674_99_fu_11567_p1 = decipher_0_i32box_q44[7:0];

assign trunc_ln674_9_fu_4649_p1 = decipher_0_i32box_q134[7:0];

assign trunc_ln674_fu_4343_p1 = decipher_0_i32box_q143[7:0];

assign trunc_ln708_1_fu_4109_p1 = state_V_20_fu_4104_p2[7:0];

assign trunc_ln708_2_fu_5296_p1 = state_V_21_fu_5291_p2[7:0];

assign trunc_ln708_3_fu_6483_p1 = state_V_22_fu_6478_p2[7:0];

assign trunc_ln708_4_fu_7670_p1 = state_V_23_fu_7665_p2[7:0];

assign trunc_ln708_5_fu_8857_p1 = state_V_24_fu_8852_p2[7:0];

assign trunc_ln708_6_fu_10044_p1 = state_V_25_fu_10039_p2[7:0];

assign trunc_ln708_7_fu_11231_p1 = state_V_fu_11226_p2[7:0];

assign trunc_ln708_8_fu_12418_p1 = state_V_26_fu_12413_p2[7:0];

assign trunc_ln708_9_fu_13605_p1 = state_V_27_fu_13600_p2[7:0];

assign trunc_ln708_fu_3834_p1 = ret_V_fu_3828_p2[7:0];

assign xor_ln1545_100_fu_7261_p2 = (tmp_145_fu_6755_p4 ^ tmp_143_fu_6741_p4);

assign xor_ln1545_101_fu_7273_p2 = (xor_ln1545_102_fu_7267_p2 ^ xor_ln1545_100_fu_7261_p2);

assign xor_ln1545_102_fu_7267_p2 = (trunc_ln674_35_fu_6819_p1 ^ tmp_150_fu_6799_p4);

assign xor_ln1545_103_fu_7279_p2 = (trunc_ln674_32_fu_6717_p1 ^ tmp_147_fu_6775_p4);

assign xor_ln1545_104_fu_7291_p2 = (xor_ln1545_105_fu_7285_p2 ^ xor_ln1545_103_fu_7279_p2);

assign xor_ln1545_105_fu_7285_p2 = (tmp_154_fu_6833_p4 ^ tmp_149_fu_6789_p4);

assign xor_ln1545_106_fu_7297_p2 = (trunc_ln674_33_fu_6751_p1 ^ tmp_142_fu_6731_p4);

assign xor_ln1545_107_fu_7309_p2 = (xor_ln1545_108_fu_7303_p2 ^ xor_ln1545_106_fu_7297_p2);

assign xor_ln1545_108_fu_7303_p2 = (tmp_153_fu_6823_p4 ^ tmp_151_fu_6809_p4);

assign xor_ln1545_109_fu_7315_p2 = (tmp_146_fu_6765_p4 ^ tmp_141_fu_6721_p4);

assign xor_ln1545_10_fu_4923_p2 = (trunc_ln674_1_fu_4377_p1 ^ tmp_16_fu_4357_p4);

assign xor_ln1545_110_fu_7321_p2 = (trunc_ln674_34_fu_6785_p1 ^ tmp_155_fu_6843_p4);

assign xor_ln1545_112_fu_7333_p2 = (tmp_161_fu_6891_p4 ^ tmp_159_fu_6877_p4);

assign xor_ln1545_113_fu_7345_p2 = (xor_ln1545_114_fu_7339_p2 ^ xor_ln1545_112_fu_7333_p2);

assign xor_ln1545_114_fu_7339_p2 = (trunc_ln674_39_fu_6955_p1 ^ tmp_166_fu_6935_p4);

assign xor_ln1545_115_fu_7351_p2 = (trunc_ln674_36_fu_6853_p1 ^ tmp_163_fu_6911_p4);

assign xor_ln1545_116_fu_7363_p2 = (xor_ln1545_117_fu_7357_p2 ^ xor_ln1545_115_fu_7351_p2);

assign xor_ln1545_117_fu_7357_p2 = (tmp_170_fu_6969_p4 ^ tmp_165_fu_6925_p4);

assign xor_ln1545_118_fu_7369_p2 = (trunc_ln674_37_fu_6887_p1 ^ tmp_158_fu_6867_p4);

assign xor_ln1545_119_fu_7381_p2 = (xor_ln1545_120_fu_7375_p2 ^ xor_ln1545_118_fu_7369_p2);

assign xor_ln1545_11_fu_4935_p2 = (xor_ln1545_12_fu_4929_p2 ^ xor_ln1545_10_fu_4923_p2);

assign xor_ln1545_120_fu_7375_p2 = (tmp_169_fu_6959_p4 ^ tmp_167_fu_6945_p4);

assign xor_ln1545_121_fu_7387_p2 = (tmp_162_fu_6901_p4 ^ tmp_157_fu_6857_p4);

assign xor_ln1545_122_fu_7399_p2 = (xor_ln1545_123_fu_7393_p2 ^ xor_ln1545_121_fu_7387_p2);

assign xor_ln1545_123_fu_7393_p2 = (trunc_ln674_38_fu_6921_p1 ^ tmp_171_fu_6979_p4);

assign xor_ln1545_124_fu_7405_p2 = (tmp_177_fu_7027_p4 ^ tmp_175_fu_7013_p4);

assign xor_ln1545_125_fu_7417_p2 = (xor_ln1545_126_fu_7411_p2 ^ xor_ln1545_124_fu_7405_p2);

assign xor_ln1545_126_fu_7411_p2 = (trunc_ln674_43_fu_7091_p1 ^ tmp_182_fu_7071_p4);

assign xor_ln1545_127_fu_7423_p2 = (trunc_ln674_40_fu_6989_p1 ^ tmp_179_fu_7047_p4);

assign xor_ln1545_128_fu_7435_p2 = (xor_ln1545_129_fu_7429_p2 ^ xor_ln1545_127_fu_7423_p2);

assign xor_ln1545_129_fu_7429_p2 = (tmp_186_fu_7105_p4 ^ tmp_181_fu_7061_p4);

assign xor_ln1545_12_fu_4929_p2 = (tmp_27_fu_4449_p4 ^ tmp_25_fu_4435_p4);

assign xor_ln1545_130_fu_7441_p2 = (trunc_ln674_41_fu_7023_p1 ^ tmp_174_fu_7003_p4);

assign xor_ln1545_131_fu_7447_p2 = (tmp_185_fu_7095_p4 ^ tmp_183_fu_7081_p4);

assign xor_ln1545_133_fu_7459_p2 = (tmp_178_fu_7037_p4 ^ tmp_173_fu_6993_p4);

assign xor_ln1545_134_fu_7471_p2 = (xor_ln1545_135_fu_7465_p2 ^ xor_ln1545_133_fu_7459_p2);

assign xor_ln1545_135_fu_7465_p2 = (trunc_ln674_42_fu_7057_p1 ^ tmp_187_fu_7115_p4);

assign xor_ln1545_136_fu_7477_p2 = (tmp_193_fu_7163_p4 ^ tmp_191_fu_7149_p4);

assign xor_ln1545_137_fu_7489_p2 = (xor_ln1545_138_fu_7483_p2 ^ xor_ln1545_136_fu_7477_p2);

assign xor_ln1545_138_fu_7483_p2 = (trunc_ln674_47_fu_7227_p1 ^ tmp_198_fu_7207_p4);

assign xor_ln1545_139_fu_7495_p2 = (trunc_ln674_44_fu_7125_p1 ^ tmp_195_fu_7183_p4);

assign xor_ln1545_13_fu_4941_p2 = (tmp_20_fu_4391_p4 ^ tmp_15_fu_4347_p4);

assign xor_ln1545_140_fu_7501_p2 = (tmp_202_fu_7241_p4 ^ tmp_197_fu_7197_p4);

assign xor_ln1545_142_fu_7513_p2 = (trunc_ln674_45_fu_7159_p1 ^ tmp_190_fu_7139_p4);

assign xor_ln1545_143_fu_7519_p2 = (tmp_201_fu_7231_p4 ^ tmp_199_fu_7217_p4);

assign xor_ln1545_145_fu_7531_p2 = (tmp_194_fu_7173_p4 ^ tmp_189_fu_7129_p4);

assign xor_ln1545_146_fu_7543_p2 = (xor_ln1545_147_fu_7537_p2 ^ xor_ln1545_145_fu_7531_p2);

assign xor_ln1545_147_fu_7537_p2 = (trunc_ln674_46_fu_7193_p1 ^ tmp_203_fu_7251_p4);

assign xor_ln1545_148_fu_8448_p2 = (tmp_208_fu_7942_p4 ^ tmp_206_fu_7928_p4);

assign xor_ln1545_149_fu_8460_p2 = (xor_ln1545_150_fu_8454_p2 ^ xor_ln1545_148_fu_8448_p2);

assign xor_ln1545_14_fu_4947_p2 = (trunc_ln674_2_fu_4411_p1 ^ tmp_29_fu_4469_p4);

assign xor_ln1545_150_fu_8454_p2 = (trunc_ln674_51_fu_8006_p1 ^ tmp_213_fu_7986_p4);

assign xor_ln1545_151_fu_8466_p2 = (trunc_ln674_48_fu_7904_p1 ^ tmp_210_fu_7962_p4);

assign xor_ln1545_152_fu_8478_p2 = (xor_ln1545_153_fu_8472_p2 ^ xor_ln1545_151_fu_8466_p2);

assign xor_ln1545_153_fu_8472_p2 = (tmp_217_fu_8020_p4 ^ tmp_212_fu_7976_p4);

assign xor_ln1545_154_fu_8484_p2 = (trunc_ln674_49_fu_7938_p1 ^ tmp_205_fu_7918_p4);

assign xor_ln1545_155_fu_8496_p2 = (xor_ln1545_156_fu_8490_p2 ^ xor_ln1545_154_fu_8484_p2);

assign xor_ln1545_156_fu_8490_p2 = (tmp_216_fu_8010_p4 ^ tmp_214_fu_7996_p4);

assign xor_ln1545_157_fu_8502_p2 = (tmp_209_fu_7952_p4 ^ tmp_204_fu_7908_p4);

assign xor_ln1545_158_fu_8508_p2 = (trunc_ln674_50_fu_7972_p1 ^ tmp_218_fu_8030_p4);

assign xor_ln1545_160_fu_8520_p2 = (tmp_224_fu_8078_p4 ^ tmp_222_fu_8064_p4);

assign xor_ln1545_161_fu_8532_p2 = (xor_ln1545_162_fu_8526_p2 ^ xor_ln1545_160_fu_8520_p2);

assign xor_ln1545_162_fu_8526_p2 = (trunc_ln674_55_fu_8142_p1 ^ tmp_229_fu_8122_p4);

assign xor_ln1545_163_fu_8538_p2 = (trunc_ln674_52_fu_8040_p1 ^ tmp_226_fu_8098_p4);

assign xor_ln1545_164_fu_8550_p2 = (xor_ln1545_165_fu_8544_p2 ^ xor_ln1545_163_fu_8538_p2);

assign xor_ln1545_165_fu_8544_p2 = (tmp_233_fu_8156_p4 ^ tmp_228_fu_8112_p4);

assign xor_ln1545_166_fu_8556_p2 = (trunc_ln674_53_fu_8074_p1 ^ tmp_221_fu_8054_p4);

assign xor_ln1545_167_fu_8568_p2 = (xor_ln1545_168_fu_8562_p2 ^ xor_ln1545_166_fu_8556_p2);

assign xor_ln1545_168_fu_8562_p2 = (tmp_232_fu_8146_p4 ^ tmp_230_fu_8132_p4);

assign xor_ln1545_169_fu_8574_p2 = (tmp_225_fu_8088_p4 ^ tmp_220_fu_8044_p4);

assign xor_ln1545_16_fu_4959_p2 = (tmp_35_fu_4517_p4 ^ tmp_33_fu_4503_p4);

assign xor_ln1545_170_fu_8586_p2 = (xor_ln1545_171_fu_8580_p2 ^ xor_ln1545_169_fu_8574_p2);

assign xor_ln1545_171_fu_8580_p2 = (trunc_ln674_54_fu_8108_p1 ^ tmp_234_fu_8166_p4);

assign xor_ln1545_172_fu_8592_p2 = (tmp_240_fu_8214_p4 ^ tmp_238_fu_8200_p4);

assign xor_ln1545_173_fu_8604_p2 = (xor_ln1545_174_fu_8598_p2 ^ xor_ln1545_172_fu_8592_p2);

assign xor_ln1545_174_fu_8598_p2 = (trunc_ln674_59_fu_8278_p1 ^ tmp_245_fu_8258_p4);

assign xor_ln1545_175_fu_8610_p2 = (trunc_ln674_56_fu_8176_p1 ^ tmp_242_fu_8234_p4);

assign xor_ln1545_176_fu_8622_p2 = (xor_ln1545_177_fu_8616_p2 ^ xor_ln1545_175_fu_8610_p2);

assign xor_ln1545_177_fu_8616_p2 = (tmp_249_fu_8292_p4 ^ tmp_244_fu_8248_p4);

assign xor_ln1545_178_fu_8628_p2 = (trunc_ln674_57_fu_8210_p1 ^ tmp_237_fu_8190_p4);

assign xor_ln1545_179_fu_8634_p2 = (tmp_248_fu_8282_p4 ^ tmp_246_fu_8268_p4);

assign xor_ln1545_17_fu_4971_p2 = (xor_ln1545_18_fu_4965_p2 ^ xor_ln1545_16_fu_4959_p2);

assign xor_ln1545_181_fu_8646_p2 = (tmp_241_fu_8224_p4 ^ tmp_236_fu_8180_p4);

assign xor_ln1545_182_fu_8658_p2 = (xor_ln1545_183_fu_8652_p2 ^ xor_ln1545_181_fu_8646_p2);

assign xor_ln1545_183_fu_8652_p2 = (trunc_ln674_58_fu_8244_p1 ^ tmp_250_fu_8302_p4);

assign xor_ln1545_184_fu_8664_p2 = (tmp_256_fu_8350_p4 ^ tmp_254_fu_8336_p4);

assign xor_ln1545_185_fu_8676_p2 = (xor_ln1545_186_fu_8670_p2 ^ xor_ln1545_184_fu_8664_p2);

assign xor_ln1545_186_fu_8670_p2 = (trunc_ln674_63_fu_8414_p1 ^ tmp_261_fu_8394_p4);

assign xor_ln1545_187_fu_8682_p2 = (trunc_ln674_60_fu_8312_p1 ^ tmp_258_fu_8370_p4);

assign xor_ln1545_188_fu_8688_p2 = (tmp_265_fu_8428_p4 ^ tmp_260_fu_8384_p4);

assign xor_ln1545_18_fu_4965_p2 = (trunc_ln674_7_fu_4581_p1 ^ tmp_40_fu_4561_p4);

assign xor_ln1545_190_fu_8700_p2 = (trunc_ln674_61_fu_8346_p1 ^ tmp_253_fu_8326_p4);

assign xor_ln1545_191_fu_8706_p2 = (tmp_264_fu_8418_p4 ^ tmp_262_fu_8404_p4);

assign xor_ln1545_193_fu_8718_p2 = (tmp_257_fu_8360_p4 ^ tmp_252_fu_8316_p4);

assign xor_ln1545_194_fu_8730_p2 = (xor_ln1545_195_fu_8724_p2 ^ xor_ln1545_193_fu_8718_p2);

assign xor_ln1545_195_fu_8724_p2 = (trunc_ln674_62_fu_8380_p1 ^ tmp_266_fu_8438_p4);

assign xor_ln1545_196_fu_9635_p2 = (tmp_271_fu_9129_p4 ^ tmp_269_fu_9115_p4);

assign xor_ln1545_197_fu_9647_p2 = (xor_ln1545_198_fu_9641_p2 ^ xor_ln1545_196_fu_9635_p2);

assign xor_ln1545_198_fu_9641_p2 = (trunc_ln674_67_fu_9193_p1 ^ tmp_276_fu_9173_p4);

assign xor_ln1545_199_fu_9653_p2 = (trunc_ln674_64_fu_9091_p1 ^ tmp_273_fu_9149_p4);

assign xor_ln1545_19_fu_4977_p2 = (trunc_ln674_4_fu_4479_p1 ^ tmp_37_fu_4537_p4);

assign xor_ln1545_200_fu_9665_p2 = (xor_ln1545_201_fu_9659_p2 ^ xor_ln1545_199_fu_9653_p2);

assign xor_ln1545_201_fu_9659_p2 = (tmp_280_fu_9207_p4 ^ tmp_275_fu_9163_p4);

assign xor_ln1545_202_fu_9671_p2 = (trunc_ln674_65_fu_9125_p1 ^ tmp_268_fu_9105_p4);

assign xor_ln1545_203_fu_9683_p2 = (xor_ln1545_204_fu_9677_p2 ^ xor_ln1545_202_fu_9671_p2);

assign xor_ln1545_204_fu_9677_p2 = (tmp_279_fu_9197_p4 ^ tmp_277_fu_9183_p4);

assign xor_ln1545_205_fu_9689_p2 = (tmp_272_fu_9139_p4 ^ tmp_267_fu_9095_p4);

assign xor_ln1545_206_fu_9695_p2 = (trunc_ln674_66_fu_9159_p1 ^ tmp_281_fu_9217_p4);

assign xor_ln1545_208_fu_9707_p2 = (tmp_287_fu_9265_p4 ^ tmp_285_fu_9251_p4);

assign xor_ln1545_209_fu_9719_p2 = (xor_ln1545_210_fu_9713_p2 ^ xor_ln1545_208_fu_9707_p2);

assign xor_ln1545_20_fu_4989_p2 = (xor_ln1545_21_fu_4983_p2 ^ xor_ln1545_19_fu_4977_p2);

assign xor_ln1545_210_fu_9713_p2 = (trunc_ln674_71_fu_9329_p1 ^ tmp_292_fu_9309_p4);

assign xor_ln1545_211_fu_9725_p2 = (trunc_ln674_68_fu_9227_p1 ^ tmp_289_fu_9285_p4);

assign xor_ln1545_212_fu_9737_p2 = (xor_ln1545_213_fu_9731_p2 ^ xor_ln1545_211_fu_9725_p2);

assign xor_ln1545_213_fu_9731_p2 = (tmp_296_fu_9343_p4 ^ tmp_291_fu_9299_p4);

assign xor_ln1545_214_fu_9743_p2 = (trunc_ln674_69_fu_9261_p1 ^ tmp_284_fu_9241_p4);

assign xor_ln1545_215_fu_9755_p2 = (xor_ln1545_216_fu_9749_p2 ^ xor_ln1545_214_fu_9743_p2);

assign xor_ln1545_216_fu_9749_p2 = (tmp_295_fu_9333_p4 ^ tmp_293_fu_9319_p4);

assign xor_ln1545_217_fu_9761_p2 = (tmp_288_fu_9275_p4 ^ tmp_283_fu_9231_p4);

assign xor_ln1545_218_fu_9773_p2 = (xor_ln1545_219_fu_9767_p2 ^ xor_ln1545_217_fu_9761_p2);

assign xor_ln1545_219_fu_9767_p2 = (trunc_ln674_70_fu_9295_p1 ^ tmp_297_fu_9353_p4);

assign xor_ln1545_21_fu_4983_p2 = (tmp_44_fu_4595_p4 ^ tmp_39_fu_4551_p4);

assign xor_ln1545_220_fu_9779_p2 = (tmp_303_fu_9401_p4 ^ tmp_301_fu_9387_p4);

assign xor_ln1545_221_fu_9791_p2 = (xor_ln1545_222_fu_9785_p2 ^ xor_ln1545_220_fu_9779_p2);

assign xor_ln1545_222_fu_9785_p2 = (trunc_ln674_75_fu_9465_p1 ^ tmp_308_fu_9445_p4);

assign xor_ln1545_223_fu_9797_p2 = (trunc_ln674_72_fu_9363_p1 ^ tmp_305_fu_9421_p4);

assign xor_ln1545_224_fu_9809_p2 = (xor_ln1545_225_fu_9803_p2 ^ xor_ln1545_223_fu_9797_p2);

assign xor_ln1545_225_fu_9803_p2 = (tmp_312_fu_9479_p4 ^ tmp_307_fu_9435_p4);

assign xor_ln1545_226_fu_9815_p2 = (trunc_ln674_73_fu_9397_p1 ^ tmp_300_fu_9377_p4);

assign xor_ln1545_227_fu_9821_p2 = (tmp_311_fu_9469_p4 ^ tmp_309_fu_9455_p4);

assign xor_ln1545_229_fu_9833_p2 = (tmp_304_fu_9411_p4 ^ tmp_299_fu_9367_p4);

assign xor_ln1545_22_fu_4995_p2 = (trunc_ln674_5_fu_4513_p1 ^ tmp_32_fu_4493_p4);

assign xor_ln1545_230_fu_9845_p2 = (xor_ln1545_231_fu_9839_p2 ^ xor_ln1545_229_fu_9833_p2);

assign xor_ln1545_231_fu_9839_p2 = (trunc_ln674_74_fu_9431_p1 ^ tmp_313_fu_9489_p4);

assign xor_ln1545_232_fu_9851_p2 = (tmp_319_fu_9537_p4 ^ tmp_317_fu_9523_p4);

assign xor_ln1545_233_fu_9863_p2 = (xor_ln1545_234_fu_9857_p2 ^ xor_ln1545_232_fu_9851_p2);

assign xor_ln1545_234_fu_9857_p2 = (trunc_ln674_79_fu_9601_p1 ^ tmp_324_fu_9581_p4);

assign xor_ln1545_235_fu_9869_p2 = (trunc_ln674_76_fu_9499_p1 ^ tmp_321_fu_9557_p4);

assign xor_ln1545_236_fu_9875_p2 = (tmp_328_fu_9615_p4 ^ tmp_323_fu_9571_p4);

assign xor_ln1545_238_fu_9887_p2 = (trunc_ln674_77_fu_9533_p1 ^ tmp_316_fu_9513_p4);

assign xor_ln1545_239_fu_9893_p2 = (tmp_327_fu_9605_p4 ^ tmp_325_fu_9591_p4);

assign xor_ln1545_23_fu_5007_p2 = (xor_ln1545_24_fu_5001_p2 ^ xor_ln1545_22_fu_4995_p2);

assign xor_ln1545_241_fu_9905_p2 = (tmp_320_fu_9547_p4 ^ tmp_315_fu_9503_p4);

assign xor_ln1545_242_fu_9917_p2 = (xor_ln1545_243_fu_9911_p2 ^ xor_ln1545_241_fu_9905_p2);

assign xor_ln1545_243_fu_9911_p2 = (trunc_ln674_78_fu_9567_p1 ^ tmp_329_fu_9625_p4);

assign xor_ln1545_244_fu_10822_p2 = (tmp_334_fu_10316_p4 ^ tmp_332_fu_10302_p4);

assign xor_ln1545_245_fu_10834_p2 = (xor_ln1545_246_fu_10828_p2 ^ xor_ln1545_244_fu_10822_p2);

assign xor_ln1545_246_fu_10828_p2 = (trunc_ln674_83_fu_10380_p1 ^ tmp_339_fu_10360_p4);

assign xor_ln1545_247_fu_10840_p2 = (trunc_ln674_80_fu_10278_p1 ^ tmp_336_fu_10336_p4);

assign xor_ln1545_248_fu_10852_p2 = (xor_ln1545_249_fu_10846_p2 ^ xor_ln1545_247_fu_10840_p2);

assign xor_ln1545_249_fu_10846_p2 = (tmp_343_fu_10394_p4 ^ tmp_338_fu_10350_p4);

assign xor_ln1545_24_fu_5001_p2 = (tmp_43_fu_4585_p4 ^ tmp_41_fu_4571_p4);

assign xor_ln1545_250_fu_10858_p2 = (trunc_ln674_81_fu_10312_p1 ^ tmp_331_fu_10292_p4);

assign xor_ln1545_251_fu_10870_p2 = (xor_ln1545_252_fu_10864_p2 ^ xor_ln1545_250_fu_10858_p2);

assign xor_ln1545_252_fu_10864_p2 = (tmp_342_fu_10384_p4 ^ tmp_340_fu_10370_p4);

assign xor_ln1545_253_fu_10876_p2 = (tmp_335_fu_10326_p4 ^ tmp_330_fu_10282_p4);

assign xor_ln1545_254_fu_10882_p2 = (trunc_ln674_82_fu_10346_p1 ^ tmp_344_fu_10404_p4);

assign xor_ln1545_256_fu_10894_p2 = (tmp_350_fu_10452_p4 ^ tmp_348_fu_10438_p4);

assign xor_ln1545_257_fu_10906_p2 = (xor_ln1545_258_fu_10900_p2 ^ xor_ln1545_256_fu_10894_p2);

assign xor_ln1545_258_fu_10900_p2 = (trunc_ln674_87_fu_10516_p1 ^ tmp_355_fu_10496_p4);

assign xor_ln1545_259_fu_10912_p2 = (trunc_ln674_84_fu_10414_p1 ^ tmp_352_fu_10472_p4);

assign xor_ln1545_25_fu_5013_p2 = (tmp_36_fu_4527_p4 ^ tmp_31_fu_4483_p4);

assign xor_ln1545_260_fu_10924_p2 = (xor_ln1545_261_fu_10918_p2 ^ xor_ln1545_259_fu_10912_p2);

assign xor_ln1545_261_fu_10918_p2 = (tmp_359_fu_10530_p4 ^ tmp_354_fu_10486_p4);

assign xor_ln1545_262_fu_10930_p2 = (trunc_ln674_85_fu_10448_p1 ^ tmp_347_fu_10428_p4);

assign xor_ln1545_263_fu_10942_p2 = (xor_ln1545_264_fu_10936_p2 ^ xor_ln1545_262_fu_10930_p2);

assign xor_ln1545_264_fu_10936_p2 = (tmp_358_fu_10520_p4 ^ tmp_356_fu_10506_p4);

assign xor_ln1545_265_fu_10948_p2 = (tmp_351_fu_10462_p4 ^ tmp_346_fu_10418_p4);

assign xor_ln1545_266_fu_10960_p2 = (xor_ln1545_267_fu_10954_p2 ^ xor_ln1545_265_fu_10948_p2);

assign xor_ln1545_267_fu_10954_p2 = (trunc_ln674_86_fu_10482_p1 ^ tmp_360_fu_10540_p4);

assign xor_ln1545_268_fu_10966_p2 = (tmp_366_fu_10588_p4 ^ tmp_364_fu_10574_p4);

assign xor_ln1545_269_fu_10978_p2 = (xor_ln1545_270_fu_10972_p2 ^ xor_ln1545_268_fu_10966_p2);

assign xor_ln1545_26_fu_5025_p2 = (xor_ln1545_27_fu_5019_p2 ^ xor_ln1545_25_fu_5013_p2);

assign xor_ln1545_270_fu_10972_p2 = (trunc_ln674_91_fu_10652_p1 ^ tmp_371_fu_10632_p4);

assign xor_ln1545_271_fu_10984_p2 = (trunc_ln674_88_fu_10550_p1 ^ tmp_368_fu_10608_p4);

assign xor_ln1545_272_fu_10996_p2 = (xor_ln1545_273_fu_10990_p2 ^ xor_ln1545_271_fu_10984_p2);

assign xor_ln1545_273_fu_10990_p2 = (tmp_375_fu_10666_p4 ^ tmp_370_fu_10622_p4);

assign xor_ln1545_274_fu_11002_p2 = (trunc_ln674_89_fu_10584_p1 ^ tmp_363_fu_10564_p4);

assign xor_ln1545_275_fu_11008_p2 = (tmp_374_fu_10656_p4 ^ tmp_372_fu_10642_p4);

assign xor_ln1545_277_fu_11020_p2 = (tmp_367_fu_10598_p4 ^ tmp_362_fu_10554_p4);

assign xor_ln1545_278_fu_11032_p2 = (xor_ln1545_279_fu_11026_p2 ^ xor_ln1545_277_fu_11020_p2);

assign xor_ln1545_279_fu_11026_p2 = (trunc_ln674_90_fu_10618_p1 ^ tmp_376_fu_10676_p4);

assign xor_ln1545_27_fu_5019_p2 = (trunc_ln674_6_fu_4547_p1 ^ tmp_45_fu_4605_p4);

assign xor_ln1545_280_fu_11038_p2 = (tmp_382_fu_10724_p4 ^ tmp_380_fu_10710_p4);

assign xor_ln1545_281_fu_11050_p2 = (xor_ln1545_282_fu_11044_p2 ^ xor_ln1545_280_fu_11038_p2);

assign xor_ln1545_282_fu_11044_p2 = (trunc_ln674_95_fu_10788_p1 ^ tmp_387_fu_10768_p4);

assign xor_ln1545_283_fu_11056_p2 = (trunc_ln674_92_fu_10686_p1 ^ tmp_384_fu_10744_p4);

assign xor_ln1545_284_fu_11062_p2 = (tmp_391_fu_10802_p4 ^ tmp_386_fu_10758_p4);

assign xor_ln1545_286_fu_11074_p2 = (trunc_ln674_93_fu_10720_p1 ^ tmp_379_fu_10700_p4);

assign xor_ln1545_287_fu_11080_p2 = (tmp_390_fu_10792_p4 ^ tmp_388_fu_10778_p4);

assign xor_ln1545_289_fu_11092_p2 = (tmp_383_fu_10734_p4 ^ tmp_378_fu_10690_p4);

assign xor_ln1545_28_fu_5031_p2 = (tmp_51_fu_4653_p4 ^ tmp_49_fu_4639_p4);

assign xor_ln1545_290_fu_11104_p2 = (xor_ln1545_291_fu_11098_p2 ^ xor_ln1545_289_fu_11092_p2);

assign xor_ln1545_291_fu_11098_p2 = (trunc_ln674_94_fu_10754_p1 ^ tmp_392_fu_10812_p4);

assign xor_ln1545_292_fu_12009_p2 = (tmp_397_fu_11503_p4 ^ tmp_395_fu_11489_p4);

assign xor_ln1545_293_fu_12021_p2 = (xor_ln1545_294_fu_12015_p2 ^ xor_ln1545_292_fu_12009_p2);

assign xor_ln1545_294_fu_12015_p2 = (trunc_ln674_99_fu_11567_p1 ^ tmp_402_fu_11547_p4);

assign xor_ln1545_295_fu_12027_p2 = (trunc_ln674_96_fu_11465_p1 ^ tmp_399_fu_11523_p4);

assign xor_ln1545_296_fu_12039_p2 = (xor_ln1545_297_fu_12033_p2 ^ xor_ln1545_295_fu_12027_p2);

assign xor_ln1545_297_fu_12033_p2 = (tmp_406_fu_11581_p4 ^ tmp_401_fu_11537_p4);

assign xor_ln1545_298_fu_12045_p2 = (trunc_ln674_97_fu_11499_p1 ^ tmp_394_fu_11479_p4);

assign xor_ln1545_299_fu_12057_p2 = (xor_ln1545_300_fu_12051_p2 ^ xor_ln1545_298_fu_12045_p2);

assign xor_ln1545_29_fu_5043_p2 = (xor_ln1545_30_fu_5037_p2 ^ xor_ln1545_28_fu_5031_p2);

assign xor_ln1545_300_fu_12051_p2 = (tmp_405_fu_11571_p4 ^ tmp_403_fu_11557_p4);

assign xor_ln1545_301_fu_12063_p2 = (tmp_398_fu_11513_p4 ^ tmp_393_fu_11469_p4);

assign xor_ln1545_302_fu_12069_p2 = (trunc_ln674_98_fu_11533_p1 ^ tmp_407_fu_11591_p4);

assign xor_ln1545_304_fu_12081_p2 = (tmp_413_fu_11639_p4 ^ tmp_411_fu_11625_p4);

assign xor_ln1545_305_fu_12093_p2 = (xor_ln1545_306_fu_12087_p2 ^ xor_ln1545_304_fu_12081_p2);

assign xor_ln1545_306_fu_12087_p2 = (trunc_ln674_103_fu_11703_p1 ^ tmp_418_fu_11683_p4);

assign xor_ln1545_307_fu_12099_p2 = (trunc_ln674_100_fu_11601_p1 ^ tmp_415_fu_11659_p4);

assign xor_ln1545_308_fu_12111_p2 = (xor_ln1545_309_fu_12105_p2 ^ xor_ln1545_307_fu_12099_p2);

assign xor_ln1545_309_fu_12105_p2 = (tmp_422_fu_11717_p4 ^ tmp_417_fu_11673_p4);

assign xor_ln1545_30_fu_5037_p2 = (trunc_ln674_11_fu_4717_p1 ^ tmp_56_fu_4697_p4);

assign xor_ln1545_310_fu_12117_p2 = (trunc_ln674_101_fu_11635_p1 ^ tmp_410_fu_11615_p4);

assign xor_ln1545_311_fu_12129_p2 = (xor_ln1545_312_fu_12123_p2 ^ xor_ln1545_310_fu_12117_p2);

assign xor_ln1545_312_fu_12123_p2 = (tmp_421_fu_11707_p4 ^ tmp_419_fu_11693_p4);

assign xor_ln1545_313_fu_12135_p2 = (tmp_414_fu_11649_p4 ^ tmp_409_fu_11605_p4);

assign xor_ln1545_314_fu_12147_p2 = (xor_ln1545_315_fu_12141_p2 ^ xor_ln1545_313_fu_12135_p2);

assign xor_ln1545_315_fu_12141_p2 = (trunc_ln674_102_fu_11669_p1 ^ tmp_423_fu_11727_p4);

assign xor_ln1545_316_fu_12153_p2 = (tmp_429_fu_11775_p4 ^ tmp_427_fu_11761_p4);

assign xor_ln1545_317_fu_12165_p2 = (xor_ln1545_318_fu_12159_p2 ^ xor_ln1545_316_fu_12153_p2);

assign xor_ln1545_318_fu_12159_p2 = (trunc_ln674_107_fu_11839_p1 ^ tmp_434_fu_11819_p4);

assign xor_ln1545_319_fu_12171_p2 = (trunc_ln674_104_fu_11737_p1 ^ tmp_431_fu_11795_p4);

assign xor_ln1545_31_fu_5049_p2 = (trunc_ln674_8_fu_4615_p1 ^ tmp_53_fu_4673_p4);

assign xor_ln1545_320_fu_12183_p2 = (xor_ln1545_321_fu_12177_p2 ^ xor_ln1545_319_fu_12171_p2);

assign xor_ln1545_321_fu_12177_p2 = (tmp_438_fu_11853_p4 ^ tmp_433_fu_11809_p4);

assign xor_ln1545_322_fu_12189_p2 = (trunc_ln674_105_fu_11771_p1 ^ tmp_426_fu_11751_p4);

assign xor_ln1545_323_fu_12195_p2 = (tmp_437_fu_11843_p4 ^ tmp_435_fu_11829_p4);

assign xor_ln1545_325_fu_12207_p2 = (tmp_430_fu_11785_p4 ^ tmp_425_fu_11741_p4);

assign xor_ln1545_326_fu_12219_p2 = (xor_ln1545_327_fu_12213_p2 ^ xor_ln1545_325_fu_12207_p2);

assign xor_ln1545_327_fu_12213_p2 = (trunc_ln674_106_fu_11805_p1 ^ tmp_439_fu_11863_p4);

assign xor_ln1545_328_fu_12225_p2 = (tmp_445_fu_11911_p4 ^ tmp_443_fu_11897_p4);

assign xor_ln1545_329_fu_12237_p2 = (xor_ln1545_330_fu_12231_p2 ^ xor_ln1545_328_fu_12225_p2);

assign xor_ln1545_32_fu_5061_p2 = (xor_ln1545_33_fu_5055_p2 ^ xor_ln1545_31_fu_5049_p2);

assign xor_ln1545_330_fu_12231_p2 = (trunc_ln674_111_fu_11975_p1 ^ tmp_450_fu_11955_p4);

assign xor_ln1545_331_fu_12243_p2 = (trunc_ln674_108_fu_11873_p1 ^ tmp_447_fu_11931_p4);

assign xor_ln1545_332_fu_12249_p2 = (tmp_454_fu_11989_p4 ^ tmp_449_fu_11945_p4);

assign xor_ln1545_334_fu_12261_p2 = (trunc_ln674_109_fu_11907_p1 ^ tmp_442_fu_11887_p4);

assign xor_ln1545_335_fu_12267_p2 = (tmp_453_fu_11979_p4 ^ tmp_451_fu_11965_p4);

assign xor_ln1545_337_fu_12279_p2 = (tmp_446_fu_11921_p4 ^ tmp_441_fu_11877_p4);

assign xor_ln1545_338_fu_12291_p2 = (xor_ln1545_339_fu_12285_p2 ^ xor_ln1545_337_fu_12279_p2);

assign xor_ln1545_339_fu_12285_p2 = (trunc_ln674_110_fu_11941_p1 ^ tmp_455_fu_11999_p4);

assign xor_ln1545_33_fu_5055_p2 = (tmp_60_fu_4731_p4 ^ tmp_55_fu_4687_p4);

assign xor_ln1545_340_fu_13196_p2 = (tmp_460_fu_12690_p4 ^ tmp_458_fu_12676_p4);

assign xor_ln1545_341_fu_13208_p2 = (xor_ln1545_342_fu_13202_p2 ^ xor_ln1545_340_fu_13196_p2);

assign xor_ln1545_342_fu_13202_p2 = (trunc_ln674_115_fu_12754_p1 ^ tmp_465_fu_12734_p4);

assign xor_ln1545_343_fu_13214_p2 = (trunc_ln674_112_fu_12652_p1 ^ tmp_462_fu_12710_p4);

assign xor_ln1545_344_fu_13226_p2 = (xor_ln1545_345_fu_13220_p2 ^ xor_ln1545_343_fu_13214_p2);

assign xor_ln1545_345_fu_13220_p2 = (tmp_469_fu_12768_p4 ^ tmp_464_fu_12724_p4);

assign xor_ln1545_346_fu_13232_p2 = (trunc_ln674_113_fu_12686_p1 ^ tmp_457_fu_12666_p4);

assign xor_ln1545_347_fu_13244_p2 = (xor_ln1545_348_fu_13238_p2 ^ xor_ln1545_346_fu_13232_p2);

assign xor_ln1545_348_fu_13238_p2 = (tmp_468_fu_12758_p4 ^ tmp_466_fu_12744_p4);

assign xor_ln1545_349_fu_13250_p2 = (tmp_461_fu_12700_p4 ^ tmp_456_fu_12656_p4);

assign xor_ln1545_34_fu_5067_p2 = (trunc_ln674_9_fu_4649_p1 ^ tmp_48_fu_4629_p4);

assign xor_ln1545_350_fu_13256_p2 = (trunc_ln674_114_fu_12720_p1 ^ tmp_470_fu_12778_p4);

assign xor_ln1545_352_fu_13268_p2 = (tmp_476_fu_12826_p4 ^ tmp_474_fu_12812_p4);

assign xor_ln1545_353_fu_13280_p2 = (xor_ln1545_354_fu_13274_p2 ^ xor_ln1545_352_fu_13268_p2);

assign xor_ln1545_354_fu_13274_p2 = (trunc_ln674_119_fu_12890_p1 ^ tmp_481_fu_12870_p4);

assign xor_ln1545_355_fu_13286_p2 = (trunc_ln674_116_fu_12788_p1 ^ tmp_478_fu_12846_p4);

assign xor_ln1545_356_fu_13298_p2 = (xor_ln1545_357_fu_13292_p2 ^ xor_ln1545_355_fu_13286_p2);

assign xor_ln1545_357_fu_13292_p2 = (tmp_485_fu_12904_p4 ^ tmp_480_fu_12860_p4);

assign xor_ln1545_358_fu_13304_p2 = (trunc_ln674_117_fu_12822_p1 ^ tmp_473_fu_12802_p4);

assign xor_ln1545_359_fu_13316_p2 = (xor_ln1545_360_fu_13310_p2 ^ xor_ln1545_358_fu_13304_p2);

assign xor_ln1545_35_fu_5073_p2 = (tmp_59_fu_4721_p4 ^ tmp_57_fu_4707_p4);

assign xor_ln1545_360_fu_13310_p2 = (tmp_484_fu_12894_p4 ^ tmp_482_fu_12880_p4);

assign xor_ln1545_361_fu_13322_p2 = (tmp_477_fu_12836_p4 ^ tmp_472_fu_12792_p4);

assign xor_ln1545_362_fu_13334_p2 = (xor_ln1545_363_fu_13328_p2 ^ xor_ln1545_361_fu_13322_p2);

assign xor_ln1545_363_fu_13328_p2 = (trunc_ln674_118_fu_12856_p1 ^ tmp_486_fu_12914_p4);

assign xor_ln1545_364_fu_13340_p2 = (tmp_492_fu_12962_p4 ^ tmp_490_fu_12948_p4);

assign xor_ln1545_365_fu_13352_p2 = (xor_ln1545_366_fu_13346_p2 ^ xor_ln1545_364_fu_13340_p2);

assign xor_ln1545_366_fu_13346_p2 = (trunc_ln674_123_fu_13026_p1 ^ tmp_497_fu_13006_p4);

assign xor_ln1545_367_fu_13358_p2 = (trunc_ln674_120_fu_12924_p1 ^ tmp_494_fu_12982_p4);

assign xor_ln1545_368_fu_13370_p2 = (xor_ln1545_369_fu_13364_p2 ^ xor_ln1545_367_fu_13358_p2);

assign xor_ln1545_369_fu_13364_p2 = (tmp_501_fu_13040_p4 ^ tmp_496_fu_12996_p4);

assign xor_ln1545_370_fu_13376_p2 = (trunc_ln674_121_fu_12958_p1 ^ tmp_489_fu_12938_p4);

assign xor_ln1545_371_fu_13382_p2 = (tmp_500_fu_13030_p4 ^ tmp_498_fu_13016_p4);

assign xor_ln1545_373_fu_13394_p2 = (tmp_493_fu_12972_p4 ^ tmp_488_fu_12928_p4);

assign xor_ln1545_374_fu_13406_p2 = (xor_ln1545_375_fu_13400_p2 ^ xor_ln1545_373_fu_13394_p2);

assign xor_ln1545_375_fu_13400_p2 = (trunc_ln674_122_fu_12992_p1 ^ tmp_502_fu_13050_p4);

assign xor_ln1545_376_fu_13412_p2 = (tmp_508_fu_13098_p4 ^ tmp_506_fu_13084_p4);

assign xor_ln1545_377_fu_13424_p2 = (xor_ln1545_378_fu_13418_p2 ^ xor_ln1545_376_fu_13412_p2);

assign xor_ln1545_378_fu_13418_p2 = (trunc_ln674_127_fu_13162_p1 ^ tmp_513_fu_13142_p4);

assign xor_ln1545_379_fu_13430_p2 = (trunc_ln674_124_fu_13060_p1 ^ tmp_510_fu_13118_p4);

assign xor_ln1545_37_fu_5085_p2 = (tmp_52_fu_4663_p4 ^ tmp_47_fu_4619_p4);

assign xor_ln1545_380_fu_13436_p2 = (tmp_517_fu_13176_p4 ^ tmp_512_fu_13132_p4);

assign xor_ln1545_382_fu_13448_p2 = (trunc_ln674_125_fu_13094_p1 ^ tmp_505_fu_13074_p4);

assign xor_ln1545_383_fu_13454_p2 = (tmp_516_fu_13166_p4 ^ tmp_514_fu_13152_p4);

assign xor_ln1545_385_fu_13466_p2 = (tmp_509_fu_13108_p4 ^ tmp_504_fu_13064_p4);

assign xor_ln1545_386_fu_13478_p2 = (xor_ln1545_387_fu_13472_p2 ^ xor_ln1545_385_fu_13466_p2);

assign xor_ln1545_387_fu_13472_p2 = (trunc_ln674_126_fu_13128_p1 ^ tmp_518_fu_13186_p4);

assign xor_ln1545_388_fu_14383_p2 = (tmp_523_fu_13877_p4 ^ tmp_521_fu_13863_p4);

assign xor_ln1545_389_fu_14395_p2 = (xor_ln1545_390_fu_14389_p2 ^ xor_ln1545_388_fu_14383_p2);

assign xor_ln1545_38_fu_5097_p2 = (xor_ln1545_39_fu_5091_p2 ^ xor_ln1545_37_fu_5085_p2);

assign xor_ln1545_390_fu_14389_p2 = (trunc_ln674_131_fu_13941_p1 ^ tmp_528_fu_13921_p4);

assign xor_ln1545_391_fu_14401_p2 = (trunc_ln674_128_fu_13839_p1 ^ tmp_525_fu_13897_p4);

assign xor_ln1545_392_fu_14413_p2 = (xor_ln1545_393_fu_14407_p2 ^ xor_ln1545_391_fu_14401_p2);

assign xor_ln1545_393_fu_14407_p2 = (tmp_532_fu_13955_p4 ^ tmp_527_fu_13911_p4);

assign xor_ln1545_394_fu_14419_p2 = (trunc_ln674_129_fu_13873_p1 ^ tmp_520_fu_13853_p4);

assign xor_ln1545_395_fu_14431_p2 = (xor_ln1545_396_fu_14425_p2 ^ xor_ln1545_394_fu_14419_p2);

assign xor_ln1545_396_fu_14425_p2 = (tmp_531_fu_13945_p4 ^ tmp_529_fu_13931_p4);

assign xor_ln1545_397_fu_14437_p2 = (tmp_524_fu_13887_p4 ^ tmp_519_fu_13843_p4);

assign xor_ln1545_398_fu_14443_p2 = (trunc_ln674_130_fu_13907_p1 ^ tmp_533_fu_13965_p4);

assign xor_ln1545_39_fu_5091_p2 = (trunc_ln674_10_fu_4683_p1 ^ tmp_61_fu_4741_p4);

assign xor_ln1545_400_fu_14455_p2 = (tmp_539_fu_14013_p4 ^ tmp_537_fu_13999_p4);

assign xor_ln1545_401_fu_14467_p2 = (xor_ln1545_402_fu_14461_p2 ^ xor_ln1545_400_fu_14455_p2);

assign xor_ln1545_402_fu_14461_p2 = (trunc_ln674_135_fu_14077_p1 ^ tmp_544_fu_14057_p4);

assign xor_ln1545_403_fu_14473_p2 = (trunc_ln674_132_fu_13975_p1 ^ tmp_541_fu_14033_p4);

assign xor_ln1545_404_fu_14485_p2 = (xor_ln1545_405_fu_14479_p2 ^ xor_ln1545_403_fu_14473_p2);

assign xor_ln1545_405_fu_14479_p2 = (tmp_548_fu_14091_p4 ^ tmp_543_fu_14047_p4);

assign xor_ln1545_406_fu_14491_p2 = (trunc_ln674_133_fu_14009_p1 ^ tmp_536_fu_13989_p4);

assign xor_ln1545_407_fu_14503_p2 = (xor_ln1545_408_fu_14497_p2 ^ xor_ln1545_406_fu_14491_p2);

assign xor_ln1545_408_fu_14497_p2 = (tmp_547_fu_14081_p4 ^ tmp_545_fu_14067_p4);

assign xor_ln1545_409_fu_14509_p2 = (tmp_540_fu_14023_p4 ^ tmp_535_fu_13979_p4);

assign xor_ln1545_40_fu_5103_p2 = (tmp_67_fu_4789_p4 ^ tmp_65_fu_4775_p4);

assign xor_ln1545_410_fu_14521_p2 = (xor_ln1545_411_fu_14515_p2 ^ xor_ln1545_409_fu_14509_p2);

assign xor_ln1545_411_fu_14515_p2 = (trunc_ln674_134_fu_14043_p1 ^ tmp_549_fu_14101_p4);

assign xor_ln1545_412_fu_14527_p2 = (tmp_555_fu_14149_p4 ^ tmp_553_fu_14135_p4);

assign xor_ln1545_413_fu_14539_p2 = (xor_ln1545_414_fu_14533_p2 ^ xor_ln1545_412_fu_14527_p2);

assign xor_ln1545_414_fu_14533_p2 = (trunc_ln674_139_fu_14213_p1 ^ tmp_560_fu_14193_p4);

assign xor_ln1545_415_fu_14545_p2 = (trunc_ln674_136_fu_14111_p1 ^ tmp_557_fu_14169_p4);

assign xor_ln1545_416_fu_14557_p2 = (xor_ln1545_417_fu_14551_p2 ^ xor_ln1545_415_fu_14545_p2);

assign xor_ln1545_417_fu_14551_p2 = (tmp_564_fu_14227_p4 ^ tmp_559_fu_14183_p4);

assign xor_ln1545_418_fu_14563_p2 = (trunc_ln674_137_fu_14145_p1 ^ tmp_552_fu_14125_p4);

assign xor_ln1545_419_fu_14569_p2 = (tmp_563_fu_14217_p4 ^ tmp_561_fu_14203_p4);

assign xor_ln1545_41_fu_5115_p2 = (xor_ln1545_42_fu_5109_p2 ^ xor_ln1545_40_fu_5103_p2);

assign xor_ln1545_421_fu_14581_p2 = (tmp_556_fu_14159_p4 ^ tmp_551_fu_14115_p4);

assign xor_ln1545_422_fu_14593_p2 = (xor_ln1545_423_fu_14587_p2 ^ xor_ln1545_421_fu_14581_p2);

assign xor_ln1545_423_fu_14587_p2 = (trunc_ln674_138_fu_14179_p1 ^ tmp_565_fu_14237_p4);

assign xor_ln1545_424_fu_14599_p2 = (tmp_571_fu_14285_p4 ^ tmp_569_fu_14271_p4);

assign xor_ln1545_425_fu_14611_p2 = (xor_ln1545_426_fu_14605_p2 ^ xor_ln1545_424_fu_14599_p2);

assign xor_ln1545_426_fu_14605_p2 = (trunc_ln674_143_fu_14349_p1 ^ tmp_576_fu_14329_p4);

assign xor_ln1545_427_fu_14617_p2 = (trunc_ln674_140_fu_14247_p1 ^ tmp_573_fu_14305_p4);

assign xor_ln1545_428_fu_14623_p2 = (tmp_580_fu_14363_p4 ^ tmp_575_fu_14319_p4);

assign xor_ln1545_42_fu_5109_p2 = (trunc_ln674_15_fu_4853_p1 ^ tmp_72_fu_4833_p4);

assign xor_ln1545_430_fu_14635_p2 = (trunc_ln674_141_fu_14281_p1 ^ tmp_568_fu_14261_p4);

assign xor_ln1545_431_fu_14641_p2 = (tmp_579_fu_14353_p4 ^ tmp_577_fu_14339_p4);

assign xor_ln1545_433_fu_14653_p2 = (tmp_572_fu_14295_p4 ^ tmp_567_fu_14251_p4);

assign xor_ln1545_434_fu_14665_p2 = (xor_ln1545_435_fu_14659_p2 ^ xor_ln1545_433_fu_14653_p2);

assign xor_ln1545_435_fu_14659_p2 = (trunc_ln674_142_fu_14315_p1 ^ tmp_581_fu_14373_p4);

assign xor_ln1545_43_fu_5121_p2 = (trunc_ln674_12_fu_4751_p1 ^ tmp_69_fu_4809_p4);

assign xor_ln1545_44_fu_5127_p2 = (tmp_76_fu_4867_p4 ^ tmp_71_fu_4823_p4);

assign xor_ln1545_46_fu_5139_p2 = (trunc_ln674_13_fu_4785_p1 ^ tmp_64_fu_4765_p4);

assign xor_ln1545_47_fu_5145_p2 = (tmp_75_fu_4857_p4 ^ tmp_73_fu_4843_p4);

assign xor_ln1545_49_fu_5157_p2 = (tmp_68_fu_4799_p4 ^ tmp_63_fu_4755_p4);

assign xor_ln1545_50_fu_5169_p2 = (xor_ln1545_51_fu_5163_p2 ^ xor_ln1545_49_fu_5157_p2);

assign xor_ln1545_51_fu_5163_p2 = (trunc_ln674_14_fu_4819_p1 ^ tmp_77_fu_4877_p4);

assign xor_ln1545_52_fu_6074_p2 = (tmp_82_fu_5568_p4 ^ tmp_80_fu_5554_p4);

assign xor_ln1545_53_fu_6086_p2 = (xor_ln1545_54_fu_6080_p2 ^ xor_ln1545_52_fu_6074_p2);

assign xor_ln1545_54_fu_6080_p2 = (trunc_ln674_19_fu_5632_p1 ^ tmp_87_fu_5612_p4);

assign xor_ln1545_55_fu_6092_p2 = (trunc_ln674_16_fu_5530_p1 ^ tmp_84_fu_5588_p4);

assign xor_ln1545_56_fu_6104_p2 = (xor_ln1545_57_fu_6098_p2 ^ xor_ln1545_55_fu_6092_p2);

assign xor_ln1545_57_fu_6098_p2 = (tmp_91_fu_5646_p4 ^ tmp_86_fu_5602_p4);

assign xor_ln1545_58_fu_6110_p2 = (trunc_ln674_17_fu_5564_p1 ^ tmp_79_fu_5544_p4);

assign xor_ln1545_59_fu_6122_p2 = (xor_ln1545_60_fu_6116_p2 ^ xor_ln1545_58_fu_6110_p2);

assign xor_ln1545_5_fu_4899_p2 = (xor_ln1545_fu_4887_p2 ^ xor_ln1545_6_fu_4893_p2);

assign xor_ln1545_60_fu_6116_p2 = (tmp_90_fu_5636_p4 ^ tmp_88_fu_5622_p4);

assign xor_ln1545_61_fu_6128_p2 = (tmp_83_fu_5578_p4 ^ tmp_78_fu_5534_p4);

assign xor_ln1545_62_fu_6134_p2 = (trunc_ln674_18_fu_5598_p1 ^ tmp_92_fu_5656_p4);

assign xor_ln1545_64_fu_6146_p2 = (tmp_98_fu_5704_p4 ^ tmp_96_fu_5690_p4);

assign xor_ln1545_65_fu_6158_p2 = (xor_ln1545_66_fu_6152_p2 ^ xor_ln1545_64_fu_6146_p2);

assign xor_ln1545_66_fu_6152_p2 = (trunc_ln674_23_fu_5768_p1 ^ tmp_103_fu_5748_p4);

assign xor_ln1545_67_fu_6164_p2 = (trunc_ln674_20_fu_5666_p1 ^ tmp_100_fu_5724_p4);

assign xor_ln1545_68_fu_6176_p2 = (xor_ln1545_69_fu_6170_p2 ^ xor_ln1545_67_fu_6164_p2);

assign xor_ln1545_69_fu_6170_p2 = (tmp_107_fu_5782_p4 ^ tmp_102_fu_5738_p4);

assign xor_ln1545_6_fu_4893_p2 = (trunc_ln674_3_fu_4445_p1 ^ tmp_24_fu_4425_p4);

assign xor_ln1545_70_fu_6182_p2 = (trunc_ln674_21_fu_5700_p1 ^ tmp_95_fu_5680_p4);

assign xor_ln1545_71_fu_6194_p2 = (xor_ln1545_72_fu_6188_p2 ^ xor_ln1545_70_fu_6182_p2);

assign xor_ln1545_72_fu_6188_p2 = (tmp_106_fu_5772_p4 ^ tmp_104_fu_5758_p4);

assign xor_ln1545_73_fu_6200_p2 = (tmp_99_fu_5714_p4 ^ tmp_94_fu_5670_p4);

assign xor_ln1545_74_fu_6212_p2 = (xor_ln1545_75_fu_6206_p2 ^ xor_ln1545_73_fu_6200_p2);

assign xor_ln1545_75_fu_6206_p2 = (trunc_ln674_22_fu_5734_p1 ^ tmp_108_fu_5792_p4);

assign xor_ln1545_76_fu_6218_p2 = (tmp_114_fu_5840_p4 ^ tmp_112_fu_5826_p4);

assign xor_ln1545_77_fu_6230_p2 = (xor_ln1545_78_fu_6224_p2 ^ xor_ln1545_76_fu_6218_p2);

assign xor_ln1545_78_fu_6224_p2 = (trunc_ln674_27_fu_5904_p1 ^ tmp_119_fu_5884_p4);

assign xor_ln1545_79_fu_6236_p2 = (trunc_ln674_24_fu_5802_p1 ^ tmp_116_fu_5860_p4);

assign xor_ln1545_7_fu_4905_p2 = (trunc_ln674_fu_4343_p1 ^ tmp_21_fu_4401_p4);

assign xor_ln1545_80_fu_6248_p2 = (xor_ln1545_81_fu_6242_p2 ^ xor_ln1545_79_fu_6236_p2);

assign xor_ln1545_81_fu_6242_p2 = (tmp_123_fu_5918_p4 ^ tmp_118_fu_5874_p4);

assign xor_ln1545_82_fu_6254_p2 = (trunc_ln674_25_fu_5836_p1 ^ tmp_111_fu_5816_p4);

assign xor_ln1545_83_fu_6260_p2 = (tmp_122_fu_5908_p4 ^ tmp_120_fu_5894_p4);

assign xor_ln1545_85_fu_6272_p2 = (tmp_115_fu_5850_p4 ^ tmp_110_fu_5806_p4);

assign xor_ln1545_86_fu_6284_p2 = (xor_ln1545_87_fu_6278_p2 ^ xor_ln1545_85_fu_6272_p2);

assign xor_ln1545_87_fu_6278_p2 = (trunc_ln674_26_fu_5870_p1 ^ tmp_124_fu_5928_p4);

assign xor_ln1545_88_fu_6290_p2 = (tmp_130_fu_5976_p4 ^ tmp_128_fu_5962_p4);

assign xor_ln1545_89_fu_6302_p2 = (xor_ln1545_90_fu_6296_p2 ^ xor_ln1545_88_fu_6290_p2);

assign xor_ln1545_8_fu_4917_p2 = (xor_ln1545_9_fu_4911_p2 ^ xor_ln1545_7_fu_4905_p2);

assign xor_ln1545_90_fu_6296_p2 = (trunc_ln674_31_fu_6040_p1 ^ tmp_135_fu_6020_p4);

assign xor_ln1545_91_fu_6308_p2 = (trunc_ln674_28_fu_5938_p1 ^ tmp_132_fu_5996_p4);

assign xor_ln1545_92_fu_6314_p2 = (tmp_139_fu_6054_p4 ^ tmp_134_fu_6010_p4);

assign xor_ln1545_94_fu_6326_p2 = (trunc_ln674_29_fu_5972_p1 ^ tmp_127_fu_5952_p4);

assign xor_ln1545_95_fu_6332_p2 = (tmp_138_fu_6044_p4 ^ tmp_136_fu_6030_p4);

assign xor_ln1545_97_fu_6344_p2 = (tmp_131_fu_5986_p4 ^ tmp_126_fu_5942_p4);

assign xor_ln1545_98_fu_6356_p2 = (xor_ln1545_99_fu_6350_p2 ^ xor_ln1545_97_fu_6344_p2);

assign xor_ln1545_99_fu_6350_p2 = (trunc_ln674_30_fu_6006_p1 ^ tmp_140_fu_6064_p4);

assign xor_ln1545_9_fu_4911_p2 = (tmp_28_fu_4459_p4 ^ tmp_23_fu_4415_p4);

assign xor_ln1545_fu_4887_p2 = (tmp_19_fu_4381_p4 ^ tmp_17_fu_4367_p4);

assign zext_ln708_100_fu_7554_p1 = tmp_1_V_2_fu_7507_p2;

assign zext_ln708_101_fu_7559_p1 = tmp_2_1_V_2_fu_7453_p2;

assign zext_ln708_102_fu_7564_p1 = xor_ln1545_122_fu_7399_p2;

assign zext_ln708_103_fu_7569_p1 = xor_ln1545_113_fu_7345_p2;

assign zext_ln708_104_fu_7574_p1 = xor_ln1545_104_fu_7291_p2;

assign zext_ln708_105_fu_7579_p1 = tmp_2_2_V_2_fu_7525_p2;

assign zext_ln708_106_fu_7584_p1 = xor_ln1545_134_fu_7471_p2;

assign zext_ln708_107_fu_7589_p1 = xor_ln1545_125_fu_7417_p2;

assign zext_ln708_108_fu_7594_p1 = xor_ln1545_116_fu_7363_p2;

assign zext_ln708_109_fu_7599_p1 = xor_ln1545_107_fu_7309_p2;

assign zext_ln708_10_fu_3943_p1 = tmp_7_fu_3933_p4;

assign zext_ln708_110_fu_7604_p1 = xor_ln1545_146_fu_7543_p2;

assign zext_ln708_111_fu_7609_p1 = xor_ln1545_137_fu_7489_p2;

assign zext_ln708_112_fu_7614_p1 = xor_ln1545_128_fu_7435_p2;

assign zext_ln708_113_fu_7619_p1 = xor_ln1545_119_fu_7381_p2;

assign zext_ln708_114_fu_7624_p1 = tmp_3_V_2_fu_7327_p2;

assign zext_ln708_115_fu_7674_p1 = trunc_ln708_4_fu_7670_p1;

assign zext_ln708_116_fu_7689_p1 = tmp_207_fu_7679_p4;

assign zext_ln708_117_fu_7704_p1 = tmp_211_fu_7694_p4;

assign zext_ln708_118_fu_7719_p1 = tmp_215_fu_7709_p4;

assign zext_ln708_119_fu_7734_p1 = tmp_219_fu_7724_p4;

assign zext_ln708_11_fu_3958_p1 = tmp_4_fu_3948_p4;

assign zext_ln708_120_fu_7749_p1 = tmp_223_fu_7739_p4;

assign zext_ln708_121_fu_7764_p1 = tmp_227_fu_7754_p4;

assign zext_ln708_122_fu_7779_p1 = tmp_231_fu_7769_p4;

assign zext_ln708_123_fu_7794_p1 = tmp_235_fu_7784_p4;

assign zext_ln708_124_fu_7809_p1 = tmp_239_fu_7799_p4;

assign zext_ln708_125_fu_7824_p1 = tmp_243_fu_7814_p4;

assign zext_ln708_126_fu_7839_p1 = tmp_247_fu_7829_p4;

assign zext_ln708_127_fu_7854_p1 = tmp_251_fu_7844_p4;

assign zext_ln708_128_fu_7869_p1 = tmp_255_fu_7859_p4;

assign zext_ln708_129_fu_7884_p1 = tmp_259_fu_7874_p4;

assign zext_ln708_12_fu_3973_p1 = tmp_9_fu_3963_p4;

assign zext_ln708_130_fu_7899_p1 = tmp_263_fu_7889_p4;

assign zext_ln708_131_fu_8736_p1 = xor_ln1545_149_fu_8460_p2;

assign zext_ln708_132_fu_8741_p1 = tmp_1_V_3_fu_8694_p2;

assign zext_ln708_133_fu_8746_p1 = tmp_2_1_V_3_fu_8640_p2;

assign zext_ln708_134_fu_8751_p1 = xor_ln1545_170_fu_8586_p2;

assign zext_ln708_135_fu_8756_p1 = xor_ln1545_161_fu_8532_p2;

assign zext_ln708_136_fu_8761_p1 = xor_ln1545_152_fu_8478_p2;

assign zext_ln708_137_fu_8766_p1 = tmp_2_2_V_3_fu_8712_p2;

assign zext_ln708_138_fu_8771_p1 = xor_ln1545_182_fu_8658_p2;

assign zext_ln708_139_fu_8776_p1 = xor_ln1545_173_fu_8604_p2;

assign zext_ln708_13_fu_3988_p1 = tmp_8_fu_3978_p4;

assign zext_ln708_140_fu_8781_p1 = xor_ln1545_164_fu_8550_p2;

assign zext_ln708_141_fu_8786_p1 = xor_ln1545_155_fu_8496_p2;

assign zext_ln708_142_fu_8791_p1 = xor_ln1545_194_fu_8730_p2;

assign zext_ln708_143_fu_8796_p1 = xor_ln1545_185_fu_8676_p2;

assign zext_ln708_144_fu_8801_p1 = xor_ln1545_176_fu_8622_p2;

assign zext_ln708_145_fu_8806_p1 = xor_ln1545_167_fu_8568_p2;

assign zext_ln708_146_fu_8811_p1 = tmp_3_V_3_fu_8514_p2;

assign zext_ln708_147_fu_8861_p1 = trunc_ln708_5_fu_8857_p1;

assign zext_ln708_148_fu_8876_p1 = tmp_270_fu_8866_p4;

assign zext_ln708_149_fu_8891_p1 = tmp_274_fu_8881_p4;

assign zext_ln708_14_fu_4003_p1 = tmp_10_fu_3993_p4;

assign zext_ln708_150_fu_8906_p1 = tmp_278_fu_8896_p4;

assign zext_ln708_151_fu_8921_p1 = tmp_282_fu_8911_p4;

assign zext_ln708_152_fu_8936_p1 = tmp_286_fu_8926_p4;

assign zext_ln708_153_fu_8951_p1 = tmp_290_fu_8941_p4;

assign zext_ln708_154_fu_8966_p1 = tmp_294_fu_8956_p4;

assign zext_ln708_155_fu_8981_p1 = tmp_298_fu_8971_p4;

assign zext_ln708_156_fu_8996_p1 = tmp_302_fu_8986_p4;

assign zext_ln708_157_fu_9011_p1 = tmp_306_fu_9001_p4;

assign zext_ln708_158_fu_9026_p1 = tmp_310_fu_9016_p4;

assign zext_ln708_159_fu_9041_p1 = tmp_314_fu_9031_p4;

assign zext_ln708_15_fu_4018_p1 = tmp_11_fu_4008_p4;

assign zext_ln708_160_fu_9056_p1 = tmp_318_fu_9046_p4;

assign zext_ln708_161_fu_9071_p1 = tmp_322_fu_9061_p4;

assign zext_ln708_162_fu_9086_p1 = tmp_326_fu_9076_p4;

assign zext_ln708_163_fu_9923_p1 = xor_ln1545_197_fu_9647_p2;

assign zext_ln708_164_fu_9928_p1 = tmp_1_V_4_fu_9881_p2;

assign zext_ln708_165_fu_9933_p1 = tmp_2_1_V_4_fu_9827_p2;

assign zext_ln708_166_fu_9938_p1 = xor_ln1545_218_fu_9773_p2;

assign zext_ln708_167_fu_9943_p1 = xor_ln1545_209_fu_9719_p2;

assign zext_ln708_168_fu_9948_p1 = xor_ln1545_200_fu_9665_p2;

assign zext_ln708_169_fu_9953_p1 = tmp_2_2_V_4_fu_9899_p2;

assign zext_ln708_16_fu_4033_p1 = tmp_12_fu_4023_p4;

assign zext_ln708_170_fu_9958_p1 = xor_ln1545_230_fu_9845_p2;

assign zext_ln708_171_fu_9963_p1 = xor_ln1545_221_fu_9791_p2;

assign zext_ln708_172_fu_9968_p1 = xor_ln1545_212_fu_9737_p2;

assign zext_ln708_173_fu_9973_p1 = xor_ln1545_203_fu_9683_p2;

assign zext_ln708_174_fu_9978_p1 = xor_ln1545_242_fu_9917_p2;

assign zext_ln708_175_fu_9983_p1 = xor_ln1545_233_fu_9863_p2;

assign zext_ln708_176_fu_9988_p1 = xor_ln1545_224_fu_9809_p2;

assign zext_ln708_177_fu_9993_p1 = xor_ln1545_215_fu_9755_p2;

assign zext_ln708_178_fu_9998_p1 = tmp_3_V_4_fu_9701_p2;

assign zext_ln708_179_fu_10048_p1 = trunc_ln708_6_fu_10044_p1;

assign zext_ln708_17_fu_4048_p1 = tmp_13_fu_4038_p4;

assign zext_ln708_180_fu_10063_p1 = tmp_333_fu_10053_p4;

assign zext_ln708_181_fu_10078_p1 = tmp_337_fu_10068_p4;

assign zext_ln708_182_fu_10093_p1 = tmp_341_fu_10083_p4;

assign zext_ln708_183_fu_10108_p1 = tmp_345_fu_10098_p4;

assign zext_ln708_184_fu_10123_p1 = tmp_349_fu_10113_p4;

assign zext_ln708_185_fu_10138_p1 = tmp_353_fu_10128_p4;

assign zext_ln708_186_fu_10153_p1 = tmp_357_fu_10143_p4;

assign zext_ln708_187_fu_10168_p1 = tmp_361_fu_10158_p4;

assign zext_ln708_188_fu_10183_p1 = tmp_365_fu_10173_p4;

assign zext_ln708_189_fu_10198_p1 = tmp_369_fu_10188_p4;

assign zext_ln708_18_fu_4063_p1 = tmp_14_fu_4053_p4;

assign zext_ln708_190_fu_10213_p1 = tmp_373_fu_10203_p4;

assign zext_ln708_191_fu_10228_p1 = tmp_377_fu_10218_p4;

assign zext_ln708_192_fu_10243_p1 = tmp_381_fu_10233_p4;

assign zext_ln708_193_fu_10258_p1 = tmp_385_fu_10248_p4;

assign zext_ln708_194_fu_10273_p1 = tmp_389_fu_10263_p4;

assign zext_ln708_195_fu_11110_p1 = xor_ln1545_245_fu_10834_p2;

assign zext_ln708_196_fu_11115_p1 = tmp_1_V_5_fu_11068_p2;

assign zext_ln708_197_fu_11120_p1 = tmp_2_1_V_5_fu_11014_p2;

assign zext_ln708_198_fu_11125_p1 = xor_ln1545_266_fu_10960_p2;

assign zext_ln708_199_fu_11130_p1 = xor_ln1545_257_fu_10906_p2;

assign zext_ln708_19_fu_4113_p1 = trunc_ln708_1_fu_4109_p1;

assign zext_ln708_200_fu_11135_p1 = xor_ln1545_248_fu_10852_p2;

assign zext_ln708_201_fu_11140_p1 = tmp_2_2_V_5_fu_11086_p2;

assign zext_ln708_202_fu_11145_p1 = xor_ln1545_278_fu_11032_p2;

assign zext_ln708_203_fu_11150_p1 = xor_ln1545_269_fu_10978_p2;

assign zext_ln708_204_fu_11155_p1 = xor_ln1545_260_fu_10924_p2;

assign zext_ln708_205_fu_11160_p1 = xor_ln1545_251_fu_10870_p2;

assign zext_ln708_206_fu_11165_p1 = xor_ln1545_290_fu_11104_p2;

assign zext_ln708_207_fu_11170_p1 = xor_ln1545_281_fu_11050_p2;

assign zext_ln708_208_fu_11175_p1 = xor_ln1545_272_fu_10996_p2;

assign zext_ln708_209_fu_11180_p1 = xor_ln1545_263_fu_10942_p2;

assign zext_ln708_20_fu_4128_p1 = tmp_18_fu_4118_p4;

assign zext_ln708_210_fu_11185_p1 = tmp_3_V_5_fu_10888_p2;

assign zext_ln708_211_fu_11235_p1 = trunc_ln708_7_fu_11231_p1;

assign zext_ln708_212_fu_11250_p1 = tmp_396_fu_11240_p4;

assign zext_ln708_213_fu_11265_p1 = tmp_400_fu_11255_p4;

assign zext_ln708_214_fu_11280_p1 = tmp_404_fu_11270_p4;

assign zext_ln708_215_fu_11295_p1 = tmp_408_fu_11285_p4;

assign zext_ln708_216_fu_11310_p1 = tmp_412_fu_11300_p4;

assign zext_ln708_217_fu_11325_p1 = tmp_416_fu_11315_p4;

assign zext_ln708_218_fu_11340_p1 = tmp_420_fu_11330_p4;

assign zext_ln708_219_fu_11355_p1 = tmp_424_fu_11345_p4;

assign zext_ln708_21_fu_4143_p1 = tmp_22_fu_4133_p4;

assign zext_ln708_220_fu_11370_p1 = tmp_428_fu_11360_p4;

assign zext_ln708_221_fu_11385_p1 = tmp_432_fu_11375_p4;

assign zext_ln708_222_fu_11400_p1 = tmp_436_fu_11390_p4;

assign zext_ln708_223_fu_11415_p1 = tmp_440_fu_11405_p4;

assign zext_ln708_224_fu_11430_p1 = tmp_444_fu_11420_p4;

assign zext_ln708_225_fu_11445_p1 = tmp_448_fu_11435_p4;

assign zext_ln708_226_fu_11460_p1 = tmp_452_fu_11450_p4;

assign zext_ln708_227_fu_12297_p1 = xor_ln1545_293_fu_12021_p2;

assign zext_ln708_228_fu_12302_p1 = tmp_1_V_6_fu_12255_p2;

assign zext_ln708_229_fu_12307_p1 = tmp_2_1_V_6_fu_12201_p2;

assign zext_ln708_22_fu_4158_p1 = tmp_26_fu_4148_p4;

assign zext_ln708_230_fu_12312_p1 = xor_ln1545_314_fu_12147_p2;

assign zext_ln708_231_fu_12317_p1 = xor_ln1545_305_fu_12093_p2;

assign zext_ln708_232_fu_12322_p1 = xor_ln1545_296_fu_12039_p2;

assign zext_ln708_233_fu_12327_p1 = tmp_2_2_V_6_fu_12273_p2;

assign zext_ln708_234_fu_12332_p1 = xor_ln1545_326_fu_12219_p2;

assign zext_ln708_235_fu_12337_p1 = xor_ln1545_317_fu_12165_p2;

assign zext_ln708_236_fu_12342_p1 = xor_ln1545_308_fu_12111_p2;

assign zext_ln708_237_fu_12347_p1 = xor_ln1545_299_fu_12057_p2;

assign zext_ln708_238_fu_12352_p1 = xor_ln1545_338_fu_12291_p2;

assign zext_ln708_239_fu_12357_p1 = xor_ln1545_329_fu_12237_p2;

assign zext_ln708_23_fu_4173_p1 = tmp_30_fu_4163_p4;

assign zext_ln708_240_fu_12362_p1 = xor_ln1545_320_fu_12183_p2;

assign zext_ln708_241_fu_12367_p1 = xor_ln1545_311_fu_12129_p2;

assign zext_ln708_242_fu_12372_p1 = tmp_3_V_6_fu_12075_p2;

assign zext_ln708_243_fu_12422_p1 = trunc_ln708_8_fu_12418_p1;

assign zext_ln708_244_fu_12437_p1 = tmp_459_fu_12427_p4;

assign zext_ln708_245_fu_12452_p1 = tmp_463_fu_12442_p4;

assign zext_ln708_246_fu_12467_p1 = tmp_467_fu_12457_p4;

assign zext_ln708_247_fu_12482_p1 = tmp_471_fu_12472_p4;

assign zext_ln708_248_fu_12497_p1 = tmp_475_fu_12487_p4;

assign zext_ln708_249_fu_12512_p1 = tmp_479_fu_12502_p4;

assign zext_ln708_24_fu_4188_p1 = tmp_34_fu_4178_p4;

assign zext_ln708_250_fu_12527_p1 = tmp_483_fu_12517_p4;

assign zext_ln708_251_fu_12542_p1 = tmp_487_fu_12532_p4;

assign zext_ln708_252_fu_12557_p1 = tmp_491_fu_12547_p4;

assign zext_ln708_253_fu_12572_p1 = tmp_495_fu_12562_p4;

assign zext_ln708_254_fu_12587_p1 = tmp_499_fu_12577_p4;

assign zext_ln708_255_fu_12602_p1 = tmp_503_fu_12592_p4;

assign zext_ln708_256_fu_12617_p1 = tmp_507_fu_12607_p4;

assign zext_ln708_257_fu_12632_p1 = tmp_511_fu_12622_p4;

assign zext_ln708_258_fu_12647_p1 = tmp_515_fu_12637_p4;

assign zext_ln708_259_fu_13484_p1 = xor_ln1545_341_fu_13208_p2;

assign zext_ln708_25_fu_4203_p1 = tmp_38_fu_4193_p4;

assign zext_ln708_260_fu_13489_p1 = tmp_1_V_7_fu_13442_p2;

assign zext_ln708_261_fu_13494_p1 = tmp_2_1_V_7_fu_13388_p2;

assign zext_ln708_262_fu_13499_p1 = xor_ln1545_362_fu_13334_p2;

assign zext_ln708_263_fu_13504_p1 = xor_ln1545_353_fu_13280_p2;

assign zext_ln708_264_fu_13509_p1 = xor_ln1545_344_fu_13226_p2;

assign zext_ln708_265_fu_13514_p1 = tmp_2_2_V_7_fu_13460_p2;

assign zext_ln708_266_fu_13519_p1 = xor_ln1545_374_fu_13406_p2;

assign zext_ln708_267_fu_13524_p1 = xor_ln1545_365_fu_13352_p2;

assign zext_ln708_268_fu_13529_p1 = xor_ln1545_356_fu_13298_p2;

assign zext_ln708_269_fu_13534_p1 = xor_ln1545_347_fu_13244_p2;

assign zext_ln708_26_fu_4218_p1 = tmp_42_fu_4208_p4;

assign zext_ln708_270_fu_13539_p1 = xor_ln1545_386_fu_13478_p2;

assign zext_ln708_271_fu_13544_p1 = xor_ln1545_377_fu_13424_p2;

assign zext_ln708_272_fu_13549_p1 = xor_ln1545_368_fu_13370_p2;

assign zext_ln708_273_fu_13554_p1 = xor_ln1545_359_fu_13316_p2;

assign zext_ln708_274_fu_13559_p1 = tmp_3_V_7_fu_13262_p2;

assign zext_ln708_275_fu_13609_p1 = trunc_ln708_9_fu_13605_p1;

assign zext_ln708_276_fu_13624_p1 = tmp_522_fu_13614_p4;

assign zext_ln708_277_fu_13639_p1 = tmp_526_fu_13629_p4;

assign zext_ln708_278_fu_13654_p1 = tmp_530_fu_13644_p4;

assign zext_ln708_279_fu_13669_p1 = tmp_534_fu_13659_p4;

assign zext_ln708_27_fu_4233_p1 = tmp_46_fu_4223_p4;

assign zext_ln708_280_fu_13684_p1 = tmp_538_fu_13674_p4;

assign zext_ln708_281_fu_13699_p1 = tmp_542_fu_13689_p4;

assign zext_ln708_282_fu_13714_p1 = tmp_546_fu_13704_p4;

assign zext_ln708_283_fu_13729_p1 = tmp_550_fu_13719_p4;

assign zext_ln708_284_fu_13744_p1 = tmp_554_fu_13734_p4;

assign zext_ln708_285_fu_13759_p1 = tmp_558_fu_13749_p4;

assign zext_ln708_286_fu_13774_p1 = tmp_562_fu_13764_p4;

assign zext_ln708_287_fu_13789_p1 = tmp_566_fu_13779_p4;

assign zext_ln708_288_fu_13804_p1 = tmp_570_fu_13794_p4;

assign zext_ln708_289_fu_13819_p1 = tmp_574_fu_13809_p4;

assign zext_ln708_28_fu_4248_p1 = tmp_50_fu_4238_p4;

assign zext_ln708_290_fu_13834_p1 = tmp_578_fu_13824_p4;

assign zext_ln708_291_fu_14671_p1 = xor_ln1545_389_fu_14395_p2;

assign zext_ln708_292_fu_14676_p1 = tmp_1_V_8_fu_14629_p2;

assign zext_ln708_293_fu_14681_p1 = tmp_2_1_V_8_fu_14575_p2;

assign zext_ln708_294_fu_14686_p1 = xor_ln1545_410_fu_14521_p2;

assign zext_ln708_295_fu_14691_p1 = xor_ln1545_401_fu_14467_p2;

assign zext_ln708_296_fu_14696_p1 = xor_ln1545_392_fu_14413_p2;

assign zext_ln708_297_fu_14701_p1 = tmp_2_2_V_8_fu_14647_p2;

assign zext_ln708_298_fu_14706_p1 = xor_ln1545_422_fu_14593_p2;

assign zext_ln708_299_fu_14711_p1 = xor_ln1545_413_fu_14539_p2;

assign zext_ln708_29_fu_4263_p1 = tmp_54_fu_4253_p4;

assign zext_ln708_300_fu_14716_p1 = xor_ln1545_404_fu_14485_p2;

assign zext_ln708_301_fu_14721_p1 = xor_ln1545_395_fu_14431_p2;

assign zext_ln708_302_fu_14726_p1 = xor_ln1545_434_fu_14665_p2;

assign zext_ln708_303_fu_14731_p1 = xor_ln1545_425_fu_14611_p2;

assign zext_ln708_304_fu_14736_p1 = xor_ln1545_416_fu_14557_p2;

assign zext_ln708_305_fu_14741_p1 = xor_ln1545_407_fu_14503_p2;

assign zext_ln708_306_fu_14746_p1 = tmp_3_V_8_fu_14449_p2;

assign zext_ln708_30_fu_4278_p1 = tmp_58_fu_4268_p4;

assign zext_ln708_31_fu_4293_p1 = tmp_62_fu_4283_p4;

assign zext_ln708_32_fu_4308_p1 = tmp_66_fu_4298_p4;

assign zext_ln708_33_fu_4323_p1 = tmp_70_fu_4313_p4;

assign zext_ln708_34_fu_4338_p1 = tmp_74_fu_4328_p4;

assign zext_ln708_35_fu_5175_p1 = xor_ln1545_5_fu_4899_p2;

assign zext_ln708_36_fu_5180_p1 = tmp_1_V_fu_5133_p2;

assign zext_ln708_37_fu_5185_p1 = tmp_2_1_V_fu_5079_p2;

assign zext_ln708_38_fu_5190_p1 = xor_ln1545_26_fu_5025_p2;

assign zext_ln708_39_fu_5195_p1 = xor_ln1545_17_fu_4971_p2;

assign zext_ln708_40_fu_5200_p1 = xor_ln1545_8_fu_4917_p2;

assign zext_ln708_41_fu_5205_p1 = tmp_2_2_V_fu_5151_p2;

assign zext_ln708_42_fu_5210_p1 = xor_ln1545_38_fu_5097_p2;

assign zext_ln708_43_fu_5215_p1 = xor_ln1545_29_fu_5043_p2;

assign zext_ln708_44_fu_5220_p1 = xor_ln1545_20_fu_4989_p2;

assign zext_ln708_45_fu_5225_p1 = xor_ln1545_11_fu_4935_p2;

assign zext_ln708_46_fu_5230_p1 = xor_ln1545_50_fu_5169_p2;

assign zext_ln708_47_fu_5235_p1 = xor_ln1545_41_fu_5115_p2;

assign zext_ln708_48_fu_5240_p1 = xor_ln1545_32_fu_5061_p2;

assign zext_ln708_49_fu_5245_p1 = xor_ln1545_23_fu_5007_p2;

assign zext_ln708_4_fu_3853_p1 = tmp_1_fu_3843_p4;

assign zext_ln708_50_fu_5250_p1 = tmp_3_V_fu_4953_p2;

assign zext_ln708_51_fu_5300_p1 = trunc_ln708_2_fu_5296_p1;

assign zext_ln708_52_fu_5315_p1 = tmp_81_fu_5305_p4;

assign zext_ln708_53_fu_5330_p1 = tmp_85_fu_5320_p4;

assign zext_ln708_54_fu_5345_p1 = tmp_89_fu_5335_p4;

assign zext_ln708_55_fu_5360_p1 = tmp_93_fu_5350_p4;

assign zext_ln708_56_fu_5375_p1 = tmp_97_fu_5365_p4;

assign zext_ln708_57_fu_5390_p1 = tmp_101_fu_5380_p4;

assign zext_ln708_58_fu_5405_p1 = tmp_105_fu_5395_p4;

assign zext_ln708_59_fu_5420_p1 = tmp_109_fu_5410_p4;

assign zext_ln708_5_fu_3868_p1 = tmp_2_fu_3858_p4;

assign zext_ln708_60_fu_5435_p1 = tmp_113_fu_5425_p4;

assign zext_ln708_61_fu_5450_p1 = tmp_117_fu_5440_p4;

assign zext_ln708_62_fu_5465_p1 = tmp_121_fu_5455_p4;

assign zext_ln708_63_fu_5480_p1 = tmp_125_fu_5470_p4;

assign zext_ln708_64_fu_5495_p1 = tmp_129_fu_5485_p4;

assign zext_ln708_65_fu_5510_p1 = tmp_133_fu_5500_p4;

assign zext_ln708_66_fu_5525_p1 = tmp_137_fu_5515_p4;

assign zext_ln708_67_fu_6362_p1 = xor_ln1545_53_fu_6086_p2;

assign zext_ln708_68_fu_6367_p1 = tmp_1_V_1_fu_6320_p2;

assign zext_ln708_69_fu_6372_p1 = tmp_2_1_V_1_fu_6266_p2;

assign zext_ln708_6_fu_3883_p1 = tmp_3_fu_3873_p4;

assign zext_ln708_70_fu_6377_p1 = xor_ln1545_74_fu_6212_p2;

assign zext_ln708_71_fu_6382_p1 = xor_ln1545_65_fu_6158_p2;

assign zext_ln708_72_fu_6387_p1 = xor_ln1545_56_fu_6104_p2;

assign zext_ln708_73_fu_6392_p1 = tmp_2_2_V_1_fu_6338_p2;

assign zext_ln708_74_fu_6397_p1 = xor_ln1545_86_fu_6284_p2;

assign zext_ln708_75_fu_6402_p1 = xor_ln1545_77_fu_6230_p2;

assign zext_ln708_76_fu_6407_p1 = xor_ln1545_68_fu_6176_p2;

assign zext_ln708_77_fu_6412_p1 = xor_ln1545_59_fu_6122_p2;

assign zext_ln708_78_fu_6417_p1 = xor_ln1545_98_fu_6356_p2;

assign zext_ln708_79_fu_6422_p1 = xor_ln1545_89_fu_6302_p2;

assign zext_ln708_7_fu_3898_p1 = tmp_s_fu_3888_p4;

assign zext_ln708_80_fu_6427_p1 = xor_ln1545_80_fu_6248_p2;

assign zext_ln708_81_fu_6432_p1 = xor_ln1545_71_fu_6194_p2;

assign zext_ln708_82_fu_6437_p1 = tmp_3_V_1_fu_6140_p2;

assign zext_ln708_83_fu_6487_p1 = trunc_ln708_3_fu_6483_p1;

assign zext_ln708_84_fu_6502_p1 = tmp_144_fu_6492_p4;

assign zext_ln708_85_fu_6517_p1 = tmp_148_fu_6507_p4;

assign zext_ln708_86_fu_6532_p1 = tmp_152_fu_6522_p4;

assign zext_ln708_87_fu_6547_p1 = tmp_156_fu_6537_p4;

assign zext_ln708_88_fu_6562_p1 = tmp_160_fu_6552_p4;

assign zext_ln708_89_fu_6577_p1 = tmp_164_fu_6567_p4;

assign zext_ln708_8_fu_3913_p1 = tmp_5_fu_3903_p4;

assign zext_ln708_90_fu_6592_p1 = tmp_168_fu_6582_p4;

assign zext_ln708_91_fu_6607_p1 = tmp_172_fu_6597_p4;

assign zext_ln708_92_fu_6622_p1 = tmp_176_fu_6612_p4;

assign zext_ln708_93_fu_6637_p1 = tmp_180_fu_6627_p4;

assign zext_ln708_94_fu_6652_p1 = tmp_184_fu_6642_p4;

assign zext_ln708_95_fu_6667_p1 = tmp_188_fu_6657_p4;

assign zext_ln708_96_fu_6682_p1 = tmp_192_fu_6672_p4;

assign zext_ln708_97_fu_6697_p1 = tmp_196_fu_6687_p4;

assign zext_ln708_98_fu_6712_p1 = tmp_200_fu_6702_p4;

assign zext_ln708_99_fu_7549_p1 = xor_ln1545_101_fu_7273_p2;

assign zext_ln708_9_fu_3928_p1 = tmp_6_fu_3918_p4;

assign zext_ln708_fu_3838_p1 = trunc_ln708_fu_3834_p1;

endmodule //testDec_process_r
