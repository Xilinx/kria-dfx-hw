
    wire reset;
    wire clock;
    assign reset = ap_rst_n;
    assign clock = ap_clk;
    wire [5:0] proc_0_data_FIFO_blk;
    wire [5:0] proc_0_data_PIPO_blk;
    wire [5:0] proc_0_start_FIFO_blk;
    wire [5:0] proc_0_TLF_FIFO_blk;
    wire [5:0] proc_0_input_sync_blk;
    wire [5:0] proc_0_output_sync_blk;
    wire [5:0] proc_dep_vld_vec_0;
    reg [5:0] proc_dep_vld_vec_0_reg;
    wire [5:0] in_chan_dep_vld_vec_0;
    wire [197:0] in_chan_dep_data_vec_0;
    wire [5:0] token_in_vec_0;
    wire [5:0] out_chan_dep_vld_vec_0;
    wire [32:0] out_chan_dep_data_0;
    wire [5:0] token_out_vec_0;
    wire dl_detect_out_0;
    wire dep_chan_vld_1_0;
    wire [32:0] dep_chan_data_1_0;
    wire token_1_0;
    wire dep_chan_vld_2_0;
    wire [32:0] dep_chan_data_2_0;
    wire token_2_0;
    wire dep_chan_vld_11_0;
    wire [32:0] dep_chan_data_11_0;
    wire token_11_0;
    wire dep_chan_vld_12_0;
    wire [32:0] dep_chan_data_12_0;
    wire token_12_0;
    wire dep_chan_vld_23_0;
    wire [32:0] dep_chan_data_23_0;
    wire token_23_0;
    wire dep_chan_vld_24_0;
    wire [32:0] dep_chan_data_24_0;
    wire token_24_0;
    wire [3:0] proc_1_data_FIFO_blk;
    wire [3:0] proc_1_data_PIPO_blk;
    wire [3:0] proc_1_start_FIFO_blk;
    wire [3:0] proc_1_TLF_FIFO_blk;
    wire [3:0] proc_1_input_sync_blk;
    wire [3:0] proc_1_output_sync_blk;
    wire [3:0] proc_dep_vld_vec_1;
    reg [3:0] proc_dep_vld_vec_1_reg;
    wire [4:0] in_chan_dep_vld_vec_1;
    wire [164:0] in_chan_dep_data_vec_1;
    wire [4:0] token_in_vec_1;
    wire [3:0] out_chan_dep_vld_vec_1;
    wire [32:0] out_chan_dep_data_1;
    wire [3:0] token_out_vec_1;
    wire dl_detect_out_1;
    wire dep_chan_vld_0_1;
    wire [32:0] dep_chan_data_0_1;
    wire token_0_1;
    wire dep_chan_vld_2_1;
    wire [32:0] dep_chan_data_2_1;
    wire token_2_1;
    wire dep_chan_vld_12_1;
    wire [32:0] dep_chan_data_12_1;
    wire token_12_1;
    wire dep_chan_vld_22_1;
    wire [32:0] dep_chan_data_22_1;
    wire token_22_1;
    wire dep_chan_vld_24_1;
    wire [32:0] dep_chan_data_24_1;
    wire token_24_1;
    wire [4:0] proc_2_data_FIFO_blk;
    wire [4:0] proc_2_data_PIPO_blk;
    wire [4:0] proc_2_start_FIFO_blk;
    wire [4:0] proc_2_TLF_FIFO_blk;
    wire [4:0] proc_2_input_sync_blk;
    wire [4:0] proc_2_output_sync_blk;
    wire [4:0] proc_dep_vld_vec_2;
    reg [4:0] proc_dep_vld_vec_2_reg;
    wire [4:0] in_chan_dep_vld_vec_2;
    wire [164:0] in_chan_dep_data_vec_2;
    wire [4:0] token_in_vec_2;
    wire [4:0] out_chan_dep_vld_vec_2;
    wire [32:0] out_chan_dep_data_2;
    wire [4:0] token_out_vec_2;
    wire dl_detect_out_2;
    wire dep_chan_vld_0_2;
    wire [32:0] dep_chan_data_0_2;
    wire token_0_2;
    wire dep_chan_vld_1_2;
    wire [32:0] dep_chan_data_1_2;
    wire token_1_2;
    wire dep_chan_vld_12_2;
    wire [32:0] dep_chan_data_12_2;
    wire token_12_2;
    wire dep_chan_vld_21_2;
    wire [32:0] dep_chan_data_21_2;
    wire token_21_2;
    wire dep_chan_vld_23_2;
    wire [32:0] dep_chan_data_23_2;
    wire token_23_2;
    wire [2:0] proc_3_data_FIFO_blk;
    wire [2:0] proc_3_data_PIPO_blk;
    wire [2:0] proc_3_start_FIFO_blk;
    wire [2:0] proc_3_TLF_FIFO_blk;
    wire [2:0] proc_3_input_sync_blk;
    wire [2:0] proc_3_output_sync_blk;
    wire [2:0] proc_dep_vld_vec_3;
    reg [2:0] proc_dep_vld_vec_3_reg;
    wire [2:0] in_chan_dep_vld_vec_3;
    wire [98:0] in_chan_dep_data_vec_3;
    wire [2:0] token_in_vec_3;
    wire [2:0] out_chan_dep_vld_vec_3;
    wire [32:0] out_chan_dep_data_3;
    wire [2:0] token_out_vec_3;
    wire dl_detect_out_3;
    wire dep_chan_vld_4_3;
    wire [32:0] dep_chan_data_4_3;
    wire token_4_3;
    wire dep_chan_vld_5_3;
    wire [32:0] dep_chan_data_5_3;
    wire token_5_3;
    wire dep_chan_vld_9_3;
    wire [32:0] dep_chan_data_9_3;
    wire token_9_3;
    wire [2:0] proc_4_data_FIFO_blk;
    wire [2:0] proc_4_data_PIPO_blk;
    wire [2:0] proc_4_start_FIFO_blk;
    wire [2:0] proc_4_TLF_FIFO_blk;
    wire [2:0] proc_4_input_sync_blk;
    wire [2:0] proc_4_output_sync_blk;
    wire [2:0] proc_dep_vld_vec_4;
    reg [2:0] proc_dep_vld_vec_4_reg;
    wire [2:0] in_chan_dep_vld_vec_4;
    wire [98:0] in_chan_dep_data_vec_4;
    wire [2:0] token_in_vec_4;
    wire [2:0] out_chan_dep_vld_vec_4;
    wire [32:0] out_chan_dep_data_4;
    wire [2:0] token_out_vec_4;
    wire dl_detect_out_4;
    wire dep_chan_vld_3_4;
    wire [32:0] dep_chan_data_3_4;
    wire token_3_4;
    wire dep_chan_vld_6_4;
    wire [32:0] dep_chan_data_6_4;
    wire token_6_4;
    wire dep_chan_vld_9_4;
    wire [32:0] dep_chan_data_9_4;
    wire token_9_4;
    wire [2:0] proc_5_data_FIFO_blk;
    wire [2:0] proc_5_data_PIPO_blk;
    wire [2:0] proc_5_start_FIFO_blk;
    wire [2:0] proc_5_TLF_FIFO_blk;
    wire [2:0] proc_5_input_sync_blk;
    wire [2:0] proc_5_output_sync_blk;
    wire [2:0] proc_dep_vld_vec_5;
    reg [2:0] proc_dep_vld_vec_5_reg;
    wire [2:0] in_chan_dep_vld_vec_5;
    wire [98:0] in_chan_dep_data_vec_5;
    wire [2:0] token_in_vec_5;
    wire [2:0] out_chan_dep_vld_vec_5;
    wire [32:0] out_chan_dep_data_5;
    wire [2:0] token_out_vec_5;
    wire dl_detect_out_5;
    wire dep_chan_vld_3_5;
    wire [32:0] dep_chan_data_3_5;
    wire token_3_5;
    wire dep_chan_vld_9_5;
    wire [32:0] dep_chan_data_9_5;
    wire token_9_5;
    wire dep_chan_vld_10_5;
    wire [32:0] dep_chan_data_10_5;
    wire token_10_5;
    wire [1:0] proc_6_data_FIFO_blk;
    wire [1:0] proc_6_data_PIPO_blk;
    wire [1:0] proc_6_start_FIFO_blk;
    wire [1:0] proc_6_TLF_FIFO_blk;
    wire [1:0] proc_6_input_sync_blk;
    wire [1:0] proc_6_output_sync_blk;
    wire [1:0] proc_dep_vld_vec_6;
    reg [1:0] proc_dep_vld_vec_6_reg;
    wire [2:0] in_chan_dep_vld_vec_6;
    wire [98:0] in_chan_dep_data_vec_6;
    wire [2:0] token_in_vec_6;
    wire [1:0] out_chan_dep_vld_vec_6;
    wire [32:0] out_chan_dep_data_6;
    wire [1:0] token_out_vec_6;
    wire dl_detect_out_6;
    wire dep_chan_vld_4_6;
    wire [32:0] dep_chan_data_4_6;
    wire token_4_6;
    wire dep_chan_vld_7_6;
    wire [32:0] dep_chan_data_7_6;
    wire token_7_6;
    wire dep_chan_vld_10_6;
    wire [32:0] dep_chan_data_10_6;
    wire token_10_6;
    wire [0:0] proc_7_data_FIFO_blk;
    wire [0:0] proc_7_data_PIPO_blk;
    wire [0:0] proc_7_start_FIFO_blk;
    wire [0:0] proc_7_TLF_FIFO_blk;
    wire [0:0] proc_7_input_sync_blk;
    wire [0:0] proc_7_output_sync_blk;
    wire [0:0] proc_dep_vld_vec_7;
    reg [0:0] proc_dep_vld_vec_7_reg;
    wire [0:0] in_chan_dep_vld_vec_7;
    wire [32:0] in_chan_dep_data_vec_7;
    wire [0:0] token_in_vec_7;
    wire [0:0] out_chan_dep_vld_vec_7;
    wire [32:0] out_chan_dep_data_7;
    wire [0:0] token_out_vec_7;
    wire dl_detect_out_7;
    wire dep_chan_vld_8_7;
    wire [32:0] dep_chan_data_8_7;
    wire token_8_7;
    wire [0:0] proc_8_data_FIFO_blk;
    wire [0:0] proc_8_data_PIPO_blk;
    wire [0:0] proc_8_start_FIFO_blk;
    wire [0:0] proc_8_TLF_FIFO_blk;
    wire [0:0] proc_8_input_sync_blk;
    wire [0:0] proc_8_output_sync_blk;
    wire [0:0] proc_dep_vld_vec_8;
    reg [0:0] proc_dep_vld_vec_8_reg;
    wire [0:0] in_chan_dep_vld_vec_8;
    wire [32:0] in_chan_dep_data_vec_8;
    wire [0:0] token_in_vec_8;
    wire [0:0] out_chan_dep_vld_vec_8;
    wire [32:0] out_chan_dep_data_8;
    wire [0:0] token_out_vec_8;
    wire dl_detect_out_8;
    wire dep_chan_vld_9_8;
    wire [32:0] dep_chan_data_9_8;
    wire token_9_8;
    wire [4:0] proc_9_data_FIFO_blk;
    wire [4:0] proc_9_data_PIPO_blk;
    wire [4:0] proc_9_start_FIFO_blk;
    wire [4:0] proc_9_TLF_FIFO_blk;
    wire [4:0] proc_9_input_sync_blk;
    wire [4:0] proc_9_output_sync_blk;
    wire [4:0] proc_dep_vld_vec_9;
    reg [4:0] proc_dep_vld_vec_9_reg;
    wire [3:0] in_chan_dep_vld_vec_9;
    wire [131:0] in_chan_dep_data_vec_9;
    wire [3:0] token_in_vec_9;
    wire [4:0] out_chan_dep_vld_vec_9;
    wire [32:0] out_chan_dep_data_9;
    wire [4:0] token_out_vec_9;
    wire dl_detect_out_9;
    wire dep_chan_vld_3_9;
    wire [32:0] dep_chan_data_3_9;
    wire token_3_9;
    wire dep_chan_vld_4_9;
    wire [32:0] dep_chan_data_4_9;
    wire token_4_9;
    wire dep_chan_vld_5_9;
    wire [32:0] dep_chan_data_5_9;
    wire token_5_9;
    wire dep_chan_vld_10_9;
    wire [32:0] dep_chan_data_10_9;
    wire token_10_9;
    wire [2:0] proc_10_data_FIFO_blk;
    wire [2:0] proc_10_data_PIPO_blk;
    wire [2:0] proc_10_start_FIFO_blk;
    wire [2:0] proc_10_TLF_FIFO_blk;
    wire [2:0] proc_10_input_sync_blk;
    wire [2:0] proc_10_output_sync_blk;
    wire [2:0] proc_dep_vld_vec_10;
    reg [2:0] proc_dep_vld_vec_10_reg;
    wire [2:0] in_chan_dep_vld_vec_10;
    wire [98:0] in_chan_dep_data_vec_10;
    wire [2:0] token_in_vec_10;
    wire [2:0] out_chan_dep_vld_vec_10;
    wire [32:0] out_chan_dep_data_10;
    wire [2:0] token_out_vec_10;
    wire dl_detect_out_10;
    wire dep_chan_vld_5_10;
    wire [32:0] dep_chan_data_5_10;
    wire token_5_10;
    wire dep_chan_vld_6_10;
    wire [32:0] dep_chan_data_6_10;
    wire token_6_10;
    wire dep_chan_vld_9_10;
    wire [32:0] dep_chan_data_9_10;
    wire token_9_10;
    wire [0:0] proc_11_data_FIFO_blk;
    wire [0:0] proc_11_data_PIPO_blk;
    wire [0:0] proc_11_start_FIFO_blk;
    wire [0:0] proc_11_TLF_FIFO_blk;
    wire [0:0] proc_11_input_sync_blk;
    wire [0:0] proc_11_output_sync_blk;
    wire [0:0] proc_dep_vld_vec_11;
    reg [0:0] proc_dep_vld_vec_11_reg;
    wire [1:0] in_chan_dep_vld_vec_11;
    wire [65:0] in_chan_dep_data_vec_11;
    wire [1:0] token_in_vec_11;
    wire [0:0] out_chan_dep_vld_vec_11;
    wire [32:0] out_chan_dep_data_11;
    wire [0:0] token_out_vec_11;
    wire dl_detect_out_11;
    wire dep_chan_vld_0_11;
    wire [32:0] dep_chan_data_0_11;
    wire token_0_11;
    wire dep_chan_vld_12_11;
    wire [32:0] dep_chan_data_12_11;
    wire token_12_11;
    wire [5:0] proc_12_data_FIFO_blk;
    wire [5:0] proc_12_data_PIPO_blk;
    wire [5:0] proc_12_start_FIFO_blk;
    wire [5:0] proc_12_TLF_FIFO_blk;
    wire [5:0] proc_12_input_sync_blk;
    wire [5:0] proc_12_output_sync_blk;
    wire [5:0] proc_dep_vld_vec_12;
    reg [5:0] proc_dep_vld_vec_12_reg;
    wire [3:0] in_chan_dep_vld_vec_12;
    wire [131:0] in_chan_dep_data_vec_12;
    wire [3:0] token_in_vec_12;
    wire [5:0] out_chan_dep_vld_vec_12;
    wire [32:0] out_chan_dep_data_12;
    wire [5:0] token_out_vec_12;
    wire dl_detect_out_12;
    wire dep_chan_vld_0_12;
    wire [32:0] dep_chan_data_0_12;
    wire token_0_12;
    wire dep_chan_vld_2_12;
    wire [32:0] dep_chan_data_2_12;
    wire token_2_12;
    wire dep_chan_vld_21_12;
    wire [32:0] dep_chan_data_21_12;
    wire token_21_12;
    wire dep_chan_vld_23_12;
    wire [32:0] dep_chan_data_23_12;
    wire token_23_12;
    wire [2:0] proc_13_data_FIFO_blk;
    wire [2:0] proc_13_data_PIPO_blk;
    wire [2:0] proc_13_start_FIFO_blk;
    wire [2:0] proc_13_TLF_FIFO_blk;
    wire [2:0] proc_13_input_sync_blk;
    wire [2:0] proc_13_output_sync_blk;
    wire [2:0] proc_dep_vld_vec_13;
    reg [2:0] proc_dep_vld_vec_13_reg;
    wire [2:0] in_chan_dep_vld_vec_13;
    wire [98:0] in_chan_dep_data_vec_13;
    wire [2:0] token_in_vec_13;
    wire [2:0] out_chan_dep_vld_vec_13;
    wire [32:0] out_chan_dep_data_13;
    wire [2:0] token_out_vec_13;
    wire dl_detect_out_13;
    wire dep_chan_vld_14_13;
    wire [32:0] dep_chan_data_14_13;
    wire token_14_13;
    wire dep_chan_vld_15_13;
    wire [32:0] dep_chan_data_15_13;
    wire token_15_13;
    wire dep_chan_vld_19_13;
    wire [32:0] dep_chan_data_19_13;
    wire token_19_13;
    wire [3:0] proc_14_data_FIFO_blk;
    wire [3:0] proc_14_data_PIPO_blk;
    wire [3:0] proc_14_start_FIFO_blk;
    wire [3:0] proc_14_TLF_FIFO_blk;
    wire [3:0] proc_14_input_sync_blk;
    wire [3:0] proc_14_output_sync_blk;
    wire [3:0] proc_dep_vld_vec_14;
    reg [3:0] proc_dep_vld_vec_14_reg;
    wire [3:0] in_chan_dep_vld_vec_14;
    wire [131:0] in_chan_dep_data_vec_14;
    wire [3:0] token_in_vec_14;
    wire [3:0] out_chan_dep_vld_vec_14;
    wire [32:0] out_chan_dep_data_14;
    wire [3:0] token_out_vec_14;
    wire dl_detect_out_14;
    wire dep_chan_vld_13_14;
    wire [32:0] dep_chan_data_13_14;
    wire token_13_14;
    wire dep_chan_vld_16_14;
    wire [32:0] dep_chan_data_16_14;
    wire token_16_14;
    wire dep_chan_vld_17_14;
    wire [32:0] dep_chan_data_17_14;
    wire token_17_14;
    wire dep_chan_vld_19_14;
    wire [32:0] dep_chan_data_19_14;
    wire token_19_14;
    wire [2:0] proc_15_data_FIFO_blk;
    wire [2:0] proc_15_data_PIPO_blk;
    wire [2:0] proc_15_start_FIFO_blk;
    wire [2:0] proc_15_TLF_FIFO_blk;
    wire [2:0] proc_15_input_sync_blk;
    wire [2:0] proc_15_output_sync_blk;
    wire [2:0] proc_dep_vld_vec_15;
    reg [2:0] proc_dep_vld_vec_15_reg;
    wire [2:0] in_chan_dep_vld_vec_15;
    wire [98:0] in_chan_dep_data_vec_15;
    wire [2:0] token_in_vec_15;
    wire [2:0] out_chan_dep_vld_vec_15;
    wire [32:0] out_chan_dep_data_15;
    wire [2:0] token_out_vec_15;
    wire dl_detect_out_15;
    wire dep_chan_vld_13_15;
    wire [32:0] dep_chan_data_13_15;
    wire token_13_15;
    wire dep_chan_vld_19_15;
    wire [32:0] dep_chan_data_19_15;
    wire token_19_15;
    wire dep_chan_vld_20_15;
    wire [32:0] dep_chan_data_20_15;
    wire token_20_15;
    wire [1:0] proc_16_data_FIFO_blk;
    wire [1:0] proc_16_data_PIPO_blk;
    wire [1:0] proc_16_start_FIFO_blk;
    wire [1:0] proc_16_TLF_FIFO_blk;
    wire [1:0] proc_16_input_sync_blk;
    wire [1:0] proc_16_output_sync_blk;
    wire [1:0] proc_dep_vld_vec_16;
    reg [1:0] proc_dep_vld_vec_16_reg;
    wire [2:0] in_chan_dep_vld_vec_16;
    wire [98:0] in_chan_dep_data_vec_16;
    wire [2:0] token_in_vec_16;
    wire [1:0] out_chan_dep_vld_vec_16;
    wire [32:0] out_chan_dep_data_16;
    wire [1:0] token_out_vec_16;
    wire dl_detect_out_16;
    wire dep_chan_vld_14_16;
    wire [32:0] dep_chan_data_14_16;
    wire token_14_16;
    wire dep_chan_vld_17_16;
    wire [32:0] dep_chan_data_17_16;
    wire token_17_16;
    wire dep_chan_vld_20_16;
    wire [32:0] dep_chan_data_20_16;
    wire token_20_16;
    wire [2:0] proc_17_data_FIFO_blk;
    wire [2:0] proc_17_data_PIPO_blk;
    wire [2:0] proc_17_start_FIFO_blk;
    wire [2:0] proc_17_TLF_FIFO_blk;
    wire [2:0] proc_17_input_sync_blk;
    wire [2:0] proc_17_output_sync_blk;
    wire [2:0] proc_dep_vld_vec_17;
    reg [2:0] proc_dep_vld_vec_17_reg;
    wire [2:0] in_chan_dep_vld_vec_17;
    wire [98:0] in_chan_dep_data_vec_17;
    wire [2:0] token_in_vec_17;
    wire [2:0] out_chan_dep_vld_vec_17;
    wire [32:0] out_chan_dep_data_17;
    wire [2:0] token_out_vec_17;
    wire dl_detect_out_17;
    wire dep_chan_vld_14_17;
    wire [32:0] dep_chan_data_14_17;
    wire token_14_17;
    wire dep_chan_vld_18_17;
    wire [32:0] dep_chan_data_18_17;
    wire token_18_17;
    wire dep_chan_vld_20_17;
    wire [32:0] dep_chan_data_20_17;
    wire token_20_17;
    wire [0:0] proc_18_data_FIFO_blk;
    wire [0:0] proc_18_data_PIPO_blk;
    wire [0:0] proc_18_start_FIFO_blk;
    wire [0:0] proc_18_TLF_FIFO_blk;
    wire [0:0] proc_18_input_sync_blk;
    wire [0:0] proc_18_output_sync_blk;
    wire [0:0] proc_dep_vld_vec_18;
    reg [0:0] proc_dep_vld_vec_18_reg;
    wire [0:0] in_chan_dep_vld_vec_18;
    wire [32:0] in_chan_dep_data_vec_18;
    wire [0:0] token_in_vec_18;
    wire [0:0] out_chan_dep_vld_vec_18;
    wire [32:0] out_chan_dep_data_18;
    wire [0:0] token_out_vec_18;
    wire dl_detect_out_18;
    wire dep_chan_vld_19_18;
    wire [32:0] dep_chan_data_19_18;
    wire token_19_18;
    wire [4:0] proc_19_data_FIFO_blk;
    wire [4:0] proc_19_data_PIPO_blk;
    wire [4:0] proc_19_start_FIFO_blk;
    wire [4:0] proc_19_TLF_FIFO_blk;
    wire [4:0] proc_19_input_sync_blk;
    wire [4:0] proc_19_output_sync_blk;
    wire [4:0] proc_dep_vld_vec_19;
    reg [4:0] proc_dep_vld_vec_19_reg;
    wire [3:0] in_chan_dep_vld_vec_19;
    wire [131:0] in_chan_dep_data_vec_19;
    wire [3:0] token_in_vec_19;
    wire [4:0] out_chan_dep_vld_vec_19;
    wire [32:0] out_chan_dep_data_19;
    wire [4:0] token_out_vec_19;
    wire dl_detect_out_19;
    wire dep_chan_vld_13_19;
    wire [32:0] dep_chan_data_13_19;
    wire token_13_19;
    wire dep_chan_vld_14_19;
    wire [32:0] dep_chan_data_14_19;
    wire token_14_19;
    wire dep_chan_vld_15_19;
    wire [32:0] dep_chan_data_15_19;
    wire token_15_19;
    wire dep_chan_vld_20_19;
    wire [32:0] dep_chan_data_20_19;
    wire token_20_19;
    wire [3:0] proc_20_data_FIFO_blk;
    wire [3:0] proc_20_data_PIPO_blk;
    wire [3:0] proc_20_start_FIFO_blk;
    wire [3:0] proc_20_TLF_FIFO_blk;
    wire [3:0] proc_20_input_sync_blk;
    wire [3:0] proc_20_output_sync_blk;
    wire [3:0] proc_dep_vld_vec_20;
    reg [3:0] proc_dep_vld_vec_20_reg;
    wire [3:0] in_chan_dep_vld_vec_20;
    wire [131:0] in_chan_dep_data_vec_20;
    wire [3:0] token_in_vec_20;
    wire [3:0] out_chan_dep_vld_vec_20;
    wire [32:0] out_chan_dep_data_20;
    wire [3:0] token_out_vec_20;
    wire dl_detect_out_20;
    wire dep_chan_vld_15_20;
    wire [32:0] dep_chan_data_15_20;
    wire token_15_20;
    wire dep_chan_vld_16_20;
    wire [32:0] dep_chan_data_16_20;
    wire token_16_20;
    wire dep_chan_vld_17_20;
    wire [32:0] dep_chan_data_17_20;
    wire token_17_20;
    wire dep_chan_vld_19_20;
    wire [32:0] dep_chan_data_19_20;
    wire token_19_20;
    wire [2:0] proc_21_data_FIFO_blk;
    wire [2:0] proc_21_data_PIPO_blk;
    wire [2:0] proc_21_start_FIFO_blk;
    wire [2:0] proc_21_TLF_FIFO_blk;
    wire [2:0] proc_21_input_sync_blk;
    wire [2:0] proc_21_output_sync_blk;
    wire [2:0] proc_dep_vld_vec_21;
    reg [2:0] proc_dep_vld_vec_21_reg;
    wire [2:0] in_chan_dep_vld_vec_21;
    wire [98:0] in_chan_dep_data_vec_21;
    wire [2:0] token_in_vec_21;
    wire [2:0] out_chan_dep_vld_vec_21;
    wire [32:0] out_chan_dep_data_21;
    wire [2:0] token_out_vec_21;
    wire dl_detect_out_21;
    wire dep_chan_vld_2_21;
    wire [32:0] dep_chan_data_2_21;
    wire token_2_21;
    wire dep_chan_vld_12_21;
    wire [32:0] dep_chan_data_12_21;
    wire token_12_21;
    wire dep_chan_vld_22_21;
    wire [32:0] dep_chan_data_22_21;
    wire token_22_21;
    wire [2:0] proc_22_data_FIFO_blk;
    wire [2:0] proc_22_data_PIPO_blk;
    wire [2:0] proc_22_start_FIFO_blk;
    wire [2:0] proc_22_TLF_FIFO_blk;
    wire [2:0] proc_22_input_sync_blk;
    wire [2:0] proc_22_output_sync_blk;
    wire [2:0] proc_dep_vld_vec_22;
    reg [2:0] proc_dep_vld_vec_22_reg;
    wire [2:0] in_chan_dep_vld_vec_22;
    wire [98:0] in_chan_dep_data_vec_22;
    wire [2:0] token_in_vec_22;
    wire [2:0] out_chan_dep_vld_vec_22;
    wire [32:0] out_chan_dep_data_22;
    wire [2:0] token_out_vec_22;
    wire dl_detect_out_22;
    wire dep_chan_vld_1_22;
    wire [32:0] dep_chan_data_1_22;
    wire token_1_22;
    wire dep_chan_vld_21_22;
    wire [32:0] dep_chan_data_21_22;
    wire token_21_22;
    wire dep_chan_vld_23_22;
    wire [32:0] dep_chan_data_23_22;
    wire token_23_22;
    wire [4:0] proc_23_data_FIFO_blk;
    wire [4:0] proc_23_data_PIPO_blk;
    wire [4:0] proc_23_start_FIFO_blk;
    wire [4:0] proc_23_TLF_FIFO_blk;
    wire [4:0] proc_23_input_sync_blk;
    wire [4:0] proc_23_output_sync_blk;
    wire [4:0] proc_dep_vld_vec_23;
    reg [4:0] proc_dep_vld_vec_23_reg;
    wire [4:0] in_chan_dep_vld_vec_23;
    wire [164:0] in_chan_dep_data_vec_23;
    wire [4:0] token_in_vec_23;
    wire [4:0] out_chan_dep_vld_vec_23;
    wire [32:0] out_chan_dep_data_23;
    wire [4:0] token_out_vec_23;
    wire dl_detect_out_23;
    wire dep_chan_vld_0_23;
    wire [32:0] dep_chan_data_0_23;
    wire token_0_23;
    wire dep_chan_vld_2_23;
    wire [32:0] dep_chan_data_2_23;
    wire token_2_23;
    wire dep_chan_vld_12_23;
    wire [32:0] dep_chan_data_12_23;
    wire token_12_23;
    wire dep_chan_vld_22_23;
    wire [32:0] dep_chan_data_22_23;
    wire token_22_23;
    wire dep_chan_vld_24_23;
    wire [32:0] dep_chan_data_24_23;
    wire token_24_23;
    wire [2:0] proc_24_data_FIFO_blk;
    wire [2:0] proc_24_data_PIPO_blk;
    wire [2:0] proc_24_start_FIFO_blk;
    wire [2:0] proc_24_TLF_FIFO_blk;
    wire [2:0] proc_24_input_sync_blk;
    wire [2:0] proc_24_output_sync_blk;
    wire [2:0] proc_dep_vld_vec_24;
    reg [2:0] proc_dep_vld_vec_24_reg;
    wire [2:0] in_chan_dep_vld_vec_24;
    wire [98:0] in_chan_dep_data_vec_24;
    wire [2:0] token_in_vec_24;
    wire [2:0] out_chan_dep_vld_vec_24;
    wire [32:0] out_chan_dep_data_24;
    wire [2:0] token_out_vec_24;
    wire dl_detect_out_24;
    wire dep_chan_vld_0_24;
    wire [32:0] dep_chan_data_0_24;
    wire token_0_24;
    wire dep_chan_vld_1_24;
    wire [32:0] dep_chan_data_1_24;
    wire token_1_24;
    wire dep_chan_vld_23_24;
    wire [32:0] dep_chan_data_23_24;
    wire token_23_24;
    wire [3:0] proc_25_data_FIFO_blk;
    wire [3:0] proc_25_data_PIPO_blk;
    wire [3:0] proc_25_start_FIFO_blk;
    wire [3:0] proc_25_TLF_FIFO_blk;
    wire [3:0] proc_25_input_sync_blk;
    wire [3:0] proc_25_output_sync_blk;
    wire [3:0] proc_dep_vld_vec_25;
    reg [3:0] proc_dep_vld_vec_25_reg;
    wire [3:0] in_chan_dep_vld_vec_25;
    wire [131:0] in_chan_dep_data_vec_25;
    wire [3:0] token_in_vec_25;
    wire [3:0] out_chan_dep_vld_vec_25;
    wire [32:0] out_chan_dep_data_25;
    wire [3:0] token_out_vec_25;
    wire dl_detect_out_25;
    wire dep_chan_vld_26_25;
    wire [32:0] dep_chan_data_26_25;
    wire token_26_25;
    wire dep_chan_vld_29_25;
    wire [32:0] dep_chan_data_29_25;
    wire token_29_25;
    wire dep_chan_vld_30_25;
    wire [32:0] dep_chan_data_30_25;
    wire token_30_25;
    wire dep_chan_vld_32_25;
    wire [32:0] dep_chan_data_32_25;
    wire token_32_25;
    wire [0:0] proc_26_data_FIFO_blk;
    wire [0:0] proc_26_data_PIPO_blk;
    wire [0:0] proc_26_start_FIFO_blk;
    wire [0:0] proc_26_TLF_FIFO_blk;
    wire [0:0] proc_26_input_sync_blk;
    wire [0:0] proc_26_output_sync_blk;
    wire [0:0] proc_dep_vld_vec_26;
    reg [0:0] proc_dep_vld_vec_26_reg;
    wire [1:0] in_chan_dep_vld_vec_26;
    wire [65:0] in_chan_dep_data_vec_26;
    wire [1:0] token_in_vec_26;
    wire [0:0] out_chan_dep_vld_vec_26;
    wire [32:0] out_chan_dep_data_26;
    wire [0:0] token_out_vec_26;
    wire dl_detect_out_26;
    wire dep_chan_vld_25_26;
    wire [32:0] dep_chan_data_25_26;
    wire token_25_26;
    wire dep_chan_vld_27_26;
    wire [32:0] dep_chan_data_27_26;
    wire token_27_26;
    wire [0:0] proc_27_data_FIFO_blk;
    wire [0:0] proc_27_data_PIPO_blk;
    wire [0:0] proc_27_start_FIFO_blk;
    wire [0:0] proc_27_TLF_FIFO_blk;
    wire [0:0] proc_27_input_sync_blk;
    wire [0:0] proc_27_output_sync_blk;
    wire [0:0] proc_dep_vld_vec_27;
    reg [0:0] proc_dep_vld_vec_27_reg;
    wire [0:0] in_chan_dep_vld_vec_27;
    wire [32:0] in_chan_dep_data_vec_27;
    wire [0:0] token_in_vec_27;
    wire [0:0] out_chan_dep_vld_vec_27;
    wire [32:0] out_chan_dep_data_27;
    wire [0:0] token_out_vec_27;
    wire dl_detect_out_27;
    wire dep_chan_vld_28_27;
    wire [32:0] dep_chan_data_28_27;
    wire token_28_27;
    wire [0:0] proc_28_data_FIFO_blk;
    wire [0:0] proc_28_data_PIPO_blk;
    wire [0:0] proc_28_start_FIFO_blk;
    wire [0:0] proc_28_TLF_FIFO_blk;
    wire [0:0] proc_28_input_sync_blk;
    wire [0:0] proc_28_output_sync_blk;
    wire [0:0] proc_dep_vld_vec_28;
    reg [0:0] proc_dep_vld_vec_28_reg;
    wire [0:0] in_chan_dep_vld_vec_28;
    wire [32:0] in_chan_dep_data_vec_28;
    wire [0:0] token_in_vec_28;
    wire [0:0] out_chan_dep_vld_vec_28;
    wire [32:0] out_chan_dep_data_28;
    wire [0:0] token_out_vec_28;
    wire dl_detect_out_28;
    wire dep_chan_vld_32_28;
    wire [32:0] dep_chan_data_32_28;
    wire token_32_28;
    wire [1:0] proc_29_data_FIFO_blk;
    wire [1:0] proc_29_data_PIPO_blk;
    wire [1:0] proc_29_start_FIFO_blk;
    wire [1:0] proc_29_TLF_FIFO_blk;
    wire [1:0] proc_29_input_sync_blk;
    wire [1:0] proc_29_output_sync_blk;
    wire [1:0] proc_dep_vld_vec_29;
    reg [1:0] proc_dep_vld_vec_29_reg;
    wire [0:0] in_chan_dep_vld_vec_29;
    wire [32:0] in_chan_dep_data_vec_29;
    wire [0:0] token_in_vec_29;
    wire [1:0] out_chan_dep_vld_vec_29;
    wire [32:0] out_chan_dep_data_29;
    wire [1:0] token_out_vec_29;
    wire dl_detect_out_29;
    wire dep_chan_vld_25_29;
    wire [32:0] dep_chan_data_25_29;
    wire token_25_29;
    wire [1:0] proc_30_data_FIFO_blk;
    wire [1:0] proc_30_data_PIPO_blk;
    wire [1:0] proc_30_start_FIFO_blk;
    wire [1:0] proc_30_TLF_FIFO_blk;
    wire [1:0] proc_30_input_sync_blk;
    wire [1:0] proc_30_output_sync_blk;
    wire [1:0] proc_dep_vld_vec_30;
    reg [1:0] proc_dep_vld_vec_30_reg;
    wire [1:0] in_chan_dep_vld_vec_30;
    wire [65:0] in_chan_dep_data_vec_30;
    wire [1:0] token_in_vec_30;
    wire [1:0] out_chan_dep_vld_vec_30;
    wire [32:0] out_chan_dep_data_30;
    wire [1:0] token_out_vec_30;
    wire dl_detect_out_30;
    wire dep_chan_vld_25_30;
    wire [32:0] dep_chan_data_25_30;
    wire token_25_30;
    wire dep_chan_vld_31_30;
    wire [32:0] dep_chan_data_31_30;
    wire token_31_30;
    wire [1:0] proc_31_data_FIFO_blk;
    wire [1:0] proc_31_data_PIPO_blk;
    wire [1:0] proc_31_start_FIFO_blk;
    wire [1:0] proc_31_TLF_FIFO_blk;
    wire [1:0] proc_31_input_sync_blk;
    wire [1:0] proc_31_output_sync_blk;
    wire [1:0] proc_dep_vld_vec_31;
    reg [1:0] proc_dep_vld_vec_31_reg;
    wire [1:0] in_chan_dep_vld_vec_31;
    wire [65:0] in_chan_dep_data_vec_31;
    wire [1:0] token_in_vec_31;
    wire [1:0] out_chan_dep_vld_vec_31;
    wire [32:0] out_chan_dep_data_31;
    wire [1:0] token_out_vec_31;
    wire dl_detect_out_31;
    wire dep_chan_vld_30_31;
    wire [32:0] dep_chan_data_30_31;
    wire token_30_31;
    wire dep_chan_vld_32_31;
    wire [32:0] dep_chan_data_32_31;
    wire token_32_31;
    wire [2:0] proc_32_data_FIFO_blk;
    wire [2:0] proc_32_data_PIPO_blk;
    wire [2:0] proc_32_start_FIFO_blk;
    wire [2:0] proc_32_TLF_FIFO_blk;
    wire [2:0] proc_32_input_sync_blk;
    wire [2:0] proc_32_output_sync_blk;
    wire [2:0] proc_dep_vld_vec_32;
    reg [2:0] proc_dep_vld_vec_32_reg;
    wire [2:0] in_chan_dep_vld_vec_32;
    wire [98:0] in_chan_dep_data_vec_32;
    wire [2:0] token_in_vec_32;
    wire [2:0] out_chan_dep_vld_vec_32;
    wire [32:0] out_chan_dep_data_32;
    wire [2:0] token_out_vec_32;
    wire dl_detect_out_32;
    wire dep_chan_vld_25_32;
    wire [32:0] dep_chan_data_25_32;
    wire token_25_32;
    wire dep_chan_vld_29_32;
    wire [32:0] dep_chan_data_29_32;
    wire token_29_32;
    wire dep_chan_vld_31_32;
    wire [32:0] dep_chan_data_31_32;
    wire token_31_32;
    wire [32:0] dl_in_vec;
    wire dl_detect_out;
    wire token_clear;
    reg [32:0] origin;

    reg ap_done_reg_0;// for module Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.addrbound_2_U0
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_0 <= 'b0;
        end
        else begin
            ap_done_reg_0 <= Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.addrbound_2_U0.ap_done & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.addrbound_2_U0.ap_continue;
        end
    end

    reg ap_done_reg_1;// for module Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split48_proc_U0
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_1 <= 'b0;
        end
        else begin
            ap_done_reg_1 <= Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split48_proc_U0.ap_done & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split48_proc_U0.ap_continue;
        end
    end

    reg ap_done_reg_2;// for module Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2AxiStream_1_U0
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_2 <= 'b0;
        end
        else begin
            ap_done_reg_2 <= Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2AxiStream_1_U0.ap_done & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2AxiStream_1_U0.ap_continue;
        end
    end

    reg ap_done_reg_3;// for module Array2xfMat_64_6_1080_1920_1_U0
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_3 <= 'b0;
        end
        else begin
            ap_done_reg_3 <= Array2xfMat_64_6_1080_1920_1_U0.ap_done & ~Array2xfMat_64_6_1080_1920_1_U0.ap_continue;
        end
    end

    reg ap_done_reg_4;// for module Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.addrbound_1_U0
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_4 <= 'b0;
        end
        else begin
            ap_done_reg_4 <= Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.addrbound_1_U0.ap_done & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.addrbound_1_U0.ap_continue;
        end
    end

    reg ap_done_reg_5;// for module Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split37_proc_U0
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_5 <= 'b0;
        end
        else begin
            ap_done_reg_5 <= Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split37_proc_U0.ap_done & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split37_proc_U0.ap_continue;
        end
    end

    reg ap_done_reg_6;// for module Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2AxiStream_U0
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_6 <= 'b0;
        end
        else begin
            ap_done_reg_6 <= Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2AxiStream_U0.ap_done & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2AxiStream_U0.ap_continue;
        end
    end

    reg ap_done_reg_7;// for module xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.addrbound_U0
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_7 <= 'b0;
        end
        else begin
            ap_done_reg_7 <= xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.addrbound_U0.ap_done & ~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.addrbound_U0.ap_continue;
        end
    end

    reg ap_done_reg_8;// for module xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split24_proc_U0
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_8 <= 'b0;
        end
        else begin
            ap_done_reg_8 <= xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split24_proc_U0.ap_done & ~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split24_proc_U0.ap_continue;
        end
    end

    reg ap_done_reg_9;// for module xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.MatStream2AxiStream_U0
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_9 <= 'b0;
        end
        else begin
            ap_done_reg_9 <= xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.MatStream2AxiStream_U0.ap_done & ~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.MatStream2AxiStream_U0.ap_continue;
        end
    end

    reg ap_done_reg_10;// for module xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.AxiStream2Axi_U0
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_10 <= 'b0;
        end
        else begin
            ap_done_reg_10 <= xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.AxiStream2Axi_U0.ap_done & ~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.AxiStream2Axi_U0.ap_continue;
        end
    end

reg [15:0] trans_in_cnt_0;// for process pp_pipeline_accel_entry33_U0
always @(negedge reset or posedge clock) begin
    if (~reset) begin
         trans_in_cnt_0 <= 16'h0;
    end
    else if (pp_pipeline_accel_entry33_U0.start_write == 1'b1) begin
        trans_in_cnt_0 <= trans_in_cnt_0 + 16'h1;
    end
    else begin
        trans_in_cnt_0 <= trans_in_cnt_0;
    end
end

reg [15:0] trans_out_cnt_0;// for process pp_pipeline_accel_entry33_U0
always @(negedge reset or posedge clock) begin
    if (~reset) begin
         trans_out_cnt_0 <= 16'h0;
    end
    else if (pp_pipeline_accel_entry33_U0.ap_done == 1'b1 && pp_pipeline_accel_entry33_U0.ap_continue == 1'b1) begin
        trans_out_cnt_0 <= trans_out_cnt_0 + 16'h1;
    end
    else begin
        trans_out_cnt_0 <= trans_out_cnt_0;
    end
end

reg [15:0] trans_in_cnt_1;// for process Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0
always @(negedge reset or posedge clock) begin
    if (~reset) begin
         trans_in_cnt_1 <= 16'h0;
    end
    else if (Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0.start_write == 1'b1) begin
        trans_in_cnt_1 <= trans_in_cnt_1 + 16'h1;
    end
    else begin
        trans_in_cnt_1 <= trans_in_cnt_1;
    end
end

reg [15:0] trans_out_cnt_1;// for process Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0
always @(negedge reset or posedge clock) begin
    if (~reset) begin
         trans_out_cnt_1 <= 16'h0;
    end
    else if (Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0.ap_done == 1'b1 && Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0.ap_continue == 1'b1) begin
        trans_out_cnt_1 <= trans_out_cnt_1 + 16'h1;
    end
    else begin
        trans_out_cnt_1 <= trans_out_cnt_1;
    end
end

reg [15:0] trans_in_cnt_2;// for process Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0
always @(negedge reset or posedge clock) begin
    if (~reset) begin
         trans_in_cnt_2 <= 16'h0;
    end
    else if (Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0.start_write == 1'b1) begin
        trans_in_cnt_2 <= trans_in_cnt_2 + 16'h1;
    end
    else begin
        trans_in_cnt_2 <= trans_in_cnt_2;
    end
end

reg [15:0] trans_out_cnt_2;// for process Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0
always @(negedge reset or posedge clock) begin
    if (~reset) begin
         trans_out_cnt_2 <= 16'h0;
    end
    else if (Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0.ap_done == 1'b1 && Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0.ap_continue == 1'b1) begin
        trans_out_cnt_2 <= trans_out_cnt_2 + 16'h1;
    end
    else begin
        trans_out_cnt_2 <= trans_out_cnt_2;
    end
end

reg [15:0] trans_in_cnt_3;// for process Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_pxl_width_1_U0
always @(negedge reset or posedge clock) begin
    if (~reset) begin
         trans_in_cnt_3 <= 16'h0;
    end
    else if (Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_pxl_width_1_U0.start_write == 1'b1) begin
        trans_in_cnt_3 <= trans_in_cnt_3 + 16'h1;
    end
    else begin
        trans_in_cnt_3 <= trans_in_cnt_3;
    end
end

reg [15:0] trans_out_cnt_3;// for process Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_pxl_width_1_U0
always @(negedge reset or posedge clock) begin
    if (~reset) begin
         trans_out_cnt_3 <= 16'h0;
    end
    else if (Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_pxl_width_1_U0.ap_done == 1'b1 && Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_pxl_width_1_U0.ap_continue == 1'b1) begin
        trans_out_cnt_3 <= trans_out_cnt_3 + 16'h1;
    end
    else begin
        trans_out_cnt_3 <= trans_out_cnt_3;
    end
end

reg [15:0] trans_in_cnt_4;// for process Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0
always @(negedge reset or posedge clock) begin
    if (~reset) begin
         trans_in_cnt_4 <= 16'h0;
    end
    else if (Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0.start_write == 1'b1) begin
        trans_in_cnt_4 <= trans_in_cnt_4 + 16'h1;
    end
    else begin
        trans_in_cnt_4 <= trans_in_cnt_4;
    end
end

reg [15:0] trans_out_cnt_4;// for process Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0
always @(negedge reset or posedge clock) begin
    if (~reset) begin
         trans_out_cnt_4 <= 16'h0;
    end
    else if (Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0.ap_done == 1'b1 && Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0.ap_continue == 1'b1) begin
        trans_out_cnt_4 <= trans_out_cnt_4 + 16'h1;
    end
    else begin
        trans_out_cnt_4 <= trans_out_cnt_4;
    end
end

reg [15:0] trans_in_cnt_5;// for process Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0
always @(negedge reset or posedge clock) begin
    if (~reset) begin
         trans_in_cnt_5 <= 16'h0;
    end
    else if (Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0.start_write == 1'b1) begin
        trans_in_cnt_5 <= trans_in_cnt_5 + 16'h1;
    end
    else begin
        trans_in_cnt_5 <= trans_in_cnt_5;
    end
end

reg [15:0] trans_out_cnt_5;// for process Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0
always @(negedge reset or posedge clock) begin
    if (~reset) begin
         trans_out_cnt_5 <= 16'h0;
    end
    else if (Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0.ap_done == 1'b1 && Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0.ap_continue == 1'b1) begin
        trans_out_cnt_5 <= trans_out_cnt_5 + 16'h1;
    end
    else begin
        trans_out_cnt_5 <= trans_out_cnt_5;
    end
end

reg [15:0] trans_in_cnt_6;// for process Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_pxl_width_U0
always @(negedge reset or posedge clock) begin
    if (~reset) begin
         trans_in_cnt_6 <= 16'h0;
    end
    else if (Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_pxl_width_U0.start_write == 1'b1) begin
        trans_in_cnt_6 <= trans_in_cnt_6 + 16'h1;
    end
    else begin
        trans_in_cnt_6 <= trans_in_cnt_6;
    end
end

reg [15:0] trans_out_cnt_6;// for process Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_pxl_width_U0
always @(negedge reset or posedge clock) begin
    if (~reset) begin
         trans_out_cnt_6 <= 16'h0;
    end
    else if (Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_pxl_width_U0.ap_done == 1'b1 && Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_pxl_width_U0.ap_continue == 1'b1) begin
        trans_out_cnt_6 <= trans_out_cnt_6 + 16'h1;
    end
    else begin
        trans_out_cnt_6 <= trans_out_cnt_6;
    end
end

reg [15:0] trans_in_cnt_7;// for process Array2xfMat_64_0_2160_3840_1_U0
always @(negedge reset or posedge clock) begin
    if (~reset) begin
         trans_in_cnt_7 <= 16'h0;
    end
    else if (Array2xfMat_64_0_2160_3840_1_U0.start_write == 1'b1) begin
        trans_in_cnt_7 <= trans_in_cnt_7 + 16'h1;
    end
    else begin
        trans_in_cnt_7 <= trans_in_cnt_7;
    end
end

reg [15:0] trans_out_cnt_7;// for process Array2xfMat_64_0_2160_3840_1_U0
always @(negedge reset or posedge clock) begin
    if (~reset) begin
         trans_out_cnt_7 <= 16'h0;
    end
    else if (Array2xfMat_64_0_2160_3840_1_U0.ap_done == 1'b1 && Array2xfMat_64_0_2160_3840_1_U0.ap_continue == 1'b1) begin
        trans_out_cnt_7 <= trans_out_cnt_7 + 16'h1;
    end
    else begin
        trans_out_cnt_7 <= trans_out_cnt_7;
    end
end

reg [15:0] trans_in_cnt_8;// for process Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0
always @(negedge reset or posedge clock) begin
    if (~reset) begin
         trans_in_cnt_8 <= 16'h0;
    end
    else if (Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.start_write == 1'b1) begin
        trans_in_cnt_8 <= trans_in_cnt_8 + 16'h1;
    end
    else begin
        trans_in_cnt_8 <= trans_in_cnt_8;
    end
end

reg [15:0] trans_out_cnt_8;// for process Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0
always @(negedge reset or posedge clock) begin
    if (~reset) begin
         trans_out_cnt_8 <= 16'h0;
    end
    else if (Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.ap_done == 1'b1 && Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.ap_continue == 1'b1) begin
        trans_out_cnt_8 <= trans_out_cnt_8 + 16'h1;
    end
    else begin
        trans_out_cnt_8 <= trans_out_cnt_8;
    end
end

reg [15:0] trans_in_cnt_9;// for process xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0
always @(negedge reset or posedge clock) begin
    if (~reset) begin
         trans_in_cnt_9 <= 16'h0;
    end
    else if (xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0.start_write == 1'b1) begin
        trans_in_cnt_9 <= trans_in_cnt_9 + 16'h1;
    end
    else begin
        trans_in_cnt_9 <= trans_in_cnt_9;
    end
end

reg [15:0] trans_out_cnt_9;// for process xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0
always @(negedge reset or posedge clock) begin
    if (~reset) begin
         trans_out_cnt_9 <= 16'h0;
    end
    else if (xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0.ap_done == 1'b1 && xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0.ap_continue == 1'b1) begin
        trans_out_cnt_9 <= trans_out_cnt_9 + 16'h1;
    end
    else begin
        trans_out_cnt_9 <= trans_out_cnt_9;
    end
end

    // Process: pp_pipeline_accel_entry33_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 0, 6, 6) pp_pipeline_accel_hls_deadlock_detect_unit_0 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_0),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_0),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_0),
        .token_in_vec(token_in_vec_0),
        .dl_detect_in(dl_detect_out),
        .origin(origin[0]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_0),
        .out_chan_dep_data(out_chan_dep_data_0),
        .token_out_vec(token_out_vec_0),
        .dl_detect_out(dl_in_vec[0]));

    assign proc_0_data_FIFO_blk[0] = 1'b0 | (~pp_pipeline_accel_entry33_U0.img_inp_y_out_blk_n) | (~pp_pipeline_accel_entry33_U0.in_img_linestride_out_blk_n);
    assign proc_0_data_PIPO_blk[0] = 1'b0;
    assign proc_0_start_FIFO_blk[0] = 1'b0;
    assign proc_0_TLF_FIFO_blk[0] = 1'b0;
    assign proc_0_input_sync_blk[0] = 1'b0 | (ap_sync_pp_pipeline_accel_entry33_U0_ap_ready & pp_pipeline_accel_entry33_U0.ap_idle & ~ap_sync_Array2xfMat_64_0_2160_3840_1_U0_ap_ready);
    assign proc_0_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_0[0] = dl_detect_out ? proc_dep_vld_vec_0_reg[0] : (proc_0_data_FIFO_blk[0] | proc_0_data_PIPO_blk[0] | proc_0_start_FIFO_blk[0] | proc_0_TLF_FIFO_blk[0] | proc_0_input_sync_blk[0] | proc_0_output_sync_blk[0]);
    assign proc_0_data_FIFO_blk[1] = 1'b0 | (~pp_pipeline_accel_entry33_U0.img_inp_uv_out_blk_n);
    assign proc_0_data_PIPO_blk[1] = 1'b0;
    assign proc_0_start_FIFO_blk[1] = 1'b0;
    assign proc_0_TLF_FIFO_blk[1] = 1'b0;
    assign proc_0_input_sync_blk[1] = 1'b0 | (ap_sync_pp_pipeline_accel_entry33_U0_ap_ready & pp_pipeline_accel_entry33_U0.ap_idle & ~ap_sync_Array2xfMat_64_6_1080_1920_1_U0_ap_ready);
    assign proc_0_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_0[1] = dl_detect_out ? proc_dep_vld_vec_0_reg[1] : (proc_0_data_FIFO_blk[1] | proc_0_data_PIPO_blk[1] | proc_0_start_FIFO_blk[1] | proc_0_TLF_FIFO_blk[1] | proc_0_input_sync_blk[1] | proc_0_output_sync_blk[1]);
    assign proc_0_data_FIFO_blk[2] = 1'b0 | (~pp_pipeline_accel_entry33_U0.img_out_out_blk_n) | (~pp_pipeline_accel_entry33_U0.out_img_linestride_out_blk_n);
    assign proc_0_data_PIPO_blk[2] = 1'b0;
    assign proc_0_start_FIFO_blk[2] = 1'b0 | (~start_for_xfMat2Array_64_9_720_720_1_1_U0_U.if_full_n & pp_pipeline_accel_entry33_U0.ap_start & ~pp_pipeline_accel_entry33_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_xfMat2Array_64_9_720_720_1_1_U0_U.if_read);
    assign proc_0_TLF_FIFO_blk[2] = 1'b0;
    assign proc_0_input_sync_blk[2] = 1'b0;
    assign proc_0_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_0[2] = dl_detect_out ? proc_dep_vld_vec_0_reg[2] : (proc_0_data_FIFO_blk[2] | proc_0_data_PIPO_blk[2] | proc_0_start_FIFO_blk[2] | proc_0_TLF_FIFO_blk[2] | proc_0_input_sync_blk[2] | proc_0_output_sync_blk[2]);
    assign proc_0_data_FIFO_blk[3] = 1'b0 | (~pp_pipeline_accel_entry33_U0.params_out_blk_n);
    assign proc_0_data_PIPO_blk[3] = 1'b0;
    assign proc_0_start_FIFO_blk[3] = 1'b0;
    assign proc_0_TLF_FIFO_blk[3] = 1'b0;
    assign proc_0_input_sync_blk[3] = 1'b0 | (ap_sync_pp_pipeline_accel_entry33_U0_ap_ready & pp_pipeline_accel_entry33_U0.ap_idle & ~ap_sync_preProcess_9_9_720_720_1_8_8_8_4_8_8_U0_ap_ready);
    assign proc_0_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_0[3] = dl_detect_out ? proc_dep_vld_vec_0_reg[3] : (proc_0_data_FIFO_blk[3] | proc_0_data_PIPO_blk[3] | proc_0_start_FIFO_blk[3] | proc_0_TLF_FIFO_blk[3] | proc_0_input_sync_blk[3] | proc_0_output_sync_blk[3]);
    assign proc_0_data_FIFO_blk[4] = 1'b0 | (~pp_pipeline_accel_entry33_U0.in_img_width_out_blk_n) | (~pp_pipeline_accel_entry33_U0.in_img_height_out_blk_n) | (~pp_pipeline_accel_entry33_U0.out_img_width_out_blk_n) | (~pp_pipeline_accel_entry33_U0.out_img_height_out_blk_n);
    assign proc_0_data_PIPO_blk[4] = 1'b0;
    assign proc_0_start_FIFO_blk[4] = 1'b0 | (~start_for_Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0_U.if_full_n & pp_pipeline_accel_entry33_U0.ap_start & ~pp_pipeline_accel_entry33_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0_U.if_read);
    assign proc_0_TLF_FIFO_blk[4] = 1'b0;
    assign proc_0_input_sync_blk[4] = 1'b0;
    assign proc_0_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_0[4] = dl_detect_out ? proc_dep_vld_vec_0_reg[4] : (proc_0_data_FIFO_blk[4] | proc_0_data_PIPO_blk[4] | proc_0_start_FIFO_blk[4] | proc_0_TLF_FIFO_blk[4] | proc_0_input_sync_blk[4] | proc_0_output_sync_blk[4]);
    assign proc_0_data_FIFO_blk[5] = 1'b0 | (~pp_pipeline_accel_entry33_U0.in_img_linestride_out1_blk_n);
    assign proc_0_data_PIPO_blk[5] = 1'b0;
    assign proc_0_start_FIFO_blk[5] = 1'b0 | (~start_for_Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit2022_proc_U0_U.if_full_n & pp_pipeline_accel_entry33_U0.ap_start & ~pp_pipeline_accel_entry33_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit2022_proc_U0_U.if_read);
    assign proc_0_TLF_FIFO_blk[5] = 1'b0;
    assign proc_0_input_sync_blk[5] = 1'b0;
    assign proc_0_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_0[5] = dl_detect_out ? proc_dep_vld_vec_0_reg[5] : (proc_0_data_FIFO_blk[5] | proc_0_data_PIPO_blk[5] | proc_0_start_FIFO_blk[5] | proc_0_TLF_FIFO_blk[5] | proc_0_input_sync_blk[5] | proc_0_output_sync_blk[5]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_0_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_0_reg <= proc_dep_vld_vec_0;
        end
    end
    assign in_chan_dep_vld_vec_0[0] = dep_chan_vld_1_0;
    assign in_chan_dep_data_vec_0[32 : 0] = dep_chan_data_1_0;
    assign token_in_vec_0[0] = token_1_0;
    assign in_chan_dep_vld_vec_0[1] = dep_chan_vld_2_0;
    assign in_chan_dep_data_vec_0[65 : 33] = dep_chan_data_2_0;
    assign token_in_vec_0[1] = token_2_0;
    assign in_chan_dep_vld_vec_0[2] = dep_chan_vld_11_0;
    assign in_chan_dep_data_vec_0[98 : 66] = dep_chan_data_11_0;
    assign token_in_vec_0[2] = token_11_0;
    assign in_chan_dep_vld_vec_0[3] = dep_chan_vld_12_0;
    assign in_chan_dep_data_vec_0[131 : 99] = dep_chan_data_12_0;
    assign token_in_vec_0[3] = token_12_0;
    assign in_chan_dep_vld_vec_0[4] = dep_chan_vld_23_0;
    assign in_chan_dep_data_vec_0[164 : 132] = dep_chan_data_23_0;
    assign token_in_vec_0[4] = token_23_0;
    assign in_chan_dep_vld_vec_0[5] = dep_chan_vld_24_0;
    assign in_chan_dep_data_vec_0[197 : 165] = dep_chan_data_24_0;
    assign token_in_vec_0[5] = token_24_0;
    assign dep_chan_vld_0_2 = out_chan_dep_vld_vec_0[0];
    assign dep_chan_data_0_2 = out_chan_dep_data_0;
    assign token_0_2 = token_out_vec_0[0];
    assign dep_chan_vld_0_12 = out_chan_dep_vld_vec_0[1];
    assign dep_chan_data_0_12 = out_chan_dep_data_0;
    assign token_0_12 = token_out_vec_0[1];
    assign dep_chan_vld_0_24 = out_chan_dep_vld_vec_0[2];
    assign dep_chan_data_0_24 = out_chan_dep_data_0;
    assign token_0_24 = token_out_vec_0[2];
    assign dep_chan_vld_0_23 = out_chan_dep_vld_vec_0[3];
    assign dep_chan_data_0_23 = out_chan_dep_data_0;
    assign token_0_23 = token_out_vec_0[3];
    assign dep_chan_vld_0_1 = out_chan_dep_vld_vec_0[4];
    assign dep_chan_data_0_1 = out_chan_dep_data_0;
    assign token_0_1 = token_out_vec_0[4];
    assign dep_chan_vld_0_11 = out_chan_dep_vld_vec_0[5];
    assign dep_chan_data_0_11 = out_chan_dep_data_0;
    assign token_0_11 = token_out_vec_0[5];

    // Process: Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 1, 5, 4) pp_pipeline_accel_hls_deadlock_detect_unit_1 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_1),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_1),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_1),
        .token_in_vec(token_in_vec_1),
        .dl_detect_in(dl_detect_out),
        .origin(origin[1]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_1),
        .out_chan_dep_data(out_chan_dep_data_1),
        .token_out_vec(token_out_vec_1),
        .dl_detect_out(dl_in_vec[1]));

    assign proc_1_data_FIFO_blk[0] = 1'b0 | (~Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.in_img_height_blk_n) | (~Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.in_img_width_blk_n) | (~Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.out_img_height_blk_n) | (~Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.out_img_width_blk_n);
    assign proc_1_data_PIPO_blk[0] = 1'b0;
    assign proc_1_start_FIFO_blk[0] = 1'b0 | (~start_for_Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0_U.if_empty_n & Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.ap_idle & ~start_for_Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0_U.if_write);
    assign proc_1_TLF_FIFO_blk[0] = 1'b0;
    assign proc_1_input_sync_blk[0] = 1'b0;
    assign proc_1_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_1[0] = dl_detect_out ? proc_dep_vld_vec_1_reg[0] : (proc_1_data_FIFO_blk[0] | proc_1_data_PIPO_blk[0] | proc_1_start_FIFO_blk[0] | proc_1_TLF_FIFO_blk[0] | proc_1_input_sync_blk[0] | proc_1_output_sync_blk[0]);
    assign proc_1_data_FIFO_blk[1] = 1'b0 | (~Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.imgInput_y_rows_out_blk_n) | (~Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.imgInput_y_cols_out_blk_n);
    assign proc_1_data_PIPO_blk[1] = 1'b0;
    assign proc_1_start_FIFO_blk[1] = 1'b0;
    assign proc_1_TLF_FIFO_blk[1] = 1'b0;
    assign proc_1_input_sync_blk[1] = 1'b0;
    assign proc_1_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_1[1] = dl_detect_out ? proc_dep_vld_vec_1_reg[1] : (proc_1_data_FIFO_blk[1] | proc_1_data_PIPO_blk[1] | proc_1_start_FIFO_blk[1] | proc_1_TLF_FIFO_blk[1] | proc_1_input_sync_blk[1] | proc_1_output_sync_blk[1]);
    assign proc_1_data_FIFO_blk[2] = 1'b0 | (~Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.rgb_mat_rows_out_blk_n) | (~Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.rgb_mat_cols_out_blk_n) | (~Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.resize_out_mat_rows_out_blk_n) | (~Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.resize_out_mat_cols_out_blk_n);
    assign proc_1_data_PIPO_blk[2] = 1'b0;
    assign proc_1_start_FIFO_blk[2] = 1'b0 | (~start_for_resize_1_9_2160_3840_720_720_1_9_U0_U.if_full_n & Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.ap_start & ~Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.real_start & (trans_in_cnt_8 == trans_out_cnt_8) & ~start_for_resize_1_9_2160_3840_720_720_1_9_U0_U.if_read);
    assign proc_1_TLF_FIFO_blk[2] = 1'b0;
    assign proc_1_input_sync_blk[2] = 1'b0;
    assign proc_1_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_1[2] = dl_detect_out ? proc_dep_vld_vec_1_reg[2] : (proc_1_data_FIFO_blk[2] | proc_1_data_PIPO_blk[2] | proc_1_start_FIFO_blk[2] | proc_1_TLF_FIFO_blk[2] | proc_1_input_sync_blk[2] | proc_1_output_sync_blk[2]);
    assign proc_1_data_FIFO_blk[3] = 1'b0 | (~Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.out_mat_rows_out_blk_n) | (~Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit20_proc_U0.out_mat_cols_out_blk_n);
    assign proc_1_data_PIPO_blk[3] = 1'b0;
    assign proc_1_start_FIFO_blk[3] = 1'b0;
    assign proc_1_TLF_FIFO_blk[3] = 1'b0;
    assign proc_1_input_sync_blk[3] = 1'b0;
    assign proc_1_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_1[3] = dl_detect_out ? proc_dep_vld_vec_1_reg[3] : (proc_1_data_FIFO_blk[3] | proc_1_data_PIPO_blk[3] | proc_1_start_FIFO_blk[3] | proc_1_TLF_FIFO_blk[3] | proc_1_input_sync_blk[3] | proc_1_output_sync_blk[3]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_1_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_1_reg <= proc_dep_vld_vec_1;
        end
    end
    assign in_chan_dep_vld_vec_1[0] = dep_chan_vld_0_1;
    assign in_chan_dep_data_vec_1[32 : 0] = dep_chan_data_0_1;
    assign token_in_vec_1[0] = token_0_1;
    assign in_chan_dep_vld_vec_1[1] = dep_chan_vld_2_1;
    assign in_chan_dep_data_vec_1[65 : 33] = dep_chan_data_2_1;
    assign token_in_vec_1[1] = token_2_1;
    assign in_chan_dep_vld_vec_1[2] = dep_chan_vld_12_1;
    assign in_chan_dep_data_vec_1[98 : 66] = dep_chan_data_12_1;
    assign token_in_vec_1[2] = token_12_1;
    assign in_chan_dep_vld_vec_1[3] = dep_chan_vld_22_1;
    assign in_chan_dep_data_vec_1[131 : 99] = dep_chan_data_22_1;
    assign token_in_vec_1[3] = token_22_1;
    assign in_chan_dep_vld_vec_1[4] = dep_chan_vld_24_1;
    assign in_chan_dep_data_vec_1[164 : 132] = dep_chan_data_24_1;
    assign token_in_vec_1[4] = token_24_1;
    assign dep_chan_vld_1_0 = out_chan_dep_vld_vec_1[0];
    assign dep_chan_data_1_0 = out_chan_dep_data_1;
    assign token_1_0 = token_out_vec_1[0];
    assign dep_chan_vld_1_2 = out_chan_dep_vld_vec_1[1];
    assign dep_chan_data_1_2 = out_chan_dep_data_1;
    assign token_1_2 = token_out_vec_1[1];
    assign dep_chan_vld_1_22 = out_chan_dep_vld_vec_1[2];
    assign dep_chan_data_1_22 = out_chan_dep_data_1;
    assign token_1_22 = token_out_vec_1[2];
    assign dep_chan_vld_1_24 = out_chan_dep_vld_vec_1[3];
    assign dep_chan_data_1_24 = out_chan_dep_data_1;
    assign token_1_24 = token_out_vec_1[3];

    // Process: Array2xfMat_64_0_2160_3840_1_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 2, 5, 5) pp_pipeline_accel_hls_deadlock_detect_unit_2 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_2),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_2),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_2),
        .token_in_vec(token_in_vec_2),
        .dl_detect_in(dl_detect_out),
        .origin(origin[2]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_2),
        .out_chan_dep_data(out_chan_dep_data_2),
        .token_out_vec(token_out_vec_2),
        .dl_detect_out(dl_in_vec[2]));

    assign proc_2_data_FIFO_blk[0] = 1'b0 | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.AxiStream2MatStream_1_U0.imgInput_y_466_blk_n) | (~Array2xfMat_64_0_2160_3840_1_U0.dstMat_1_out_blk_n) | (~Array2xfMat_64_0_2160_3840_1_U0.dstMat_2_out_blk_n);
    assign proc_2_data_PIPO_blk[0] = 1'b0;
    assign proc_2_start_FIFO_blk[0] = 1'b0 | (~start_for_nv122bgr_0_6_9_2160_3840_1_1_U0_U.if_full_n & Array2xfMat_64_0_2160_3840_1_U0.ap_start & ~Array2xfMat_64_0_2160_3840_1_U0.real_start & (trans_in_cnt_7 == trans_out_cnt_7) & ~start_for_nv122bgr_0_6_9_2160_3840_1_1_U0_U.if_read);
    assign proc_2_TLF_FIFO_blk[0] = 1'b0;
    assign proc_2_input_sync_blk[0] = 1'b0;
    assign proc_2_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_2[0] = dl_detect_out ? proc_dep_vld_vec_2_reg[0] : (proc_2_data_FIFO_blk[0] | proc_2_data_PIPO_blk[0] | proc_2_start_FIFO_blk[0] | proc_2_TLF_FIFO_blk[0] | proc_2_input_sync_blk[0] | proc_2_output_sync_blk[0]);
    assign proc_2_data_FIFO_blk[1] = 1'b0 | (~Array2xfMat_64_0_2160_3840_1_U0.srcPtr_blk_n) | (~Array2xfMat_64_0_2160_3840_1_U0.stride_blk_n);
    assign proc_2_data_PIPO_blk[1] = 1'b0;
    assign proc_2_start_FIFO_blk[1] = 1'b0;
    assign proc_2_TLF_FIFO_blk[1] = 1'b0;
    assign proc_2_input_sync_blk[1] = 1'b0 | (ap_sync_Array2xfMat_64_0_2160_3840_1_U0_ap_ready & Array2xfMat_64_0_2160_3840_1_U0.ap_idle & ~ap_sync_pp_pipeline_accel_entry33_U0_ap_ready);
    assign proc_2_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_2[1] = dl_detect_out ? proc_dep_vld_vec_2_reg[1] : (proc_2_data_FIFO_blk[1] | proc_2_data_PIPO_blk[1] | proc_2_start_FIFO_blk[1] | proc_2_TLF_FIFO_blk[1] | proc_2_input_sync_blk[1] | proc_2_output_sync_blk[1]);
    assign proc_2_data_FIFO_blk[2] = 1'b0 | (~Array2xfMat_64_0_2160_3840_1_U0.dstMat_1_blk_n) | (~Array2xfMat_64_0_2160_3840_1_U0.dstMat_2_blk_n);
    assign proc_2_data_PIPO_blk[2] = 1'b0;
    assign proc_2_start_FIFO_blk[2] = 1'b0;
    assign proc_2_TLF_FIFO_blk[2] = 1'b0;
    assign proc_2_input_sync_blk[2] = 1'b0;
    assign proc_2_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_2[2] = dl_detect_out ? proc_dep_vld_vec_2_reg[2] : (proc_2_data_FIFO_blk[2] | proc_2_data_PIPO_blk[2] | proc_2_start_FIFO_blk[2] | proc_2_TLF_FIFO_blk[2] | proc_2_input_sync_blk[2] | proc_2_output_sync_blk[2]);
    assign proc_2_data_FIFO_blk[3] = 1'b0;
    assign proc_2_data_PIPO_blk[3] = 1'b0;
    assign proc_2_start_FIFO_blk[3] = 1'b0;
    assign proc_2_TLF_FIFO_blk[3] = 1'b0;
    assign proc_2_input_sync_blk[3] = 1'b0 | (ap_sync_Array2xfMat_64_0_2160_3840_1_U0_ap_ready & Array2xfMat_64_0_2160_3840_1_U0.ap_idle & ~ap_sync_Array2xfMat_64_6_1080_1920_1_U0_ap_ready);
    assign proc_2_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_2[3] = dl_detect_out ? proc_dep_vld_vec_2_reg[3] : (proc_2_data_FIFO_blk[3] | proc_2_data_PIPO_blk[3] | proc_2_start_FIFO_blk[3] | proc_2_TLF_FIFO_blk[3] | proc_2_input_sync_blk[3] | proc_2_output_sync_blk[3]);
    assign proc_2_data_FIFO_blk[4] = 1'b0;
    assign proc_2_data_PIPO_blk[4] = 1'b0;
    assign proc_2_start_FIFO_blk[4] = 1'b0;
    assign proc_2_TLF_FIFO_blk[4] = 1'b0;
    assign proc_2_input_sync_blk[4] = 1'b0 | (ap_sync_Array2xfMat_64_0_2160_3840_1_U0_ap_ready & Array2xfMat_64_0_2160_3840_1_U0.ap_idle & ~ap_sync_preProcess_9_9_720_720_1_8_8_8_4_8_8_U0_ap_ready);
    assign proc_2_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_2[4] = dl_detect_out ? proc_dep_vld_vec_2_reg[4] : (proc_2_data_FIFO_blk[4] | proc_2_data_PIPO_blk[4] | proc_2_start_FIFO_blk[4] | proc_2_TLF_FIFO_blk[4] | proc_2_input_sync_blk[4] | proc_2_output_sync_blk[4]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_2_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_2_reg <= proc_dep_vld_vec_2;
        end
    end
    assign in_chan_dep_vld_vec_2[0] = dep_chan_vld_0_2;
    assign in_chan_dep_data_vec_2[32 : 0] = dep_chan_data_0_2;
    assign token_in_vec_2[0] = token_0_2;
    assign in_chan_dep_vld_vec_2[1] = dep_chan_vld_1_2;
    assign in_chan_dep_data_vec_2[65 : 33] = dep_chan_data_1_2;
    assign token_in_vec_2[1] = token_1_2;
    assign in_chan_dep_vld_vec_2[2] = dep_chan_vld_12_2;
    assign in_chan_dep_data_vec_2[98 : 66] = dep_chan_data_12_2;
    assign token_in_vec_2[2] = token_12_2;
    assign in_chan_dep_vld_vec_2[3] = dep_chan_vld_21_2;
    assign in_chan_dep_data_vec_2[131 : 99] = dep_chan_data_21_2;
    assign token_in_vec_2[3] = token_21_2;
    assign in_chan_dep_vld_vec_2[4] = dep_chan_vld_23_2;
    assign in_chan_dep_data_vec_2[164 : 132] = dep_chan_data_23_2;
    assign token_in_vec_2[4] = token_23_2;
    assign dep_chan_vld_2_21 = out_chan_dep_vld_vec_2[0];
    assign dep_chan_data_2_21 = out_chan_dep_data_2;
    assign token_2_21 = token_out_vec_2[0];
    assign dep_chan_vld_2_0 = out_chan_dep_vld_vec_2[1];
    assign dep_chan_data_2_0 = out_chan_dep_data_2;
    assign token_2_0 = token_out_vec_2[1];
    assign dep_chan_vld_2_1 = out_chan_dep_vld_vec_2[2];
    assign dep_chan_data_2_1 = out_chan_dep_data_2;
    assign token_2_1 = token_out_vec_2[2];
    assign dep_chan_vld_2_12 = out_chan_dep_vld_vec_2[3];
    assign dep_chan_data_2_12 = out_chan_dep_data_2;
    assign token_2_12 = token_out_vec_2[3];
    assign dep_chan_vld_2_23 = out_chan_dep_vld_vec_2[4];
    assign dep_chan_data_2_23 = out_chan_dep_data_2;
    assign token_2_23 = token_out_vec_2[4];

    // Process: Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 3, 3, 3) pp_pipeline_accel_hls_deadlock_detect_unit_3 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_3),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_3),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_3),
        .token_in_vec(token_in_vec_3),
        .dl_detect_in(dl_detect_out),
        .origin(origin[3]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_3),
        .out_chan_dep_data(out_chan_dep_data_3),
        .token_out_vec(token_out_vec_3),
        .dl_detect_out(dl_in_vec[3]));

    assign proc_3_data_FIFO_blk[0] = 1'b0 | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0.din_out_blk_n) | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0.rows_out_blk_n) | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0.cols_out_blk_n) | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0.stride_out_blk_n);
    assign proc_3_data_PIPO_blk[0] = 1'b0;
    assign proc_3_start_FIFO_blk[0] = 1'b0 | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_Axi2Mat_entry12_U0_U.if_full_n & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0.ap_start & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0.real_start & (trans_in_cnt_1 == trans_out_cnt_1) & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_Axi2Mat_entry12_U0_U.if_read);
    assign proc_3_TLF_FIFO_blk[0] = 1'b0;
    assign proc_3_input_sync_blk[0] = 1'b0;
    assign proc_3_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_3[0] = dl_detect_out ? proc_dep_vld_vec_3_reg[0] : (proc_3_data_FIFO_blk[0] | proc_3_data_PIPO_blk[0] | proc_3_start_FIFO_blk[0] | proc_3_TLF_FIFO_blk[0] | proc_3_input_sync_blk[0] | proc_3_output_sync_blk[0]);
    assign proc_3_data_FIFO_blk[1] = 1'b0;
    assign proc_3_data_PIPO_blk[1] = 1'b0;
    assign proc_3_start_FIFO_blk[1] = 1'b0;
    assign proc_3_TLF_FIFO_blk[1] = 1'b0;
    assign proc_3_input_sync_blk[1] = 1'b0 | (Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ap_sync_Axi2Mat_1_entry3_U0_ap_ready & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0.ap_idle & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ap_sync_last_blk_pxl_width_1_U0_ap_ready);
    assign proc_3_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_3[1] = dl_detect_out ? proc_dep_vld_vec_3_reg[1] : (proc_3_data_FIFO_blk[1] | proc_3_data_PIPO_blk[1] | proc_3_start_FIFO_blk[1] | proc_3_TLF_FIFO_blk[1] | proc_3_input_sync_blk[1] | proc_3_output_sync_blk[1]);
    assign proc_3_data_FIFO_blk[2] = 1'b0;
    assign proc_3_data_PIPO_blk[2] = 1'b0;
    assign proc_3_start_FIFO_blk[2] = 1'b0;
    assign proc_3_TLF_FIFO_blk[2] = 1'b0;
    assign proc_3_input_sync_blk[2] = 1'b0 | (Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ap_sync_Axi2Mat_1_entry3_U0_ap_ready & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_1_entry3_U0.ap_idle & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ap_sync_Axi2AxiStream_1_U0_ap_ready);
    assign proc_3_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_3[2] = dl_detect_out ? proc_dep_vld_vec_3_reg[2] : (proc_3_data_FIFO_blk[2] | proc_3_data_PIPO_blk[2] | proc_3_start_FIFO_blk[2] | proc_3_TLF_FIFO_blk[2] | proc_3_input_sync_blk[2] | proc_3_output_sync_blk[2]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_3_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_3_reg <= proc_dep_vld_vec_3;
        end
    end
    assign in_chan_dep_vld_vec_3[0] = dep_chan_vld_4_3;
    assign in_chan_dep_data_vec_3[32 : 0] = dep_chan_data_4_3;
    assign token_in_vec_3[0] = token_4_3;
    assign in_chan_dep_vld_vec_3[1] = dep_chan_vld_5_3;
    assign in_chan_dep_data_vec_3[65 : 33] = dep_chan_data_5_3;
    assign token_in_vec_3[1] = token_5_3;
    assign in_chan_dep_vld_vec_3[2] = dep_chan_vld_9_3;
    assign in_chan_dep_data_vec_3[98 : 66] = dep_chan_data_9_3;
    assign token_in_vec_3[2] = token_9_3;
    assign dep_chan_vld_3_4 = out_chan_dep_vld_vec_3[0];
    assign dep_chan_data_3_4 = out_chan_dep_data_3;
    assign token_3_4 = token_out_vec_3[0];
    assign dep_chan_vld_3_5 = out_chan_dep_vld_vec_3[1];
    assign dep_chan_data_3_5 = out_chan_dep_data_3;
    assign token_3_5 = token_out_vec_3[1];
    assign dep_chan_vld_3_9 = out_chan_dep_vld_vec_3[2];
    assign dep_chan_data_3_9 = out_chan_dep_data_3;
    assign token_3_9 = token_out_vec_3[2];

    // Process: Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 4, 3, 3) pp_pipeline_accel_hls_deadlock_detect_unit_4 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_4),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_4),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_4),
        .token_in_vec(token_in_vec_4),
        .dl_detect_in(dl_detect_out),
        .origin(origin[4]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_4),
        .out_chan_dep_data(out_chan_dep_data_4),
        .token_out_vec(token_out_vec_4),
        .dl_detect_out(dl_in_vec[4]));

    assign proc_4_data_FIFO_blk[0] = 1'b0 | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0.din_blk_n) | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0.rows_blk_n) | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0.cols_blk_n) | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0.stride_blk_n);
    assign proc_4_data_PIPO_blk[0] = 1'b0;
    assign proc_4_start_FIFO_blk[0] = 1'b0 | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_Axi2Mat_entry12_U0_U.if_empty_n & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0.ap_idle & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_Axi2Mat_entry12_U0_U.if_write);
    assign proc_4_TLF_FIFO_blk[0] = 1'b0;
    assign proc_4_input_sync_blk[0] = 1'b0;
    assign proc_4_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_4[0] = dl_detect_out ? proc_dep_vld_vec_4_reg[0] : (proc_4_data_FIFO_blk[0] | proc_4_data_PIPO_blk[0] | proc_4_start_FIFO_blk[0] | proc_4_TLF_FIFO_blk[0] | proc_4_input_sync_blk[0] | proc_4_output_sync_blk[0]);
    assign proc_4_data_FIFO_blk[1] = 1'b0 | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0.din_out_blk_n);
    assign proc_4_data_PIPO_blk[1] = 1'b0;
    assign proc_4_start_FIFO_blk[1] = 1'b0;
    assign proc_4_TLF_FIFO_blk[1] = 1'b0;
    assign proc_4_input_sync_blk[1] = 1'b0;
    assign proc_4_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_4[1] = dl_detect_out ? proc_dep_vld_vec_4_reg[1] : (proc_4_data_FIFO_blk[1] | proc_4_data_PIPO_blk[1] | proc_4_start_FIFO_blk[1] | proc_4_TLF_FIFO_blk[1] | proc_4_input_sync_blk[1] | proc_4_output_sync_blk[1]);
    assign proc_4_data_FIFO_blk[2] = 1'b0 | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0.rows_out_blk_n) | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0.cols_out_blk_n) | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0.stride_out_blk_n);
    assign proc_4_data_PIPO_blk[2] = 1'b0;
    assign proc_4_start_FIFO_blk[2] = 1'b0 | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_Axi2Mat_Block_split46_proc_U0_U.if_full_n & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0.ap_start & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_entry12_U0.real_start & (trans_in_cnt_2 == trans_out_cnt_2) & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_Axi2Mat_Block_split46_proc_U0_U.if_read);
    assign proc_4_TLF_FIFO_blk[2] = 1'b0;
    assign proc_4_input_sync_blk[2] = 1'b0;
    assign proc_4_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_4[2] = dl_detect_out ? proc_dep_vld_vec_4_reg[2] : (proc_4_data_FIFO_blk[2] | proc_4_data_PIPO_blk[2] | proc_4_start_FIFO_blk[2] | proc_4_TLF_FIFO_blk[2] | proc_4_input_sync_blk[2] | proc_4_output_sync_blk[2]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_4_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_4_reg <= proc_dep_vld_vec_4;
        end
    end
    assign in_chan_dep_vld_vec_4[0] = dep_chan_vld_3_4;
    assign in_chan_dep_data_vec_4[32 : 0] = dep_chan_data_3_4;
    assign token_in_vec_4[0] = token_3_4;
    assign in_chan_dep_vld_vec_4[1] = dep_chan_vld_6_4;
    assign in_chan_dep_data_vec_4[65 : 33] = dep_chan_data_6_4;
    assign token_in_vec_4[1] = token_6_4;
    assign in_chan_dep_vld_vec_4[2] = dep_chan_vld_9_4;
    assign in_chan_dep_data_vec_4[98 : 66] = dep_chan_data_9_4;
    assign token_in_vec_4[2] = token_9_4;
    assign dep_chan_vld_4_3 = out_chan_dep_vld_vec_4[0];
    assign dep_chan_data_4_3 = out_chan_dep_data_4;
    assign token_4_3 = token_out_vec_4[0];
    assign dep_chan_vld_4_9 = out_chan_dep_vld_vec_4[1];
    assign dep_chan_data_4_9 = out_chan_dep_data_4;
    assign token_4_9 = token_out_vec_4[1];
    assign dep_chan_vld_4_6 = out_chan_dep_vld_vec_4[2];
    assign dep_chan_data_4_6 = out_chan_dep_data_4;
    assign token_4_6 = token_out_vec_4[2];

    // Process: Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_pxl_width_1_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 5, 3, 3) pp_pipeline_accel_hls_deadlock_detect_unit_5 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_5),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_5),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_5),
        .token_in_vec(token_in_vec_5),
        .dl_detect_in(dl_detect_out),
        .origin(origin[5]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_5),
        .out_chan_dep_data(out_chan_dep_data_5),
        .token_out_vec(token_out_vec_5),
        .dl_detect_out(dl_in_vec[5]));

    assign proc_5_data_FIFO_blk[0] = 1'b0 | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_pxl_width_1_U0.ret_out_blk_n);
    assign proc_5_data_PIPO_blk[0] = 1'b0;
    assign proc_5_start_FIFO_blk[0] = 1'b0 | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_AxiStream2MatStream_1_U0_U.if_full_n & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_pxl_width_1_U0.ap_start & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_pxl_width_1_U0.real_start & (trans_in_cnt_3 == trans_out_cnt_3) & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_AxiStream2MatStream_1_U0_U.if_read);
    assign proc_5_TLF_FIFO_blk[0] = 1'b0;
    assign proc_5_input_sync_blk[0] = 1'b0;
    assign proc_5_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_5[0] = dl_detect_out ? proc_dep_vld_vec_5_reg[0] : (proc_5_data_FIFO_blk[0] | proc_5_data_PIPO_blk[0] | proc_5_start_FIFO_blk[0] | proc_5_TLF_FIFO_blk[0] | proc_5_input_sync_blk[0] | proc_5_output_sync_blk[0]);
    assign proc_5_data_FIFO_blk[1] = 1'b0;
    assign proc_5_data_PIPO_blk[1] = 1'b0;
    assign proc_5_start_FIFO_blk[1] = 1'b0;
    assign proc_5_TLF_FIFO_blk[1] = 1'b0;
    assign proc_5_input_sync_blk[1] = 1'b0 | (Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ap_sync_last_blk_pxl_width_1_U0_ap_ready & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_pxl_width_1_U0.ap_idle & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ap_sync_Axi2Mat_1_entry3_U0_ap_ready);
    assign proc_5_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_5[1] = dl_detect_out ? proc_dep_vld_vec_5_reg[1] : (proc_5_data_FIFO_blk[1] | proc_5_data_PIPO_blk[1] | proc_5_start_FIFO_blk[1] | proc_5_TLF_FIFO_blk[1] | proc_5_input_sync_blk[1] | proc_5_output_sync_blk[1]);
    assign proc_5_data_FIFO_blk[2] = 1'b0;
    assign proc_5_data_PIPO_blk[2] = 1'b0;
    assign proc_5_start_FIFO_blk[2] = 1'b0;
    assign proc_5_TLF_FIFO_blk[2] = 1'b0;
    assign proc_5_input_sync_blk[2] = 1'b0 | (Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ap_sync_last_blk_pxl_width_1_U0_ap_ready & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.last_blk_pxl_width_1_U0.ap_idle & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ap_sync_Axi2AxiStream_1_U0_ap_ready);
    assign proc_5_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_5[2] = dl_detect_out ? proc_dep_vld_vec_5_reg[2] : (proc_5_data_FIFO_blk[2] | proc_5_data_PIPO_blk[2] | proc_5_start_FIFO_blk[2] | proc_5_TLF_FIFO_blk[2] | proc_5_input_sync_blk[2] | proc_5_output_sync_blk[2]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_5_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_5_reg <= proc_dep_vld_vec_5;
        end
    end
    assign in_chan_dep_vld_vec_5[0] = dep_chan_vld_3_5;
    assign in_chan_dep_data_vec_5[32 : 0] = dep_chan_data_3_5;
    assign token_in_vec_5[0] = token_3_5;
    assign in_chan_dep_vld_vec_5[1] = dep_chan_vld_9_5;
    assign in_chan_dep_data_vec_5[65 : 33] = dep_chan_data_9_5;
    assign token_in_vec_5[1] = token_9_5;
    assign in_chan_dep_vld_vec_5[2] = dep_chan_vld_10_5;
    assign in_chan_dep_data_vec_5[98 : 66] = dep_chan_data_10_5;
    assign token_in_vec_5[2] = token_10_5;
    assign dep_chan_vld_5_10 = out_chan_dep_vld_vec_5[0];
    assign dep_chan_data_5_10 = out_chan_dep_data_5;
    assign token_5_10 = token_out_vec_5[0];
    assign dep_chan_vld_5_3 = out_chan_dep_vld_vec_5[1];
    assign dep_chan_data_5_3 = out_chan_dep_data_5;
    assign token_5_3 = token_out_vec_5[1];
    assign dep_chan_vld_5_9 = out_chan_dep_vld_vec_5[2];
    assign dep_chan_data_5_9 = out_chan_dep_data_5;
    assign token_5_9 = token_out_vec_5[2];

    // Process: Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 6, 3, 2) pp_pipeline_accel_hls_deadlock_detect_unit_6 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_6),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_6),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_6),
        .token_in_vec(token_in_vec_6),
        .dl_detect_in(dl_detect_out),
        .origin(origin[6]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_6),
        .out_chan_dep_data(out_chan_dep_data_6),
        .token_out_vec(token_out_vec_6),
        .dl_detect_out(dl_in_vec[6]));

    assign proc_6_data_FIFO_blk[0] = 1'b0 | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0.stride_blk_n) | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0.cols_blk_n) | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0.rows_blk_n);
    assign proc_6_data_PIPO_blk[0] = 1'b0;
    assign proc_6_start_FIFO_blk[0] = 1'b0 | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_Axi2Mat_Block_split46_proc_U0_U.if_empty_n & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0.ap_idle & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_Axi2Mat_Block_split46_proc_U0_U.if_write);
    assign proc_6_TLF_FIFO_blk[0] = 1'b0;
    assign proc_6_input_sync_blk[0] = 1'b0;
    assign proc_6_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_6[0] = dl_detect_out ? proc_dep_vld_vec_6_reg[0] : (proc_6_data_FIFO_blk[0] | proc_6_data_PIPO_blk[0] | proc_6_start_FIFO_blk[0] | proc_6_TLF_FIFO_blk[0] | proc_6_input_sync_blk[0] | proc_6_output_sync_blk[0]);
    assign proc_6_data_FIFO_blk[1] = 1'b0 | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0.stride_out_blk_n) | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0.cols_out_blk_n) | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split46_proc_U0.rows_out_blk_n);
    assign proc_6_data_PIPO_blk[1] = 1'b0;
    assign proc_6_start_FIFO_blk[1] = 1'b0;
    assign proc_6_TLF_FIFO_blk[1] = 1'b0;
    assign proc_6_input_sync_blk[1] = 1'b0;
    assign proc_6_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_6[1] = dl_detect_out ? proc_dep_vld_vec_6_reg[1] : (proc_6_data_FIFO_blk[1] | proc_6_data_PIPO_blk[1] | proc_6_start_FIFO_blk[1] | proc_6_TLF_FIFO_blk[1] | proc_6_input_sync_blk[1] | proc_6_output_sync_blk[1]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_6_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_6_reg <= proc_dep_vld_vec_6;
        end
    end
    assign in_chan_dep_vld_vec_6[0] = dep_chan_vld_4_6;
    assign in_chan_dep_data_vec_6[32 : 0] = dep_chan_data_4_6;
    assign token_in_vec_6[0] = token_4_6;
    assign in_chan_dep_vld_vec_6[1] = dep_chan_vld_7_6;
    assign in_chan_dep_data_vec_6[65 : 33] = dep_chan_data_7_6;
    assign token_in_vec_6[1] = token_7_6;
    assign in_chan_dep_vld_vec_6[2] = dep_chan_vld_10_6;
    assign in_chan_dep_data_vec_6[98 : 66] = dep_chan_data_10_6;
    assign token_in_vec_6[2] = token_10_6;
    assign dep_chan_vld_6_4 = out_chan_dep_vld_vec_6[0];
    assign dep_chan_data_6_4 = out_chan_dep_data_6;
    assign token_6_4 = token_out_vec_6[0];
    assign dep_chan_vld_6_10 = out_chan_dep_vld_vec_6[1];
    assign dep_chan_data_6_10 = out_chan_dep_data_6;
    assign token_6_10 = token_out_vec_6[1];

    // Process: Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.addrbound_2_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 7, 1, 1) pp_pipeline_accel_hls_deadlock_detect_unit_7 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_7),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_7),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_7),
        .token_in_vec(token_in_vec_7),
        .dl_detect_in(dl_detect_out),
        .origin(origin[7]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_7),
        .out_chan_dep_data(out_chan_dep_data_7),
        .token_out_vec(token_out_vec_7),
        .dl_detect_out(dl_in_vec[7]));

    assign proc_7_data_FIFO_blk[0] = 1'b0;
    assign proc_7_data_PIPO_blk[0] = 1'b0;
    assign proc_7_start_FIFO_blk[0] = 1'b0;
    assign proc_7_TLF_FIFO_blk[0] = 1'b0 | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_cast_loc_channel_U.if_empty_n & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.addrbound_2_U0.ap_idle & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.rows_cast_loc_channel_U.if_write) | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_tmp_loc_channel_U.if_empty_n & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.addrbound_2_U0.ap_idle & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.cols_tmp_loc_channel_U.if_write);
    assign proc_7_input_sync_blk[0] = 1'b0;
    assign proc_7_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_7[0] = dl_detect_out ? proc_dep_vld_vec_7_reg[0] : (proc_7_data_FIFO_blk[0] | proc_7_data_PIPO_blk[0] | proc_7_start_FIFO_blk[0] | proc_7_TLF_FIFO_blk[0] | proc_7_input_sync_blk[0] | proc_7_output_sync_blk[0]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_7_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_7_reg <= proc_dep_vld_vec_7;
        end
    end
    assign in_chan_dep_vld_vec_7[0] = dep_chan_vld_8_7;
    assign in_chan_dep_data_vec_7[32 : 0] = dep_chan_data_8_7;
    assign token_in_vec_7[0] = token_8_7;
    assign dep_chan_vld_7_6 = out_chan_dep_vld_vec_7[0];
    assign dep_chan_data_7_6 = out_chan_dep_data_7;
    assign token_7_6 = token_out_vec_7[0];

    // Process: Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split48_proc_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 8, 1, 1) pp_pipeline_accel_hls_deadlock_detect_unit_8 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_8),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_8),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_8),
        .token_in_vec(token_in_vec_8),
        .dl_detect_in(dl_detect_out),
        .origin(origin[8]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_8),
        .out_chan_dep_data(out_chan_dep_data_8),
        .token_out_vec(token_out_vec_8),
        .dl_detect_out(dl_in_vec[8]));

    assign proc_8_data_FIFO_blk[0] = 1'b0;
    assign proc_8_data_PIPO_blk[0] = 1'b0;
    assign proc_8_start_FIFO_blk[0] = 1'b0;
    assign proc_8_TLF_FIFO_blk[0] = 1'b0 | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.p_channel_U.if_empty_n & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2Mat_Block_split48_proc_U0.ap_idle & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.p_channel_U.if_write);
    assign proc_8_input_sync_blk[0] = 1'b0;
    assign proc_8_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_8[0] = dl_detect_out ? proc_dep_vld_vec_8_reg[0] : (proc_8_data_FIFO_blk[0] | proc_8_data_PIPO_blk[0] | proc_8_start_FIFO_blk[0] | proc_8_TLF_FIFO_blk[0] | proc_8_input_sync_blk[0] | proc_8_output_sync_blk[0]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_8_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_8_reg <= proc_dep_vld_vec_8;
        end
    end
    assign in_chan_dep_vld_vec_8[0] = dep_chan_vld_9_8;
    assign in_chan_dep_data_vec_8[32 : 0] = dep_chan_data_9_8;
    assign token_in_vec_8[0] = token_9_8;
    assign dep_chan_vld_8_7 = out_chan_dep_vld_vec_8[0];
    assign dep_chan_data_8_7 = out_chan_dep_data_8;
    assign token_8_7 = token_out_vec_8[0];

    // Process: Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2AxiStream_1_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 9, 4, 5) pp_pipeline_accel_hls_deadlock_detect_unit_9 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_9),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_9),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_9),
        .token_in_vec(token_in_vec_9),
        .dl_detect_in(dl_detect_out),
        .origin(origin[9]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_9),
        .out_chan_dep_data(out_chan_dep_data_9),
        .token_out_vec(token_out_vec_9),
        .dl_detect_out(dl_in_vec[9]));

    assign proc_9_data_FIFO_blk[0] = 1'b0 | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2AxiStream_1_U0.ldata1_blk_n);
    assign proc_9_data_PIPO_blk[0] = 1'b0;
    assign proc_9_start_FIFO_blk[0] = 1'b0;
    assign proc_9_TLF_FIFO_blk[0] = 1'b0;
    assign proc_9_input_sync_blk[0] = 1'b0;
    assign proc_9_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_9[0] = dl_detect_out ? proc_dep_vld_vec_9_reg[0] : (proc_9_data_FIFO_blk[0] | proc_9_data_PIPO_blk[0] | proc_9_start_FIFO_blk[0] | proc_9_TLF_FIFO_blk[0] | proc_9_input_sync_blk[0] | proc_9_output_sync_blk[0]);
    assign proc_9_data_FIFO_blk[1] = 1'b0 | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2AxiStream_1_U0.din_blk_n);
    assign proc_9_data_PIPO_blk[1] = 1'b0;
    assign proc_9_start_FIFO_blk[1] = 1'b0;
    assign proc_9_TLF_FIFO_blk[1] = 1'b0;
    assign proc_9_input_sync_blk[1] = 1'b0;
    assign proc_9_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_9[1] = dl_detect_out ? proc_dep_vld_vec_9_reg[1] : (proc_9_data_FIFO_blk[1] | proc_9_data_PIPO_blk[1] | proc_9_start_FIFO_blk[1] | proc_9_TLF_FIFO_blk[1] | proc_9_input_sync_blk[1] | proc_9_output_sync_blk[1]);
    assign proc_9_data_FIFO_blk[2] = 1'b0;
    assign proc_9_data_PIPO_blk[2] = 1'b0;
    assign proc_9_start_FIFO_blk[2] = 1'b0;
    assign proc_9_TLF_FIFO_blk[2] = 1'b0 | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.axibound_V_U.if_empty_n & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2AxiStream_1_U0.ap_idle & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.axibound_V_U.if_write);
    assign proc_9_input_sync_blk[2] = 1'b0;
    assign proc_9_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_9[2] = dl_detect_out ? proc_dep_vld_vec_9_reg[2] : (proc_9_data_FIFO_blk[2] | proc_9_data_PIPO_blk[2] | proc_9_start_FIFO_blk[2] | proc_9_TLF_FIFO_blk[2] | proc_9_input_sync_blk[2] | proc_9_output_sync_blk[2]);
    assign proc_9_data_FIFO_blk[3] = 1'b0;
    assign proc_9_data_PIPO_blk[3] = 1'b0;
    assign proc_9_start_FIFO_blk[3] = 1'b0;
    assign proc_9_TLF_FIFO_blk[3] = 1'b0;
    assign proc_9_input_sync_blk[3] = 1'b0 | (Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ap_sync_Axi2AxiStream_1_U0_ap_ready & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2AxiStream_1_U0.ap_idle & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ap_sync_Axi2Mat_1_entry3_U0_ap_ready);
    assign proc_9_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_9[3] = dl_detect_out ? proc_dep_vld_vec_9_reg[3] : (proc_9_data_FIFO_blk[3] | proc_9_data_PIPO_blk[3] | proc_9_start_FIFO_blk[3] | proc_9_TLF_FIFO_blk[3] | proc_9_input_sync_blk[3] | proc_9_output_sync_blk[3]);
    assign proc_9_data_FIFO_blk[4] = 1'b0;
    assign proc_9_data_PIPO_blk[4] = 1'b0;
    assign proc_9_start_FIFO_blk[4] = 1'b0;
    assign proc_9_TLF_FIFO_blk[4] = 1'b0;
    assign proc_9_input_sync_blk[4] = 1'b0 | (Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ap_sync_Axi2AxiStream_1_U0_ap_ready & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.Axi2AxiStream_1_U0.ap_idle & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.ap_sync_last_blk_pxl_width_1_U0_ap_ready);
    assign proc_9_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_9[4] = dl_detect_out ? proc_dep_vld_vec_9_reg[4] : (proc_9_data_FIFO_blk[4] | proc_9_data_PIPO_blk[4] | proc_9_start_FIFO_blk[4] | proc_9_TLF_FIFO_blk[4] | proc_9_input_sync_blk[4] | proc_9_output_sync_blk[4]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_9_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_9_reg <= proc_dep_vld_vec_9;
        end
    end
    assign in_chan_dep_vld_vec_9[0] = dep_chan_vld_3_9;
    assign in_chan_dep_data_vec_9[32 : 0] = dep_chan_data_3_9;
    assign token_in_vec_9[0] = token_3_9;
    assign in_chan_dep_vld_vec_9[1] = dep_chan_vld_4_9;
    assign in_chan_dep_data_vec_9[65 : 33] = dep_chan_data_4_9;
    assign token_in_vec_9[1] = token_4_9;
    assign in_chan_dep_vld_vec_9[2] = dep_chan_vld_5_9;
    assign in_chan_dep_data_vec_9[98 : 66] = dep_chan_data_5_9;
    assign token_in_vec_9[2] = token_5_9;
    assign in_chan_dep_vld_vec_9[3] = dep_chan_vld_10_9;
    assign in_chan_dep_data_vec_9[131 : 99] = dep_chan_data_10_9;
    assign token_in_vec_9[3] = token_10_9;
    assign dep_chan_vld_9_10 = out_chan_dep_vld_vec_9[0];
    assign dep_chan_data_9_10 = out_chan_dep_data_9;
    assign token_9_10 = token_out_vec_9[0];
    assign dep_chan_vld_9_4 = out_chan_dep_vld_vec_9[1];
    assign dep_chan_data_9_4 = out_chan_dep_data_9;
    assign token_9_4 = token_out_vec_9[1];
    assign dep_chan_vld_9_8 = out_chan_dep_vld_vec_9[2];
    assign dep_chan_data_9_8 = out_chan_dep_data_9;
    assign token_9_8 = token_out_vec_9[2];
    assign dep_chan_vld_9_3 = out_chan_dep_vld_vec_9[3];
    assign dep_chan_data_9_3 = out_chan_dep_data_9;
    assign token_9_3 = token_out_vec_9[3];
    assign dep_chan_vld_9_5 = out_chan_dep_vld_vec_9[4];
    assign dep_chan_data_9_5 = out_chan_dep_data_9;
    assign token_9_5 = token_out_vec_9[4];

    // Process: Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.AxiStream2MatStream_1_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 10, 3, 3) pp_pipeline_accel_hls_deadlock_detect_unit_10 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_10),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_10),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_10),
        .token_in_vec(token_in_vec_10),
        .dl_detect_in(dl_detect_out),
        .origin(origin[10]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_10),
        .out_chan_dep_data(out_chan_dep_data_10),
        .token_out_vec(token_out_vec_10),
        .dl_detect_out(dl_in_vec[10]));

    assign proc_10_data_FIFO_blk[0] = 1'b0 | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.AxiStream2MatStream_1_U0.ldata1_blk_n);
    assign proc_10_data_PIPO_blk[0] = 1'b0;
    assign proc_10_start_FIFO_blk[0] = 1'b0;
    assign proc_10_TLF_FIFO_blk[0] = 1'b0;
    assign proc_10_input_sync_blk[0] = 1'b0;
    assign proc_10_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_10[0] = dl_detect_out ? proc_dep_vld_vec_10_reg[0] : (proc_10_data_FIFO_blk[0] | proc_10_data_PIPO_blk[0] | proc_10_start_FIFO_blk[0] | proc_10_TLF_FIFO_blk[0] | proc_10_input_sync_blk[0] | proc_10_output_sync_blk[0]);
    assign proc_10_data_FIFO_blk[1] = 1'b0 | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.AxiStream2MatStream_1_U0.rows_blk_n) | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.AxiStream2MatStream_1_U0.cols_bound_per_npc_blk_n) | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.AxiStream2MatStream_1_U0.stride_blk_n);
    assign proc_10_data_PIPO_blk[1] = 1'b0;
    assign proc_10_start_FIFO_blk[1] = 1'b0;
    assign proc_10_TLF_FIFO_blk[1] = 1'b0;
    assign proc_10_input_sync_blk[1] = 1'b0;
    assign proc_10_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_10[1] = dl_detect_out ? proc_dep_vld_vec_10_reg[1] : (proc_10_data_FIFO_blk[1] | proc_10_data_PIPO_blk[1] | proc_10_start_FIFO_blk[1] | proc_10_TLF_FIFO_blk[1] | proc_10_input_sync_blk[1] | proc_10_output_sync_blk[1]);
    assign proc_10_data_FIFO_blk[2] = 1'b0 | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.AxiStream2MatStream_1_U0.last_blk_width_blk_n);
    assign proc_10_data_PIPO_blk[2] = 1'b0;
    assign proc_10_start_FIFO_blk[2] = 1'b0 | (~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_AxiStream2MatStream_1_U0_U.if_empty_n & Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.AxiStream2MatStream_1_U0.ap_idle & ~Array2xfMat_64_0_2160_3840_1_U0.grp_Axi2Mat_1_fu_90.start_for_AxiStream2MatStream_1_U0_U.if_write);
    assign proc_10_TLF_FIFO_blk[2] = 1'b0;
    assign proc_10_input_sync_blk[2] = 1'b0;
    assign proc_10_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_10[2] = dl_detect_out ? proc_dep_vld_vec_10_reg[2] : (proc_10_data_FIFO_blk[2] | proc_10_data_PIPO_blk[2] | proc_10_start_FIFO_blk[2] | proc_10_TLF_FIFO_blk[2] | proc_10_input_sync_blk[2] | proc_10_output_sync_blk[2]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_10_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_10_reg <= proc_dep_vld_vec_10;
        end
    end
    assign in_chan_dep_vld_vec_10[0] = dep_chan_vld_5_10;
    assign in_chan_dep_data_vec_10[32 : 0] = dep_chan_data_5_10;
    assign token_in_vec_10[0] = token_5_10;
    assign in_chan_dep_vld_vec_10[1] = dep_chan_vld_6_10;
    assign in_chan_dep_data_vec_10[65 : 33] = dep_chan_data_6_10;
    assign token_in_vec_10[1] = token_6_10;
    assign in_chan_dep_vld_vec_10[2] = dep_chan_vld_9_10;
    assign in_chan_dep_data_vec_10[98 : 66] = dep_chan_data_9_10;
    assign token_in_vec_10[2] = token_9_10;
    assign dep_chan_vld_10_9 = out_chan_dep_vld_vec_10[0];
    assign dep_chan_data_10_9 = out_chan_dep_data_10;
    assign token_10_9 = token_out_vec_10[0];
    assign dep_chan_vld_10_6 = out_chan_dep_vld_vec_10[1];
    assign dep_chan_data_10_6 = out_chan_dep_data_10;
    assign token_10_6 = token_out_vec_10[1];
    assign dep_chan_vld_10_5 = out_chan_dep_vld_vec_10[2];
    assign dep_chan_data_10_5 = out_chan_dep_data_10;
    assign token_10_5 = token_out_vec_10[2];

    // Process: Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit2022_proc_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 11, 2, 1) pp_pipeline_accel_hls_deadlock_detect_unit_11 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_11),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_11),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_11),
        .token_in_vec(token_in_vec_11),
        .dl_detect_in(dl_detect_out),
        .origin(origin[11]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_11),
        .out_chan_dep_data(out_chan_dep_data_11),
        .token_out_vec(token_out_vec_11),
        .dl_detect_out(dl_in_vec[11]));

    assign proc_11_data_FIFO_blk[0] = 1'b0 | (~Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit2022_proc_U0.in_img_linestride_blk_n);
    assign proc_11_data_PIPO_blk[0] = 1'b0;
    assign proc_11_start_FIFO_blk[0] = 1'b0 | (~start_for_Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit2022_proc_U0_U.if_empty_n & Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit2022_proc_U0.ap_idle & ~start_for_Block_ZN2xf2cv3MatILi0ELi2160ELi3840ELi1ELi2EEC2Eii_exit2022_proc_U0_U.if_write);
    assign proc_11_TLF_FIFO_blk[0] = 1'b0;
    assign proc_11_input_sync_blk[0] = 1'b0;
    assign proc_11_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_11[0] = dl_detect_out ? proc_dep_vld_vec_11_reg[0] : (proc_11_data_FIFO_blk[0] | proc_11_data_PIPO_blk[0] | proc_11_start_FIFO_blk[0] | proc_11_TLF_FIFO_blk[0] | proc_11_input_sync_blk[0] | proc_11_output_sync_blk[0]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_11_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_11_reg <= proc_dep_vld_vec_11;
        end
    end
    assign in_chan_dep_vld_vec_11[0] = dep_chan_vld_0_11;
    assign in_chan_dep_data_vec_11[32 : 0] = dep_chan_data_0_11;
    assign token_in_vec_11[0] = token_0_11;
    assign in_chan_dep_vld_vec_11[1] = dep_chan_vld_12_11;
    assign in_chan_dep_data_vec_11[65 : 33] = dep_chan_data_12_11;
    assign token_in_vec_11[1] = token_12_11;
    assign dep_chan_vld_11_0 = out_chan_dep_vld_vec_11[0];
    assign dep_chan_data_11_0 = out_chan_dep_data_11;
    assign token_11_0 = token_out_vec_11[0];

    // Process: Array2xfMat_64_6_1080_1920_1_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 12, 4, 6) pp_pipeline_accel_hls_deadlock_detect_unit_12 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_12),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_12),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_12),
        .token_in_vec(token_in_vec_12),
        .dl_detect_in(dl_detect_out),
        .origin(origin[12]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_12),
        .out_chan_dep_data(out_chan_dep_data_12),
        .token_out_vec(token_out_vec_12),
        .dl_detect_out(dl_in_vec[12]));

    assign proc_12_data_FIFO_blk[0] = 1'b0 | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.AxiStream2MatStream_U0.imgInput_uv_467_blk_n);
    assign proc_12_data_PIPO_blk[0] = 1'b0;
    assign proc_12_start_FIFO_blk[0] = 1'b0;
    assign proc_12_TLF_FIFO_blk[0] = 1'b0;
    assign proc_12_input_sync_blk[0] = 1'b0;
    assign proc_12_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_12[0] = dl_detect_out ? proc_dep_vld_vec_12_reg[0] : (proc_12_data_FIFO_blk[0] | proc_12_data_PIPO_blk[0] | proc_12_start_FIFO_blk[0] | proc_12_TLF_FIFO_blk[0] | proc_12_input_sync_blk[0] | proc_12_output_sync_blk[0]);
    assign proc_12_data_FIFO_blk[1] = 1'b0 | (~Array2xfMat_64_6_1080_1920_1_U0.img_inp_uv_blk_n);
    assign proc_12_data_PIPO_blk[1] = 1'b0;
    assign proc_12_start_FIFO_blk[1] = 1'b0;
    assign proc_12_TLF_FIFO_blk[1] = 1'b0;
    assign proc_12_input_sync_blk[1] = 1'b0 | (ap_sync_Array2xfMat_64_6_1080_1920_1_U0_ap_ready & Array2xfMat_64_6_1080_1920_1_U0.ap_idle & ~ap_sync_pp_pipeline_accel_entry33_U0_ap_ready);
    assign proc_12_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_12[1] = dl_detect_out ? proc_dep_vld_vec_12_reg[1] : (proc_12_data_FIFO_blk[1] | proc_12_data_PIPO_blk[1] | proc_12_start_FIFO_blk[1] | proc_12_TLF_FIFO_blk[1] | proc_12_input_sync_blk[1] | proc_12_output_sync_blk[1]);
    assign proc_12_data_FIFO_blk[2] = 1'b0;
    assign proc_12_data_PIPO_blk[2] = 1'b0;
    assign proc_12_start_FIFO_blk[2] = 1'b0;
    assign proc_12_TLF_FIFO_blk[2] = 1'b0 | (~imgInput_uv_rows_channel_U.if_empty_n & Array2xfMat_64_6_1080_1920_1_U0.ap_idle & ~imgInput_uv_rows_channel_U.if_write) | (~imgInput_uv_cols_channel_U.if_empty_n & Array2xfMat_64_6_1080_1920_1_U0.ap_idle & ~imgInput_uv_cols_channel_U.if_write);
    assign proc_12_input_sync_blk[2] = 1'b0;
    assign proc_12_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_12[2] = dl_detect_out ? proc_dep_vld_vec_12_reg[2] : (proc_12_data_FIFO_blk[2] | proc_12_data_PIPO_blk[2] | proc_12_start_FIFO_blk[2] | proc_12_TLF_FIFO_blk[2] | proc_12_input_sync_blk[2] | proc_12_output_sync_blk[2]);
    assign proc_12_data_FIFO_blk[3] = 1'b0;
    assign proc_12_data_PIPO_blk[3] = 1'b0;
    assign proc_12_start_FIFO_blk[3] = 1'b0;
    assign proc_12_TLF_FIFO_blk[3] = 1'b0 | (~select_ln59_loc_channel_U.if_empty_n & Array2xfMat_64_6_1080_1920_1_U0.ap_idle & ~select_ln59_loc_channel_U.if_write);
    assign proc_12_input_sync_blk[3] = 1'b0;
    assign proc_12_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_12[3] = dl_detect_out ? proc_dep_vld_vec_12_reg[3] : (proc_12_data_FIFO_blk[3] | proc_12_data_PIPO_blk[3] | proc_12_start_FIFO_blk[3] | proc_12_TLF_FIFO_blk[3] | proc_12_input_sync_blk[3] | proc_12_output_sync_blk[3]);
    assign proc_12_data_FIFO_blk[4] = 1'b0;
    assign proc_12_data_PIPO_blk[4] = 1'b0;
    assign proc_12_start_FIFO_blk[4] = 1'b0;
    assign proc_12_TLF_FIFO_blk[4] = 1'b0;
    assign proc_12_input_sync_blk[4] = 1'b0 | (ap_sync_Array2xfMat_64_6_1080_1920_1_U0_ap_ready & Array2xfMat_64_6_1080_1920_1_U0.ap_idle & ~ap_sync_Array2xfMat_64_0_2160_3840_1_U0_ap_ready);
    assign proc_12_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_12[4] = dl_detect_out ? proc_dep_vld_vec_12_reg[4] : (proc_12_data_FIFO_blk[4] | proc_12_data_PIPO_blk[4] | proc_12_start_FIFO_blk[4] | proc_12_TLF_FIFO_blk[4] | proc_12_input_sync_blk[4] | proc_12_output_sync_blk[4]);
    assign proc_12_data_FIFO_blk[5] = 1'b0;
    assign proc_12_data_PIPO_blk[5] = 1'b0;
    assign proc_12_start_FIFO_blk[5] = 1'b0;
    assign proc_12_TLF_FIFO_blk[5] = 1'b0;
    assign proc_12_input_sync_blk[5] = 1'b0 | (ap_sync_Array2xfMat_64_6_1080_1920_1_U0_ap_ready & Array2xfMat_64_6_1080_1920_1_U0.ap_idle & ~ap_sync_preProcess_9_9_720_720_1_8_8_8_4_8_8_U0_ap_ready);
    assign proc_12_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_12[5] = dl_detect_out ? proc_dep_vld_vec_12_reg[5] : (proc_12_data_FIFO_blk[5] | proc_12_data_PIPO_blk[5] | proc_12_start_FIFO_blk[5] | proc_12_TLF_FIFO_blk[5] | proc_12_input_sync_blk[5] | proc_12_output_sync_blk[5]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_12_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_12_reg <= proc_dep_vld_vec_12;
        end
    end
    assign in_chan_dep_vld_vec_12[0] = dep_chan_vld_0_12;
    assign in_chan_dep_data_vec_12[32 : 0] = dep_chan_data_0_12;
    assign token_in_vec_12[0] = token_0_12;
    assign in_chan_dep_vld_vec_12[1] = dep_chan_vld_2_12;
    assign in_chan_dep_data_vec_12[65 : 33] = dep_chan_data_2_12;
    assign token_in_vec_12[1] = token_2_12;
    assign in_chan_dep_vld_vec_12[2] = dep_chan_vld_21_12;
    assign in_chan_dep_data_vec_12[98 : 66] = dep_chan_data_21_12;
    assign token_in_vec_12[2] = token_21_12;
    assign in_chan_dep_vld_vec_12[3] = dep_chan_vld_23_12;
    assign in_chan_dep_data_vec_12[131 : 99] = dep_chan_data_23_12;
    assign token_in_vec_12[3] = token_23_12;
    assign dep_chan_vld_12_21 = out_chan_dep_vld_vec_12[0];
    assign dep_chan_data_12_21 = out_chan_dep_data_12;
    assign token_12_21 = token_out_vec_12[0];
    assign dep_chan_vld_12_0 = out_chan_dep_vld_vec_12[1];
    assign dep_chan_data_12_0 = out_chan_dep_data_12;
    assign token_12_0 = token_out_vec_12[1];
    assign dep_chan_vld_12_1 = out_chan_dep_vld_vec_12[2];
    assign dep_chan_data_12_1 = out_chan_dep_data_12;
    assign token_12_1 = token_out_vec_12[2];
    assign dep_chan_vld_12_11 = out_chan_dep_vld_vec_12[3];
    assign dep_chan_data_12_11 = out_chan_dep_data_12;
    assign token_12_11 = token_out_vec_12[3];
    assign dep_chan_vld_12_2 = out_chan_dep_vld_vec_12[4];
    assign dep_chan_data_12_2 = out_chan_dep_data_12;
    assign token_12_2 = token_out_vec_12[4];
    assign dep_chan_vld_12_23 = out_chan_dep_vld_vec_12[5];
    assign dep_chan_data_12_23 = out_chan_dep_data_12;
    assign token_12_23 = token_out_vec_12[5];

    // Process: Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 13, 3, 3) pp_pipeline_accel_hls_deadlock_detect_unit_13 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_13),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_13),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_13),
        .token_in_vec(token_in_vec_13),
        .dl_detect_in(dl_detect_out),
        .origin(origin[13]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_13),
        .out_chan_dep_data(out_chan_dep_data_13),
        .token_out_vec(token_out_vec_13),
        .dl_detect_out(dl_in_vec[13]));

    assign proc_13_data_FIFO_blk[0] = 1'b0 | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0.din_out_blk_n) | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0.rows_out_blk_n) | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0.cols_out_blk_n) | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0.stride_out_blk_n);
    assign proc_13_data_PIPO_blk[0] = 1'b0;
    assign proc_13_start_FIFO_blk[0] = 1'b0 | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_Axi2Mat_entry18_U0_U.if_full_n & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0.ap_start & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0.real_start & (trans_in_cnt_4 == trans_out_cnt_4) & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_Axi2Mat_entry18_U0_U.if_read);
    assign proc_13_TLF_FIFO_blk[0] = 1'b0;
    assign proc_13_input_sync_blk[0] = 1'b0;
    assign proc_13_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_13[0] = dl_detect_out ? proc_dep_vld_vec_13_reg[0] : (proc_13_data_FIFO_blk[0] | proc_13_data_PIPO_blk[0] | proc_13_start_FIFO_blk[0] | proc_13_TLF_FIFO_blk[0] | proc_13_input_sync_blk[0] | proc_13_output_sync_blk[0]);
    assign proc_13_data_FIFO_blk[1] = 1'b0;
    assign proc_13_data_PIPO_blk[1] = 1'b0;
    assign proc_13_start_FIFO_blk[1] = 1'b0;
    assign proc_13_TLF_FIFO_blk[1] = 1'b0;
    assign proc_13_input_sync_blk[1] = 1'b0 | (Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ap_sync_Axi2Mat_entry6_U0_ap_ready & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0.ap_idle & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ap_sync_last_blk_pxl_width_U0_ap_ready);
    assign proc_13_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_13[1] = dl_detect_out ? proc_dep_vld_vec_13_reg[1] : (proc_13_data_FIFO_blk[1] | proc_13_data_PIPO_blk[1] | proc_13_start_FIFO_blk[1] | proc_13_TLF_FIFO_blk[1] | proc_13_input_sync_blk[1] | proc_13_output_sync_blk[1]);
    assign proc_13_data_FIFO_blk[2] = 1'b0;
    assign proc_13_data_PIPO_blk[2] = 1'b0;
    assign proc_13_start_FIFO_blk[2] = 1'b0;
    assign proc_13_TLF_FIFO_blk[2] = 1'b0;
    assign proc_13_input_sync_blk[2] = 1'b0 | (Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ap_sync_Axi2Mat_entry6_U0_ap_ready & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry6_U0.ap_idle & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ap_sync_Axi2AxiStream_U0_ap_ready);
    assign proc_13_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_13[2] = dl_detect_out ? proc_dep_vld_vec_13_reg[2] : (proc_13_data_FIFO_blk[2] | proc_13_data_PIPO_blk[2] | proc_13_start_FIFO_blk[2] | proc_13_TLF_FIFO_blk[2] | proc_13_input_sync_blk[2] | proc_13_output_sync_blk[2]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_13_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_13_reg <= proc_dep_vld_vec_13;
        end
    end
    assign in_chan_dep_vld_vec_13[0] = dep_chan_vld_14_13;
    assign in_chan_dep_data_vec_13[32 : 0] = dep_chan_data_14_13;
    assign token_in_vec_13[0] = token_14_13;
    assign in_chan_dep_vld_vec_13[1] = dep_chan_vld_15_13;
    assign in_chan_dep_data_vec_13[65 : 33] = dep_chan_data_15_13;
    assign token_in_vec_13[1] = token_15_13;
    assign in_chan_dep_vld_vec_13[2] = dep_chan_vld_19_13;
    assign in_chan_dep_data_vec_13[98 : 66] = dep_chan_data_19_13;
    assign token_in_vec_13[2] = token_19_13;
    assign dep_chan_vld_13_14 = out_chan_dep_vld_vec_13[0];
    assign dep_chan_data_13_14 = out_chan_dep_data_13;
    assign token_13_14 = token_out_vec_13[0];
    assign dep_chan_vld_13_15 = out_chan_dep_vld_vec_13[1];
    assign dep_chan_data_13_15 = out_chan_dep_data_13;
    assign token_13_15 = token_out_vec_13[1];
    assign dep_chan_vld_13_19 = out_chan_dep_vld_vec_13[2];
    assign dep_chan_data_13_19 = out_chan_dep_data_13;
    assign token_13_19 = token_out_vec_13[2];

    // Process: Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 14, 4, 4) pp_pipeline_accel_hls_deadlock_detect_unit_14 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_14),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_14),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_14),
        .token_in_vec(token_in_vec_14),
        .dl_detect_in(dl_detect_out),
        .origin(origin[14]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_14),
        .out_chan_dep_data(out_chan_dep_data_14),
        .token_out_vec(token_out_vec_14),
        .dl_detect_out(dl_in_vec[14]));

    assign proc_14_data_FIFO_blk[0] = 1'b0 | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0.din_blk_n) | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0.rows_blk_n) | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0.cols_blk_n) | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0.stride_blk_n);
    assign proc_14_data_PIPO_blk[0] = 1'b0;
    assign proc_14_start_FIFO_blk[0] = 1'b0 | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_Axi2Mat_entry18_U0_U.if_empty_n & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0.ap_idle & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_Axi2Mat_entry18_U0_U.if_write);
    assign proc_14_TLF_FIFO_blk[0] = 1'b0;
    assign proc_14_input_sync_blk[0] = 1'b0;
    assign proc_14_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_14[0] = dl_detect_out ? proc_dep_vld_vec_14_reg[0] : (proc_14_data_FIFO_blk[0] | proc_14_data_PIPO_blk[0] | proc_14_start_FIFO_blk[0] | proc_14_TLF_FIFO_blk[0] | proc_14_input_sync_blk[0] | proc_14_output_sync_blk[0]);
    assign proc_14_data_FIFO_blk[1] = 1'b0 | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0.din_out_blk_n);
    assign proc_14_data_PIPO_blk[1] = 1'b0;
    assign proc_14_start_FIFO_blk[1] = 1'b0;
    assign proc_14_TLF_FIFO_blk[1] = 1'b0;
    assign proc_14_input_sync_blk[1] = 1'b0;
    assign proc_14_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_14[1] = dl_detect_out ? proc_dep_vld_vec_14_reg[1] : (proc_14_data_FIFO_blk[1] | proc_14_data_PIPO_blk[1] | proc_14_start_FIFO_blk[1] | proc_14_TLF_FIFO_blk[1] | proc_14_input_sync_blk[1] | proc_14_output_sync_blk[1]);
    assign proc_14_data_FIFO_blk[2] = 1'b0 | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0.rows_out_blk_n);
    assign proc_14_data_PIPO_blk[2] = 1'b0;
    assign proc_14_start_FIFO_blk[2] = 1'b0;
    assign proc_14_TLF_FIFO_blk[2] = 1'b0;
    assign proc_14_input_sync_blk[2] = 1'b0;
    assign proc_14_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_14[2] = dl_detect_out ? proc_dep_vld_vec_14_reg[2] : (proc_14_data_FIFO_blk[2] | proc_14_data_PIPO_blk[2] | proc_14_start_FIFO_blk[2] | proc_14_TLF_FIFO_blk[2] | proc_14_input_sync_blk[2] | proc_14_output_sync_blk[2]);
    assign proc_14_data_FIFO_blk[3] = 1'b0 | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0.cols_out_blk_n) | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0.stride_out_blk_n);
    assign proc_14_data_PIPO_blk[3] = 1'b0;
    assign proc_14_start_FIFO_blk[3] = 1'b0 | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_Axi2Mat_Block_split35_proc_U0_U.if_full_n & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0.ap_start & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_entry18_U0.real_start & (trans_in_cnt_5 == trans_out_cnt_5) & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_Axi2Mat_Block_split35_proc_U0_U.if_read);
    assign proc_14_TLF_FIFO_blk[3] = 1'b0;
    assign proc_14_input_sync_blk[3] = 1'b0;
    assign proc_14_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_14[3] = dl_detect_out ? proc_dep_vld_vec_14_reg[3] : (proc_14_data_FIFO_blk[3] | proc_14_data_PIPO_blk[3] | proc_14_start_FIFO_blk[3] | proc_14_TLF_FIFO_blk[3] | proc_14_input_sync_blk[3] | proc_14_output_sync_blk[3]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_14_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_14_reg <= proc_dep_vld_vec_14;
        end
    end
    assign in_chan_dep_vld_vec_14[0] = dep_chan_vld_13_14;
    assign in_chan_dep_data_vec_14[32 : 0] = dep_chan_data_13_14;
    assign token_in_vec_14[0] = token_13_14;
    assign in_chan_dep_vld_vec_14[1] = dep_chan_vld_16_14;
    assign in_chan_dep_data_vec_14[65 : 33] = dep_chan_data_16_14;
    assign token_in_vec_14[1] = token_16_14;
    assign in_chan_dep_vld_vec_14[2] = dep_chan_vld_17_14;
    assign in_chan_dep_data_vec_14[98 : 66] = dep_chan_data_17_14;
    assign token_in_vec_14[2] = token_17_14;
    assign in_chan_dep_vld_vec_14[3] = dep_chan_vld_19_14;
    assign in_chan_dep_data_vec_14[131 : 99] = dep_chan_data_19_14;
    assign token_in_vec_14[3] = token_19_14;
    assign dep_chan_vld_14_13 = out_chan_dep_vld_vec_14[0];
    assign dep_chan_data_14_13 = out_chan_dep_data_14;
    assign token_14_13 = token_out_vec_14[0];
    assign dep_chan_vld_14_19 = out_chan_dep_vld_vec_14[1];
    assign dep_chan_data_14_19 = out_chan_dep_data_14;
    assign token_14_19 = token_out_vec_14[1];
    assign dep_chan_vld_14_17 = out_chan_dep_vld_vec_14[2];
    assign dep_chan_data_14_17 = out_chan_dep_data_14;
    assign token_14_17 = token_out_vec_14[2];
    assign dep_chan_vld_14_16 = out_chan_dep_vld_vec_14[3];
    assign dep_chan_data_14_16 = out_chan_dep_data_14;
    assign token_14_16 = token_out_vec_14[3];

    // Process: Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_pxl_width_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 15, 3, 3) pp_pipeline_accel_hls_deadlock_detect_unit_15 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_15),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_15),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_15),
        .token_in_vec(token_in_vec_15),
        .dl_detect_in(dl_detect_out),
        .origin(origin[15]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_15),
        .out_chan_dep_data(out_chan_dep_data_15),
        .token_out_vec(token_out_vec_15),
        .dl_detect_out(dl_in_vec[15]));

    assign proc_15_data_FIFO_blk[0] = 1'b0 | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_pxl_width_U0.ret_out_blk_n);
    assign proc_15_data_PIPO_blk[0] = 1'b0;
    assign proc_15_start_FIFO_blk[0] = 1'b0 | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_AxiStream2MatStream_U0_U.if_full_n & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_pxl_width_U0.ap_start & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_pxl_width_U0.real_start & (trans_in_cnt_6 == trans_out_cnt_6) & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_AxiStream2MatStream_U0_U.if_read);
    assign proc_15_TLF_FIFO_blk[0] = 1'b0;
    assign proc_15_input_sync_blk[0] = 1'b0;
    assign proc_15_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_15[0] = dl_detect_out ? proc_dep_vld_vec_15_reg[0] : (proc_15_data_FIFO_blk[0] | proc_15_data_PIPO_blk[0] | proc_15_start_FIFO_blk[0] | proc_15_TLF_FIFO_blk[0] | proc_15_input_sync_blk[0] | proc_15_output_sync_blk[0]);
    assign proc_15_data_FIFO_blk[1] = 1'b0;
    assign proc_15_data_PIPO_blk[1] = 1'b0;
    assign proc_15_start_FIFO_blk[1] = 1'b0;
    assign proc_15_TLF_FIFO_blk[1] = 1'b0;
    assign proc_15_input_sync_blk[1] = 1'b0 | (Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ap_sync_last_blk_pxl_width_U0_ap_ready & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_pxl_width_U0.ap_idle & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ap_sync_Axi2Mat_entry6_U0_ap_ready);
    assign proc_15_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_15[1] = dl_detect_out ? proc_dep_vld_vec_15_reg[1] : (proc_15_data_FIFO_blk[1] | proc_15_data_PIPO_blk[1] | proc_15_start_FIFO_blk[1] | proc_15_TLF_FIFO_blk[1] | proc_15_input_sync_blk[1] | proc_15_output_sync_blk[1]);
    assign proc_15_data_FIFO_blk[2] = 1'b0;
    assign proc_15_data_PIPO_blk[2] = 1'b0;
    assign proc_15_start_FIFO_blk[2] = 1'b0;
    assign proc_15_TLF_FIFO_blk[2] = 1'b0;
    assign proc_15_input_sync_blk[2] = 1'b0 | (Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ap_sync_last_blk_pxl_width_U0_ap_ready & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.last_blk_pxl_width_U0.ap_idle & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ap_sync_Axi2AxiStream_U0_ap_ready);
    assign proc_15_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_15[2] = dl_detect_out ? proc_dep_vld_vec_15_reg[2] : (proc_15_data_FIFO_blk[2] | proc_15_data_PIPO_blk[2] | proc_15_start_FIFO_blk[2] | proc_15_TLF_FIFO_blk[2] | proc_15_input_sync_blk[2] | proc_15_output_sync_blk[2]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_15_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_15_reg <= proc_dep_vld_vec_15;
        end
    end
    assign in_chan_dep_vld_vec_15[0] = dep_chan_vld_13_15;
    assign in_chan_dep_data_vec_15[32 : 0] = dep_chan_data_13_15;
    assign token_in_vec_15[0] = token_13_15;
    assign in_chan_dep_vld_vec_15[1] = dep_chan_vld_19_15;
    assign in_chan_dep_data_vec_15[65 : 33] = dep_chan_data_19_15;
    assign token_in_vec_15[1] = token_19_15;
    assign in_chan_dep_vld_vec_15[2] = dep_chan_vld_20_15;
    assign in_chan_dep_data_vec_15[98 : 66] = dep_chan_data_20_15;
    assign token_in_vec_15[2] = token_20_15;
    assign dep_chan_vld_15_20 = out_chan_dep_vld_vec_15[0];
    assign dep_chan_data_15_20 = out_chan_dep_data_15;
    assign token_15_20 = token_out_vec_15[0];
    assign dep_chan_vld_15_13 = out_chan_dep_vld_vec_15[1];
    assign dep_chan_data_15_13 = out_chan_dep_data_15;
    assign token_15_13 = token_out_vec_15[1];
    assign dep_chan_vld_15_19 = out_chan_dep_vld_vec_15[2];
    assign dep_chan_data_15_19 = out_chan_dep_data_15;
    assign token_15_19 = token_out_vec_15[2];

    // Process: Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split35_proc_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 16, 3, 2) pp_pipeline_accel_hls_deadlock_detect_unit_16 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_16),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_16),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_16),
        .token_in_vec(token_in_vec_16),
        .dl_detect_in(dl_detect_out),
        .origin(origin[16]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_16),
        .out_chan_dep_data(out_chan_dep_data_16),
        .token_out_vec(token_out_vec_16),
        .dl_detect_out(dl_in_vec[16]));

    assign proc_16_data_FIFO_blk[0] = 1'b0 | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split35_proc_U0.stride_blk_n) | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split35_proc_U0.cols_blk_n);
    assign proc_16_data_PIPO_blk[0] = 1'b0;
    assign proc_16_start_FIFO_blk[0] = 1'b0 | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_Axi2Mat_Block_split35_proc_U0_U.if_empty_n & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split35_proc_U0.ap_idle & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_Axi2Mat_Block_split35_proc_U0_U.if_write);
    assign proc_16_TLF_FIFO_blk[0] = 1'b0;
    assign proc_16_input_sync_blk[0] = 1'b0;
    assign proc_16_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_16[0] = dl_detect_out ? proc_dep_vld_vec_16_reg[0] : (proc_16_data_FIFO_blk[0] | proc_16_data_PIPO_blk[0] | proc_16_start_FIFO_blk[0] | proc_16_TLF_FIFO_blk[0] | proc_16_input_sync_blk[0] | proc_16_output_sync_blk[0]);
    assign proc_16_data_FIFO_blk[1] = 1'b0 | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split35_proc_U0.stride_out_blk_n) | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split35_proc_U0.cols_out_blk_n);
    assign proc_16_data_PIPO_blk[1] = 1'b0;
    assign proc_16_start_FIFO_blk[1] = 1'b0;
    assign proc_16_TLF_FIFO_blk[1] = 1'b0;
    assign proc_16_input_sync_blk[1] = 1'b0;
    assign proc_16_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_16[1] = dl_detect_out ? proc_dep_vld_vec_16_reg[1] : (proc_16_data_FIFO_blk[1] | proc_16_data_PIPO_blk[1] | proc_16_start_FIFO_blk[1] | proc_16_TLF_FIFO_blk[1] | proc_16_input_sync_blk[1] | proc_16_output_sync_blk[1]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_16_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_16_reg <= proc_dep_vld_vec_16;
        end
    end
    assign in_chan_dep_vld_vec_16[0] = dep_chan_vld_14_16;
    assign in_chan_dep_data_vec_16[32 : 0] = dep_chan_data_14_16;
    assign token_in_vec_16[0] = token_14_16;
    assign in_chan_dep_vld_vec_16[1] = dep_chan_vld_17_16;
    assign in_chan_dep_data_vec_16[65 : 33] = dep_chan_data_17_16;
    assign token_in_vec_16[1] = token_17_16;
    assign in_chan_dep_vld_vec_16[2] = dep_chan_vld_20_16;
    assign in_chan_dep_data_vec_16[98 : 66] = dep_chan_data_20_16;
    assign token_in_vec_16[2] = token_20_16;
    assign dep_chan_vld_16_14 = out_chan_dep_vld_vec_16[0];
    assign dep_chan_data_16_14 = out_chan_dep_data_16;
    assign token_16_14 = token_out_vec_16[0];
    assign dep_chan_vld_16_20 = out_chan_dep_vld_vec_16[1];
    assign dep_chan_data_16_20 = out_chan_dep_data_16;
    assign token_16_20 = token_out_vec_16[1];

    // Process: Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.addrbound_1_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 17, 3, 3) pp_pipeline_accel_hls_deadlock_detect_unit_17 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_17),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_17),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_17),
        .token_in_vec(token_in_vec_17),
        .dl_detect_in(dl_detect_out),
        .origin(origin[17]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_17),
        .out_chan_dep_data(out_chan_dep_data_17),
        .token_out_vec(token_out_vec_17),
        .dl_detect_out(dl_in_vec[17]));

    assign proc_17_data_FIFO_blk[0] = 1'b0 | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.addrbound_1_U0.rows_blk_n);
    assign proc_17_data_PIPO_blk[0] = 1'b0;
    assign proc_17_start_FIFO_blk[0] = 1'b0;
    assign proc_17_TLF_FIFO_blk[0] = 1'b0;
    assign proc_17_input_sync_blk[0] = 1'b0;
    assign proc_17_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_17[0] = dl_detect_out ? proc_dep_vld_vec_17_reg[0] : (proc_17_data_FIFO_blk[0] | proc_17_data_PIPO_blk[0] | proc_17_start_FIFO_blk[0] | proc_17_TLF_FIFO_blk[0] | proc_17_input_sync_blk[0] | proc_17_output_sync_blk[0]);
    assign proc_17_data_FIFO_blk[1] = 1'b0;
    assign proc_17_data_PIPO_blk[1] = 1'b0;
    assign proc_17_start_FIFO_blk[1] = 1'b0;
    assign proc_17_TLF_FIFO_blk[1] = 1'b0 | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_tmp_loc_channel_U.if_empty_n & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.addrbound_1_U0.ap_idle & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.cols_tmp_loc_channel_U.if_write);
    assign proc_17_input_sync_blk[1] = 1'b0;
    assign proc_17_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_17[1] = dl_detect_out ? proc_dep_vld_vec_17_reg[1] : (proc_17_data_FIFO_blk[1] | proc_17_data_PIPO_blk[1] | proc_17_start_FIFO_blk[1] | proc_17_TLF_FIFO_blk[1] | proc_17_input_sync_blk[1] | proc_17_output_sync_blk[1]);
    assign proc_17_data_FIFO_blk[2] = 1'b0 | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.addrbound_1_U0.rows_out_blk_n);
    assign proc_17_data_PIPO_blk[2] = 1'b0;
    assign proc_17_start_FIFO_blk[2] = 1'b0;
    assign proc_17_TLF_FIFO_blk[2] = 1'b0;
    assign proc_17_input_sync_blk[2] = 1'b0;
    assign proc_17_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_17[2] = dl_detect_out ? proc_dep_vld_vec_17_reg[2] : (proc_17_data_FIFO_blk[2] | proc_17_data_PIPO_blk[2] | proc_17_start_FIFO_blk[2] | proc_17_TLF_FIFO_blk[2] | proc_17_input_sync_blk[2] | proc_17_output_sync_blk[2]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_17_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_17_reg <= proc_dep_vld_vec_17;
        end
    end
    assign in_chan_dep_vld_vec_17[0] = dep_chan_vld_14_17;
    assign in_chan_dep_data_vec_17[32 : 0] = dep_chan_data_14_17;
    assign token_in_vec_17[0] = token_14_17;
    assign in_chan_dep_vld_vec_17[1] = dep_chan_vld_18_17;
    assign in_chan_dep_data_vec_17[65 : 33] = dep_chan_data_18_17;
    assign token_in_vec_17[1] = token_18_17;
    assign in_chan_dep_vld_vec_17[2] = dep_chan_vld_20_17;
    assign in_chan_dep_data_vec_17[98 : 66] = dep_chan_data_20_17;
    assign token_in_vec_17[2] = token_20_17;
    assign dep_chan_vld_17_14 = out_chan_dep_vld_vec_17[0];
    assign dep_chan_data_17_14 = out_chan_dep_data_17;
    assign token_17_14 = token_out_vec_17[0];
    assign dep_chan_vld_17_16 = out_chan_dep_vld_vec_17[1];
    assign dep_chan_data_17_16 = out_chan_dep_data_17;
    assign token_17_16 = token_out_vec_17[1];
    assign dep_chan_vld_17_20 = out_chan_dep_vld_vec_17[2];
    assign dep_chan_data_17_20 = out_chan_dep_data_17;
    assign token_17_20 = token_out_vec_17[2];

    // Process: Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split37_proc_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 18, 1, 1) pp_pipeline_accel_hls_deadlock_detect_unit_18 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_18),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_18),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_18),
        .token_in_vec(token_in_vec_18),
        .dl_detect_in(dl_detect_out),
        .origin(origin[18]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_18),
        .out_chan_dep_data(out_chan_dep_data_18),
        .token_out_vec(token_out_vec_18),
        .dl_detect_out(dl_in_vec[18]));

    assign proc_18_data_FIFO_blk[0] = 1'b0;
    assign proc_18_data_PIPO_blk[0] = 1'b0;
    assign proc_18_start_FIFO_blk[0] = 1'b0;
    assign proc_18_TLF_FIFO_blk[0] = 1'b0 | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.p_channel_U.if_empty_n & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2Mat_Block_split37_proc_U0.ap_idle & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.p_channel_U.if_write);
    assign proc_18_input_sync_blk[0] = 1'b0;
    assign proc_18_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_18[0] = dl_detect_out ? proc_dep_vld_vec_18_reg[0] : (proc_18_data_FIFO_blk[0] | proc_18_data_PIPO_blk[0] | proc_18_start_FIFO_blk[0] | proc_18_TLF_FIFO_blk[0] | proc_18_input_sync_blk[0] | proc_18_output_sync_blk[0]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_18_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_18_reg <= proc_dep_vld_vec_18;
        end
    end
    assign in_chan_dep_vld_vec_18[0] = dep_chan_vld_19_18;
    assign in_chan_dep_data_vec_18[32 : 0] = dep_chan_data_19_18;
    assign token_in_vec_18[0] = token_19_18;
    assign dep_chan_vld_18_17 = out_chan_dep_vld_vec_18[0];
    assign dep_chan_data_18_17 = out_chan_dep_data_18;
    assign token_18_17 = token_out_vec_18[0];

    // Process: Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2AxiStream_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 19, 4, 5) pp_pipeline_accel_hls_deadlock_detect_unit_19 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_19),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_19),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_19),
        .token_in_vec(token_in_vec_19),
        .dl_detect_in(dl_detect_out),
        .origin(origin[19]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_19),
        .out_chan_dep_data(out_chan_dep_data_19),
        .token_out_vec(token_out_vec_19),
        .dl_detect_out(dl_in_vec[19]));

    assign proc_19_data_FIFO_blk[0] = 1'b0 | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2AxiStream_U0.ldata1_blk_n);
    assign proc_19_data_PIPO_blk[0] = 1'b0;
    assign proc_19_start_FIFO_blk[0] = 1'b0;
    assign proc_19_TLF_FIFO_blk[0] = 1'b0;
    assign proc_19_input_sync_blk[0] = 1'b0;
    assign proc_19_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_19[0] = dl_detect_out ? proc_dep_vld_vec_19_reg[0] : (proc_19_data_FIFO_blk[0] | proc_19_data_PIPO_blk[0] | proc_19_start_FIFO_blk[0] | proc_19_TLF_FIFO_blk[0] | proc_19_input_sync_blk[0] | proc_19_output_sync_blk[0]);
    assign proc_19_data_FIFO_blk[1] = 1'b0 | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2AxiStream_U0.din_blk_n);
    assign proc_19_data_PIPO_blk[1] = 1'b0;
    assign proc_19_start_FIFO_blk[1] = 1'b0;
    assign proc_19_TLF_FIFO_blk[1] = 1'b0;
    assign proc_19_input_sync_blk[1] = 1'b0;
    assign proc_19_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_19[1] = dl_detect_out ? proc_dep_vld_vec_19_reg[1] : (proc_19_data_FIFO_blk[1] | proc_19_data_PIPO_blk[1] | proc_19_start_FIFO_blk[1] | proc_19_TLF_FIFO_blk[1] | proc_19_input_sync_blk[1] | proc_19_output_sync_blk[1]);
    assign proc_19_data_FIFO_blk[2] = 1'b0;
    assign proc_19_data_PIPO_blk[2] = 1'b0;
    assign proc_19_start_FIFO_blk[2] = 1'b0;
    assign proc_19_TLF_FIFO_blk[2] = 1'b0 | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.axibound_V_U.if_empty_n & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2AxiStream_U0.ap_idle & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.axibound_V_U.if_write);
    assign proc_19_input_sync_blk[2] = 1'b0;
    assign proc_19_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_19[2] = dl_detect_out ? proc_dep_vld_vec_19_reg[2] : (proc_19_data_FIFO_blk[2] | proc_19_data_PIPO_blk[2] | proc_19_start_FIFO_blk[2] | proc_19_TLF_FIFO_blk[2] | proc_19_input_sync_blk[2] | proc_19_output_sync_blk[2]);
    assign proc_19_data_FIFO_blk[3] = 1'b0;
    assign proc_19_data_PIPO_blk[3] = 1'b0;
    assign proc_19_start_FIFO_blk[3] = 1'b0;
    assign proc_19_TLF_FIFO_blk[3] = 1'b0;
    assign proc_19_input_sync_blk[3] = 1'b0 | (Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ap_sync_Axi2AxiStream_U0_ap_ready & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2AxiStream_U0.ap_idle & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ap_sync_Axi2Mat_entry6_U0_ap_ready);
    assign proc_19_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_19[3] = dl_detect_out ? proc_dep_vld_vec_19_reg[3] : (proc_19_data_FIFO_blk[3] | proc_19_data_PIPO_blk[3] | proc_19_start_FIFO_blk[3] | proc_19_TLF_FIFO_blk[3] | proc_19_input_sync_blk[3] | proc_19_output_sync_blk[3]);
    assign proc_19_data_FIFO_blk[4] = 1'b0;
    assign proc_19_data_PIPO_blk[4] = 1'b0;
    assign proc_19_start_FIFO_blk[4] = 1'b0;
    assign proc_19_TLF_FIFO_blk[4] = 1'b0;
    assign proc_19_input_sync_blk[4] = 1'b0 | (Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ap_sync_Axi2AxiStream_U0_ap_ready & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.Axi2AxiStream_U0.ap_idle & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.ap_sync_last_blk_pxl_width_U0_ap_ready);
    assign proc_19_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_19[4] = dl_detect_out ? proc_dep_vld_vec_19_reg[4] : (proc_19_data_FIFO_blk[4] | proc_19_data_PIPO_blk[4] | proc_19_start_FIFO_blk[4] | proc_19_TLF_FIFO_blk[4] | proc_19_input_sync_blk[4] | proc_19_output_sync_blk[4]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_19_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_19_reg <= proc_dep_vld_vec_19;
        end
    end
    assign in_chan_dep_vld_vec_19[0] = dep_chan_vld_13_19;
    assign in_chan_dep_data_vec_19[32 : 0] = dep_chan_data_13_19;
    assign token_in_vec_19[0] = token_13_19;
    assign in_chan_dep_vld_vec_19[1] = dep_chan_vld_14_19;
    assign in_chan_dep_data_vec_19[65 : 33] = dep_chan_data_14_19;
    assign token_in_vec_19[1] = token_14_19;
    assign in_chan_dep_vld_vec_19[2] = dep_chan_vld_15_19;
    assign in_chan_dep_data_vec_19[98 : 66] = dep_chan_data_15_19;
    assign token_in_vec_19[2] = token_15_19;
    assign in_chan_dep_vld_vec_19[3] = dep_chan_vld_20_19;
    assign in_chan_dep_data_vec_19[131 : 99] = dep_chan_data_20_19;
    assign token_in_vec_19[3] = token_20_19;
    assign dep_chan_vld_19_20 = out_chan_dep_vld_vec_19[0];
    assign dep_chan_data_19_20 = out_chan_dep_data_19;
    assign token_19_20 = token_out_vec_19[0];
    assign dep_chan_vld_19_14 = out_chan_dep_vld_vec_19[1];
    assign dep_chan_data_19_14 = out_chan_dep_data_19;
    assign token_19_14 = token_out_vec_19[1];
    assign dep_chan_vld_19_18 = out_chan_dep_vld_vec_19[2];
    assign dep_chan_data_19_18 = out_chan_dep_data_19;
    assign token_19_18 = token_out_vec_19[2];
    assign dep_chan_vld_19_13 = out_chan_dep_vld_vec_19[3];
    assign dep_chan_data_19_13 = out_chan_dep_data_19;
    assign token_19_13 = token_out_vec_19[3];
    assign dep_chan_vld_19_15 = out_chan_dep_vld_vec_19[4];
    assign dep_chan_data_19_15 = out_chan_dep_data_19;
    assign token_19_15 = token_out_vec_19[4];

    // Process: Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.AxiStream2MatStream_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 20, 4, 4) pp_pipeline_accel_hls_deadlock_detect_unit_20 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_20),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_20),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_20),
        .token_in_vec(token_in_vec_20),
        .dl_detect_in(dl_detect_out),
        .origin(origin[20]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_20),
        .out_chan_dep_data(out_chan_dep_data_20),
        .token_out_vec(token_out_vec_20),
        .dl_detect_out(dl_in_vec[20]));

    assign proc_20_data_FIFO_blk[0] = 1'b0 | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.AxiStream2MatStream_U0.ldata1_blk_n);
    assign proc_20_data_PIPO_blk[0] = 1'b0;
    assign proc_20_start_FIFO_blk[0] = 1'b0;
    assign proc_20_TLF_FIFO_blk[0] = 1'b0;
    assign proc_20_input_sync_blk[0] = 1'b0;
    assign proc_20_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_20[0] = dl_detect_out ? proc_dep_vld_vec_20_reg[0] : (proc_20_data_FIFO_blk[0] | proc_20_data_PIPO_blk[0] | proc_20_start_FIFO_blk[0] | proc_20_TLF_FIFO_blk[0] | proc_20_input_sync_blk[0] | proc_20_output_sync_blk[0]);
    assign proc_20_data_FIFO_blk[1] = 1'b0 | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.AxiStream2MatStream_U0.rows_blk_n);
    assign proc_20_data_PIPO_blk[1] = 1'b0;
    assign proc_20_start_FIFO_blk[1] = 1'b0;
    assign proc_20_TLF_FIFO_blk[1] = 1'b0;
    assign proc_20_input_sync_blk[1] = 1'b0;
    assign proc_20_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_20[1] = dl_detect_out ? proc_dep_vld_vec_20_reg[1] : (proc_20_data_FIFO_blk[1] | proc_20_data_PIPO_blk[1] | proc_20_start_FIFO_blk[1] | proc_20_TLF_FIFO_blk[1] | proc_20_input_sync_blk[1] | proc_20_output_sync_blk[1]);
    assign proc_20_data_FIFO_blk[2] = 1'b0 | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.AxiStream2MatStream_U0.cols_bound_per_npc_blk_n) | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.AxiStream2MatStream_U0.stride_blk_n);
    assign proc_20_data_PIPO_blk[2] = 1'b0;
    assign proc_20_start_FIFO_blk[2] = 1'b0;
    assign proc_20_TLF_FIFO_blk[2] = 1'b0;
    assign proc_20_input_sync_blk[2] = 1'b0;
    assign proc_20_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_20[2] = dl_detect_out ? proc_dep_vld_vec_20_reg[2] : (proc_20_data_FIFO_blk[2] | proc_20_data_PIPO_blk[2] | proc_20_start_FIFO_blk[2] | proc_20_TLF_FIFO_blk[2] | proc_20_input_sync_blk[2] | proc_20_output_sync_blk[2]);
    assign proc_20_data_FIFO_blk[3] = 1'b0 | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.AxiStream2MatStream_U0.last_blk_width_blk_n);
    assign proc_20_data_PIPO_blk[3] = 1'b0;
    assign proc_20_start_FIFO_blk[3] = 1'b0 | (~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_AxiStream2MatStream_U0_U.if_empty_n & Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.AxiStream2MatStream_U0.ap_idle & ~Array2xfMat_64_6_1080_1920_1_U0.grp_Axi2Mat_fu_70.start_for_AxiStream2MatStream_U0_U.if_write);
    assign proc_20_TLF_FIFO_blk[3] = 1'b0;
    assign proc_20_input_sync_blk[3] = 1'b0;
    assign proc_20_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_20[3] = dl_detect_out ? proc_dep_vld_vec_20_reg[3] : (proc_20_data_FIFO_blk[3] | proc_20_data_PIPO_blk[3] | proc_20_start_FIFO_blk[3] | proc_20_TLF_FIFO_blk[3] | proc_20_input_sync_blk[3] | proc_20_output_sync_blk[3]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_20_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_20_reg <= proc_dep_vld_vec_20;
        end
    end
    assign in_chan_dep_vld_vec_20[0] = dep_chan_vld_15_20;
    assign in_chan_dep_data_vec_20[32 : 0] = dep_chan_data_15_20;
    assign token_in_vec_20[0] = token_15_20;
    assign in_chan_dep_vld_vec_20[1] = dep_chan_vld_16_20;
    assign in_chan_dep_data_vec_20[65 : 33] = dep_chan_data_16_20;
    assign token_in_vec_20[1] = token_16_20;
    assign in_chan_dep_vld_vec_20[2] = dep_chan_vld_17_20;
    assign in_chan_dep_data_vec_20[98 : 66] = dep_chan_data_17_20;
    assign token_in_vec_20[2] = token_17_20;
    assign in_chan_dep_vld_vec_20[3] = dep_chan_vld_19_20;
    assign in_chan_dep_data_vec_20[131 : 99] = dep_chan_data_19_20;
    assign token_in_vec_20[3] = token_19_20;
    assign dep_chan_vld_20_19 = out_chan_dep_vld_vec_20[0];
    assign dep_chan_data_20_19 = out_chan_dep_data_20;
    assign token_20_19 = token_out_vec_20[0];
    assign dep_chan_vld_20_17 = out_chan_dep_vld_vec_20[1];
    assign dep_chan_data_20_17 = out_chan_dep_data_20;
    assign token_20_17 = token_out_vec_20[1];
    assign dep_chan_vld_20_16 = out_chan_dep_vld_vec_20[2];
    assign dep_chan_data_20_16 = out_chan_dep_data_20;
    assign token_20_16 = token_out_vec_20[2];
    assign dep_chan_vld_20_15 = out_chan_dep_vld_vec_20[3];
    assign dep_chan_data_20_15 = out_chan_dep_data_20;
    assign token_20_15 = token_out_vec_20[3];

    // Process: nv122bgr_0_6_9_2160_3840_1_1_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 21, 3, 3) pp_pipeline_accel_hls_deadlock_detect_unit_21 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_21),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_21),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_21),
        .token_in_vec(token_in_vec_21),
        .dl_detect_in(dl_detect_out),
        .origin(origin[21]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_21),
        .out_chan_dep_data(out_chan_dep_data_21),
        .token_out_vec(token_out_vec_21),
        .dl_detect_out(dl_in_vec[21]));

    assign proc_21_data_FIFO_blk[0] = 1'b0 | (~nv122bgr_0_6_9_2160_3840_1_1_U0.grp_KernNv122bgr_0_6_9_2160_3840_1_1_1_5_9_s_fu_44.imgInput_y_466_blk_n) | (~nv122bgr_0_6_9_2160_3840_1_1_U0.src_y_rows_blk_n) | (~nv122bgr_0_6_9_2160_3840_1_1_U0.src_y_cols_blk_n);
    assign proc_21_data_PIPO_blk[0] = 1'b0;
    assign proc_21_start_FIFO_blk[0] = 1'b0 | (~start_for_nv122bgr_0_6_9_2160_3840_1_1_U0_U.if_empty_n & nv122bgr_0_6_9_2160_3840_1_1_U0.ap_idle & ~start_for_nv122bgr_0_6_9_2160_3840_1_1_U0_U.if_write);
    assign proc_21_TLF_FIFO_blk[0] = 1'b0;
    assign proc_21_input_sync_blk[0] = 1'b0;
    assign proc_21_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_21[0] = dl_detect_out ? proc_dep_vld_vec_21_reg[0] : (proc_21_data_FIFO_blk[0] | proc_21_data_PIPO_blk[0] | proc_21_start_FIFO_blk[0] | proc_21_TLF_FIFO_blk[0] | proc_21_input_sync_blk[0] | proc_21_output_sync_blk[0]);
    assign proc_21_data_FIFO_blk[1] = 1'b0 | (~nv122bgr_0_6_9_2160_3840_1_1_U0.grp_KernNv122bgr_0_6_9_2160_3840_1_1_1_5_9_s_fu_44.imgInput_uv_467_blk_n);
    assign proc_21_data_PIPO_blk[1] = 1'b0;
    assign proc_21_start_FIFO_blk[1] = 1'b0;
    assign proc_21_TLF_FIFO_blk[1] = 1'b0;
    assign proc_21_input_sync_blk[1] = 1'b0;
    assign proc_21_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_21[1] = dl_detect_out ? proc_dep_vld_vec_21_reg[1] : (proc_21_data_FIFO_blk[1] | proc_21_data_PIPO_blk[1] | proc_21_start_FIFO_blk[1] | proc_21_TLF_FIFO_blk[1] | proc_21_input_sync_blk[1] | proc_21_output_sync_blk[1]);
    assign proc_21_data_FIFO_blk[2] = 1'b0 | (~nv122bgr_0_6_9_2160_3840_1_1_U0.grp_KernNv122bgr_0_6_9_2160_3840_1_1_1_5_9_s_fu_44.rgb_mat_468_blk_n);
    assign proc_21_data_PIPO_blk[2] = 1'b0;
    assign proc_21_start_FIFO_blk[2] = 1'b0;
    assign proc_21_TLF_FIFO_blk[2] = 1'b0;
    assign proc_21_input_sync_blk[2] = 1'b0;
    assign proc_21_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_21[2] = dl_detect_out ? proc_dep_vld_vec_21_reg[2] : (proc_21_data_FIFO_blk[2] | proc_21_data_PIPO_blk[2] | proc_21_start_FIFO_blk[2] | proc_21_TLF_FIFO_blk[2] | proc_21_input_sync_blk[2] | proc_21_output_sync_blk[2]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_21_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_21_reg <= proc_dep_vld_vec_21;
        end
    end
    assign in_chan_dep_vld_vec_21[0] = dep_chan_vld_2_21;
    assign in_chan_dep_data_vec_21[32 : 0] = dep_chan_data_2_21;
    assign token_in_vec_21[0] = token_2_21;
    assign in_chan_dep_vld_vec_21[1] = dep_chan_vld_12_21;
    assign in_chan_dep_data_vec_21[65 : 33] = dep_chan_data_12_21;
    assign token_in_vec_21[1] = token_12_21;
    assign in_chan_dep_vld_vec_21[2] = dep_chan_vld_22_21;
    assign in_chan_dep_data_vec_21[98 : 66] = dep_chan_data_22_21;
    assign token_in_vec_21[2] = token_22_21;
    assign dep_chan_vld_21_2 = out_chan_dep_vld_vec_21[0];
    assign dep_chan_data_21_2 = out_chan_dep_data_21;
    assign token_21_2 = token_out_vec_21[0];
    assign dep_chan_vld_21_12 = out_chan_dep_vld_vec_21[1];
    assign dep_chan_data_21_12 = out_chan_dep_data_21;
    assign token_21_12 = token_out_vec_21[1];
    assign dep_chan_vld_21_22 = out_chan_dep_vld_vec_21[2];
    assign dep_chan_data_21_22 = out_chan_dep_data_21;
    assign token_21_22 = token_out_vec_21[2];

    // Process: resize_1_9_2160_3840_720_720_1_9_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 22, 3, 3) pp_pipeline_accel_hls_deadlock_detect_unit_22 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_22),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_22),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_22),
        .token_in_vec(token_in_vec_22),
        .dl_detect_in(dl_detect_out),
        .origin(origin[22]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_22),
        .out_chan_dep_data(out_chan_dep_data_22),
        .token_out_vec(token_out_vec_22),
        .dl_detect_out(dl_in_vec[22]));

    assign proc_22_data_FIFO_blk[0] = 1'b0 | (~resize_1_9_2160_3840_720_720_1_9_U0.grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_80.rgb_mat_468_blk_n);
    assign proc_22_data_PIPO_blk[0] = 1'b0;
    assign proc_22_start_FIFO_blk[0] = 1'b0;
    assign proc_22_TLF_FIFO_blk[0] = 1'b0;
    assign proc_22_input_sync_blk[0] = 1'b0;
    assign proc_22_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_22[0] = dl_detect_out ? proc_dep_vld_vec_22_reg[0] : (proc_22_data_FIFO_blk[0] | proc_22_data_PIPO_blk[0] | proc_22_start_FIFO_blk[0] | proc_22_TLF_FIFO_blk[0] | proc_22_input_sync_blk[0] | proc_22_output_sync_blk[0]);
    assign proc_22_data_FIFO_blk[1] = 1'b0 | (~resize_1_9_2160_3840_720_720_1_9_U0.grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_80.resize_out_mat_469_blk_n) | (~resize_1_9_2160_3840_720_720_1_9_U0.p_dst_rows_out_blk_n) | (~resize_1_9_2160_3840_720_720_1_9_U0.p_dst_cols_out_blk_n);
    assign proc_22_data_PIPO_blk[1] = 1'b0;
    assign proc_22_start_FIFO_blk[1] = 1'b0;
    assign proc_22_TLF_FIFO_blk[1] = 1'b0;
    assign proc_22_input_sync_blk[1] = 1'b0;
    assign proc_22_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_22[1] = dl_detect_out ? proc_dep_vld_vec_22_reg[1] : (proc_22_data_FIFO_blk[1] | proc_22_data_PIPO_blk[1] | proc_22_start_FIFO_blk[1] | proc_22_TLF_FIFO_blk[1] | proc_22_input_sync_blk[1] | proc_22_output_sync_blk[1]);
    assign proc_22_data_FIFO_blk[2] = 1'b0 | (~resize_1_9_2160_3840_720_720_1_9_U0.p_src_rows_blk_n) | (~resize_1_9_2160_3840_720_720_1_9_U0.p_src_cols_blk_n) | (~resize_1_9_2160_3840_720_720_1_9_U0.p_dst_rows_blk_n) | (~resize_1_9_2160_3840_720_720_1_9_U0.p_dst_cols_blk_n);
    assign proc_22_data_PIPO_blk[2] = 1'b0;
    assign proc_22_start_FIFO_blk[2] = 1'b0 | (~start_for_resize_1_9_2160_3840_720_720_1_9_U0_U.if_empty_n & resize_1_9_2160_3840_720_720_1_9_U0.ap_idle & ~start_for_resize_1_9_2160_3840_720_720_1_9_U0_U.if_write);
    assign proc_22_TLF_FIFO_blk[2] = 1'b0;
    assign proc_22_input_sync_blk[2] = 1'b0;
    assign proc_22_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_22[2] = dl_detect_out ? proc_dep_vld_vec_22_reg[2] : (proc_22_data_FIFO_blk[2] | proc_22_data_PIPO_blk[2] | proc_22_start_FIFO_blk[2] | proc_22_TLF_FIFO_blk[2] | proc_22_input_sync_blk[2] | proc_22_output_sync_blk[2]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_22_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_22_reg <= proc_dep_vld_vec_22;
        end
    end
    assign in_chan_dep_vld_vec_22[0] = dep_chan_vld_1_22;
    assign in_chan_dep_data_vec_22[32 : 0] = dep_chan_data_1_22;
    assign token_in_vec_22[0] = token_1_22;
    assign in_chan_dep_vld_vec_22[1] = dep_chan_vld_21_22;
    assign in_chan_dep_data_vec_22[65 : 33] = dep_chan_data_21_22;
    assign token_in_vec_22[1] = token_21_22;
    assign in_chan_dep_vld_vec_22[2] = dep_chan_vld_23_22;
    assign in_chan_dep_data_vec_22[98 : 66] = dep_chan_data_23_22;
    assign token_in_vec_22[2] = token_23_22;
    assign dep_chan_vld_22_21 = out_chan_dep_vld_vec_22[0];
    assign dep_chan_data_22_21 = out_chan_dep_data_22;
    assign token_22_21 = token_out_vec_22[0];
    assign dep_chan_vld_22_23 = out_chan_dep_vld_vec_22[1];
    assign dep_chan_data_22_23 = out_chan_dep_data_22;
    assign token_22_23 = token_out_vec_22[1];
    assign dep_chan_vld_22_1 = out_chan_dep_vld_vec_22[2];
    assign dep_chan_data_22_1 = out_chan_dep_data_22;
    assign token_22_1 = token_out_vec_22[2];

    // Process: preProcess_9_9_720_720_1_8_8_8_4_8_8_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 23, 5, 5) pp_pipeline_accel_hls_deadlock_detect_unit_23 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_23),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_23),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_23),
        .token_in_vec(token_in_vec_23),
        .dl_detect_in(dl_detect_out),
        .origin(origin[23]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_23),
        .out_chan_dep_data(out_chan_dep_data_23),
        .token_out_vec(token_out_vec_23),
        .dl_detect_out(dl_in_vec[23]));

    assign proc_23_data_FIFO_blk[0] = 1'b0 | (~preProcess_9_9_720_720_1_8_8_8_4_8_8_U0.resize_out_mat_469_blk_n) | (~preProcess_9_9_720_720_1_8_8_8_4_8_8_U0.in_mat_rows_blk_n) | (~preProcess_9_9_720_720_1_8_8_8_4_8_8_U0.in_mat_cols_blk_n);
    assign proc_23_data_PIPO_blk[0] = 1'b0;
    assign proc_23_start_FIFO_blk[0] = 1'b0;
    assign proc_23_TLF_FIFO_blk[0] = 1'b0;
    assign proc_23_input_sync_blk[0] = 1'b0;
    assign proc_23_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_23[0] = dl_detect_out ? proc_dep_vld_vec_23_reg[0] : (proc_23_data_FIFO_blk[0] | proc_23_data_PIPO_blk[0] | proc_23_start_FIFO_blk[0] | proc_23_TLF_FIFO_blk[0] | proc_23_input_sync_blk[0] | proc_23_output_sync_blk[0]);
    assign proc_23_data_FIFO_blk[1] = 1'b0 | (~preProcess_9_9_720_720_1_8_8_8_4_8_8_U0.out_mat_470_blk_n);
    assign proc_23_data_PIPO_blk[1] = 1'b0;
    assign proc_23_start_FIFO_blk[1] = 1'b0;
    assign proc_23_TLF_FIFO_blk[1] = 1'b0;
    assign proc_23_input_sync_blk[1] = 1'b0;
    assign proc_23_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_23[1] = dl_detect_out ? proc_dep_vld_vec_23_reg[1] : (proc_23_data_FIFO_blk[1] | proc_23_data_PIPO_blk[1] | proc_23_start_FIFO_blk[1] | proc_23_TLF_FIFO_blk[1] | proc_23_input_sync_blk[1] | proc_23_output_sync_blk[1]);
    assign proc_23_data_FIFO_blk[2] = 1'b0 | (~preProcess_9_9_720_720_1_8_8_8_4_8_8_U0.params_blk_n);
    assign proc_23_data_PIPO_blk[2] = 1'b0;
    assign proc_23_start_FIFO_blk[2] = 1'b0;
    assign proc_23_TLF_FIFO_blk[2] = 1'b0;
    assign proc_23_input_sync_blk[2] = 1'b0 | (ap_sync_preProcess_9_9_720_720_1_8_8_8_4_8_8_U0_ap_ready & preProcess_9_9_720_720_1_8_8_8_4_8_8_U0.ap_idle & ~ap_sync_pp_pipeline_accel_entry33_U0_ap_ready);
    assign proc_23_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_23[2] = dl_detect_out ? proc_dep_vld_vec_23_reg[2] : (proc_23_data_FIFO_blk[2] | proc_23_data_PIPO_blk[2] | proc_23_start_FIFO_blk[2] | proc_23_TLF_FIFO_blk[2] | proc_23_input_sync_blk[2] | proc_23_output_sync_blk[2]);
    assign proc_23_data_FIFO_blk[3] = 1'b0;
    assign proc_23_data_PIPO_blk[3] = 1'b0;
    assign proc_23_start_FIFO_blk[3] = 1'b0;
    assign proc_23_TLF_FIFO_blk[3] = 1'b0;
    assign proc_23_input_sync_blk[3] = 1'b0 | (ap_sync_preProcess_9_9_720_720_1_8_8_8_4_8_8_U0_ap_ready & preProcess_9_9_720_720_1_8_8_8_4_8_8_U0.ap_idle & ~ap_sync_Array2xfMat_64_0_2160_3840_1_U0_ap_ready);
    assign proc_23_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_23[3] = dl_detect_out ? proc_dep_vld_vec_23_reg[3] : (proc_23_data_FIFO_blk[3] | proc_23_data_PIPO_blk[3] | proc_23_start_FIFO_blk[3] | proc_23_TLF_FIFO_blk[3] | proc_23_input_sync_blk[3] | proc_23_output_sync_blk[3]);
    assign proc_23_data_FIFO_blk[4] = 1'b0;
    assign proc_23_data_PIPO_blk[4] = 1'b0;
    assign proc_23_start_FIFO_blk[4] = 1'b0;
    assign proc_23_TLF_FIFO_blk[4] = 1'b0;
    assign proc_23_input_sync_blk[4] = 1'b0 | (ap_sync_preProcess_9_9_720_720_1_8_8_8_4_8_8_U0_ap_ready & preProcess_9_9_720_720_1_8_8_8_4_8_8_U0.ap_idle & ~ap_sync_Array2xfMat_64_6_1080_1920_1_U0_ap_ready);
    assign proc_23_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_23[4] = dl_detect_out ? proc_dep_vld_vec_23_reg[4] : (proc_23_data_FIFO_blk[4] | proc_23_data_PIPO_blk[4] | proc_23_start_FIFO_blk[4] | proc_23_TLF_FIFO_blk[4] | proc_23_input_sync_blk[4] | proc_23_output_sync_blk[4]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_23_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_23_reg <= proc_dep_vld_vec_23;
        end
    end
    assign in_chan_dep_vld_vec_23[0] = dep_chan_vld_0_23;
    assign in_chan_dep_data_vec_23[32 : 0] = dep_chan_data_0_23;
    assign token_in_vec_23[0] = token_0_23;
    assign in_chan_dep_vld_vec_23[1] = dep_chan_vld_2_23;
    assign in_chan_dep_data_vec_23[65 : 33] = dep_chan_data_2_23;
    assign token_in_vec_23[1] = token_2_23;
    assign in_chan_dep_vld_vec_23[2] = dep_chan_vld_12_23;
    assign in_chan_dep_data_vec_23[98 : 66] = dep_chan_data_12_23;
    assign token_in_vec_23[2] = token_12_23;
    assign in_chan_dep_vld_vec_23[3] = dep_chan_vld_22_23;
    assign in_chan_dep_data_vec_23[131 : 99] = dep_chan_data_22_23;
    assign token_in_vec_23[3] = token_22_23;
    assign in_chan_dep_vld_vec_23[4] = dep_chan_vld_24_23;
    assign in_chan_dep_data_vec_23[164 : 132] = dep_chan_data_24_23;
    assign token_in_vec_23[4] = token_24_23;
    assign dep_chan_vld_23_22 = out_chan_dep_vld_vec_23[0];
    assign dep_chan_data_23_22 = out_chan_dep_data_23;
    assign token_23_22 = token_out_vec_23[0];
    assign dep_chan_vld_23_24 = out_chan_dep_vld_vec_23[1];
    assign dep_chan_data_23_24 = out_chan_dep_data_23;
    assign token_23_24 = token_out_vec_23[1];
    assign dep_chan_vld_23_0 = out_chan_dep_vld_vec_23[2];
    assign dep_chan_data_23_0 = out_chan_dep_data_23;
    assign token_23_0 = token_out_vec_23[2];
    assign dep_chan_vld_23_2 = out_chan_dep_vld_vec_23[3];
    assign dep_chan_data_23_2 = out_chan_dep_data_23;
    assign token_23_2 = token_out_vec_23[3];
    assign dep_chan_vld_23_12 = out_chan_dep_vld_vec_23[4];
    assign dep_chan_data_23_12 = out_chan_dep_data_23;
    assign token_23_12 = token_out_vec_23[4];

    // Process: xfMat2Array_64_9_720_720_1_1_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 24, 3, 3) pp_pipeline_accel_hls_deadlock_detect_unit_24 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_24),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_24),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_24),
        .token_in_vec(token_in_vec_24),
        .dl_detect_in(dl_detect_out),
        .origin(origin[24]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_24),
        .out_chan_dep_data(out_chan_dep_data_24),
        .token_out_vec(token_out_vec_24),
        .dl_detect_out(dl_in_vec[24]));

    assign proc_24_data_FIFO_blk[0] = 1'b0 | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.MatStream2AxiStream_U0.out_mat_470_blk_n);
    assign proc_24_data_PIPO_blk[0] = 1'b0;
    assign proc_24_start_FIFO_blk[0] = 1'b0;
    assign proc_24_TLF_FIFO_blk[0] = 1'b0;
    assign proc_24_input_sync_blk[0] = 1'b0;
    assign proc_24_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_24[0] = dl_detect_out ? proc_dep_vld_vec_24_reg[0] : (proc_24_data_FIFO_blk[0] | proc_24_data_PIPO_blk[0] | proc_24_start_FIFO_blk[0] | proc_24_TLF_FIFO_blk[0] | proc_24_input_sync_blk[0] | proc_24_output_sync_blk[0]);
    assign proc_24_data_FIFO_blk[1] = 1'b0 | (~xfMat2Array_64_9_720_720_1_1_U0.srcMat_rows_blk_n) | (~xfMat2Array_64_9_720_720_1_1_U0.srcMat_cols_blk_n);
    assign proc_24_data_PIPO_blk[1] = 1'b0;
    assign proc_24_start_FIFO_blk[1] = 1'b0;
    assign proc_24_TLF_FIFO_blk[1] = 1'b0;
    assign proc_24_input_sync_blk[1] = 1'b0;
    assign proc_24_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_24[1] = dl_detect_out ? proc_dep_vld_vec_24_reg[1] : (proc_24_data_FIFO_blk[1] | proc_24_data_PIPO_blk[1] | proc_24_start_FIFO_blk[1] | proc_24_TLF_FIFO_blk[1] | proc_24_input_sync_blk[1] | proc_24_output_sync_blk[1]);
    assign proc_24_data_FIFO_blk[2] = 1'b0 | (~xfMat2Array_64_9_720_720_1_1_U0.dstPtr_blk_n) | (~xfMat2Array_64_9_720_720_1_1_U0.stride_blk_n);
    assign proc_24_data_PIPO_blk[2] = 1'b0;
    assign proc_24_start_FIFO_blk[2] = 1'b0 | (~start_for_xfMat2Array_64_9_720_720_1_1_U0_U.if_empty_n & xfMat2Array_64_9_720_720_1_1_U0.ap_idle & ~start_for_xfMat2Array_64_9_720_720_1_1_U0_U.if_write);
    assign proc_24_TLF_FIFO_blk[2] = 1'b0;
    assign proc_24_input_sync_blk[2] = 1'b0;
    assign proc_24_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_24[2] = dl_detect_out ? proc_dep_vld_vec_24_reg[2] : (proc_24_data_FIFO_blk[2] | proc_24_data_PIPO_blk[2] | proc_24_start_FIFO_blk[2] | proc_24_TLF_FIFO_blk[2] | proc_24_input_sync_blk[2] | proc_24_output_sync_blk[2]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_24_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_24_reg <= proc_dep_vld_vec_24;
        end
    end
    assign in_chan_dep_vld_vec_24[0] = dep_chan_vld_0_24;
    assign in_chan_dep_data_vec_24[32 : 0] = dep_chan_data_0_24;
    assign token_in_vec_24[0] = token_0_24;
    assign in_chan_dep_vld_vec_24[1] = dep_chan_vld_1_24;
    assign in_chan_dep_data_vec_24[65 : 33] = dep_chan_data_1_24;
    assign token_in_vec_24[1] = token_1_24;
    assign in_chan_dep_vld_vec_24[2] = dep_chan_vld_23_24;
    assign in_chan_dep_data_vec_24[98 : 66] = dep_chan_data_23_24;
    assign token_in_vec_24[2] = token_23_24;
    assign dep_chan_vld_24_23 = out_chan_dep_vld_vec_24[0];
    assign dep_chan_data_24_23 = out_chan_dep_data_24;
    assign token_24_23 = token_out_vec_24[0];
    assign dep_chan_vld_24_1 = out_chan_dep_vld_vec_24[1];
    assign dep_chan_data_24_1 = out_chan_dep_data_24;
    assign token_24_1 = token_out_vec_24[1];
    assign dep_chan_vld_24_0 = out_chan_dep_vld_vec_24[2];
    assign dep_chan_data_24_0 = out_chan_dep_data_24;
    assign token_24_0 = token_out_vec_24[2];

    // Process: xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 25, 4, 4) pp_pipeline_accel_hls_deadlock_detect_unit_25 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_25),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_25),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_25),
        .token_in_vec(token_in_vec_25),
        .dl_detect_in(dl_detect_out),
        .origin(origin[25]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_25),
        .out_chan_dep_data(out_chan_dep_data_25),
        .token_out_vec(token_out_vec_25),
        .dl_detect_out(dl_in_vec[25]));

    assign proc_25_data_FIFO_blk[0] = 1'b0 | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0.dout_out_blk_n);
    assign proc_25_data_PIPO_blk[0] = 1'b0;
    assign proc_25_start_FIFO_blk[0] = 1'b0;
    assign proc_25_TLF_FIFO_blk[0] = 1'b0;
    assign proc_25_input_sync_blk[0] = 1'b0;
    assign proc_25_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_25[0] = dl_detect_out ? proc_dep_vld_vec_25_reg[0] : (proc_25_data_FIFO_blk[0] | proc_25_data_PIPO_blk[0] | proc_25_start_FIFO_blk[0] | proc_25_TLF_FIFO_blk[0] | proc_25_input_sync_blk[0] | proc_25_output_sync_blk[0]);
    assign proc_25_data_FIFO_blk[1] = 1'b0 | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0.rows_out_blk_n) | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0.cols_out_blk_n) | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0.stride_out_blk_n);
    assign proc_25_data_PIPO_blk[1] = 1'b0;
    assign proc_25_start_FIFO_blk[1] = 1'b0 | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.start_for_Mat2Axi_Block_split2_proc_U0_U.if_full_n & xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0.ap_start & ~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0.real_start & (trans_in_cnt_9 == trans_out_cnt_9) & ~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.start_for_Mat2Axi_Block_split2_proc_U0_U.if_read);
    assign proc_25_TLF_FIFO_blk[1] = 1'b0;
    assign proc_25_input_sync_blk[1] = 1'b0;
    assign proc_25_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_25[1] = dl_detect_out ? proc_dep_vld_vec_25_reg[1] : (proc_25_data_FIFO_blk[1] | proc_25_data_PIPO_blk[1] | proc_25_start_FIFO_blk[1] | proc_25_TLF_FIFO_blk[1] | proc_25_input_sync_blk[1] | proc_25_output_sync_blk[1]);
    assign proc_25_data_FIFO_blk[2] = 1'b0 | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0.rows_out1_blk_n) | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0.cols_out2_blk_n) | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0.stride_out3_blk_n);
    assign proc_25_data_PIPO_blk[2] = 1'b0;
    assign proc_25_start_FIFO_blk[2] = 1'b0;
    assign proc_25_TLF_FIFO_blk[2] = 1'b0;
    assign proc_25_input_sync_blk[2] = 1'b0;
    assign proc_25_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_25[2] = dl_detect_out ? proc_dep_vld_vec_25_reg[2] : (proc_25_data_FIFO_blk[2] | proc_25_data_PIPO_blk[2] | proc_25_start_FIFO_blk[2] | proc_25_TLF_FIFO_blk[2] | proc_25_input_sync_blk[2] | proc_25_output_sync_blk[2]);
    assign proc_25_data_FIFO_blk[3] = 1'b0;
    assign proc_25_data_PIPO_blk[3] = 1'b0;
    assign proc_25_start_FIFO_blk[3] = 1'b0 | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.start_for_Mat2AxiStream_U0_U.if_full_n & xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0.ap_start & ~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_entry28_U0.real_start & (trans_in_cnt_9 == trans_out_cnt_9) & ~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.start_for_Mat2AxiStream_U0_U.if_read);
    assign proc_25_TLF_FIFO_blk[3] = 1'b0;
    assign proc_25_input_sync_blk[3] = 1'b0;
    assign proc_25_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_25[3] = dl_detect_out ? proc_dep_vld_vec_25_reg[3] : (proc_25_data_FIFO_blk[3] | proc_25_data_PIPO_blk[3] | proc_25_start_FIFO_blk[3] | proc_25_TLF_FIFO_blk[3] | proc_25_input_sync_blk[3] | proc_25_output_sync_blk[3]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_25_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_25_reg <= proc_dep_vld_vec_25;
        end
    end
    assign in_chan_dep_vld_vec_25[0] = dep_chan_vld_26_25;
    assign in_chan_dep_data_vec_25[32 : 0] = dep_chan_data_26_25;
    assign token_in_vec_25[0] = token_26_25;
    assign in_chan_dep_vld_vec_25[1] = dep_chan_vld_29_25;
    assign in_chan_dep_data_vec_25[65 : 33] = dep_chan_data_29_25;
    assign token_in_vec_25[1] = token_29_25;
    assign in_chan_dep_vld_vec_25[2] = dep_chan_vld_30_25;
    assign in_chan_dep_data_vec_25[98 : 66] = dep_chan_data_30_25;
    assign token_in_vec_25[2] = token_30_25;
    assign in_chan_dep_vld_vec_25[3] = dep_chan_vld_32_25;
    assign in_chan_dep_data_vec_25[131 : 99] = dep_chan_data_32_25;
    assign token_in_vec_25[3] = token_32_25;
    assign dep_chan_vld_25_32 = out_chan_dep_vld_vec_25[0];
    assign dep_chan_data_25_32 = out_chan_dep_data_25;
    assign token_25_32 = token_out_vec_25[0];
    assign dep_chan_vld_25_26 = out_chan_dep_vld_vec_25[1];
    assign dep_chan_data_25_26 = out_chan_dep_data_25;
    assign token_25_26 = token_out_vec_25[1];
    assign dep_chan_vld_25_30 = out_chan_dep_vld_vec_25[2];
    assign dep_chan_data_25_30 = out_chan_dep_data_25;
    assign token_25_30 = token_out_vec_25[2];
    assign dep_chan_vld_25_29 = out_chan_dep_vld_vec_25[3];
    assign dep_chan_data_25_29 = out_chan_dep_data_25;
    assign token_25_29 = token_out_vec_25[3];

    // Process: xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split2_proc_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 26, 2, 1) pp_pipeline_accel_hls_deadlock_detect_unit_26 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_26),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_26),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_26),
        .token_in_vec(token_in_vec_26),
        .dl_detect_in(dl_detect_out),
        .origin(origin[26]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_26),
        .out_chan_dep_data(out_chan_dep_data_26),
        .token_out_vec(token_out_vec_26),
        .dl_detect_out(dl_in_vec[26]));

    assign proc_26_data_FIFO_blk[0] = 1'b0 | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split2_proc_U0.stride_blk_n) | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split2_proc_U0.cols_blk_n) | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split2_proc_U0.rows_blk_n);
    assign proc_26_data_PIPO_blk[0] = 1'b0;
    assign proc_26_start_FIFO_blk[0] = 1'b0 | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.start_for_Mat2Axi_Block_split2_proc_U0_U.if_empty_n & xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split2_proc_U0.ap_idle & ~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.start_for_Mat2Axi_Block_split2_proc_U0_U.if_write);
    assign proc_26_TLF_FIFO_blk[0] = 1'b0;
    assign proc_26_input_sync_blk[0] = 1'b0;
    assign proc_26_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_26[0] = dl_detect_out ? proc_dep_vld_vec_26_reg[0] : (proc_26_data_FIFO_blk[0] | proc_26_data_PIPO_blk[0] | proc_26_start_FIFO_blk[0] | proc_26_TLF_FIFO_blk[0] | proc_26_input_sync_blk[0] | proc_26_output_sync_blk[0]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_26_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_26_reg <= proc_dep_vld_vec_26;
        end
    end
    assign in_chan_dep_vld_vec_26[0] = dep_chan_vld_25_26;
    assign in_chan_dep_data_vec_26[32 : 0] = dep_chan_data_25_26;
    assign token_in_vec_26[0] = token_25_26;
    assign in_chan_dep_vld_vec_26[1] = dep_chan_vld_27_26;
    assign in_chan_dep_data_vec_26[65 : 33] = dep_chan_data_27_26;
    assign token_in_vec_26[1] = token_27_26;
    assign dep_chan_vld_26_25 = out_chan_dep_vld_vec_26[0];
    assign dep_chan_data_26_25 = out_chan_dep_data_26;
    assign token_26_25 = token_out_vec_26[0];

    // Process: xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.addrbound_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 27, 1, 1) pp_pipeline_accel_hls_deadlock_detect_unit_27 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_27),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_27),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_27),
        .token_in_vec(token_in_vec_27),
        .dl_detect_in(dl_detect_out),
        .origin(origin[27]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_27),
        .out_chan_dep_data(out_chan_dep_data_27),
        .token_out_vec(token_out_vec_27),
        .dl_detect_out(dl_in_vec[27]));

    assign proc_27_data_FIFO_blk[0] = 1'b0;
    assign proc_27_data_PIPO_blk[0] = 1'b0;
    assign proc_27_start_FIFO_blk[0] = 1'b0;
    assign proc_27_TLF_FIFO_blk[0] = 1'b0 | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_cast_loc_channel_U.if_empty_n & xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.addrbound_U0.ap_idle & ~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.rows_cast_loc_channel_U.if_write) | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_tmp_loc_channel_U.if_empty_n & xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.addrbound_U0.ap_idle & ~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.cols_tmp_loc_channel_U.if_write);
    assign proc_27_input_sync_blk[0] = 1'b0;
    assign proc_27_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_27[0] = dl_detect_out ? proc_dep_vld_vec_27_reg[0] : (proc_27_data_FIFO_blk[0] | proc_27_data_PIPO_blk[0] | proc_27_start_FIFO_blk[0] | proc_27_TLF_FIFO_blk[0] | proc_27_input_sync_blk[0] | proc_27_output_sync_blk[0]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_27_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_27_reg <= proc_dep_vld_vec_27;
        end
    end
    assign in_chan_dep_vld_vec_27[0] = dep_chan_vld_28_27;
    assign in_chan_dep_data_vec_27[32 : 0] = dep_chan_data_28_27;
    assign token_in_vec_27[0] = token_28_27;
    assign dep_chan_vld_27_26 = out_chan_dep_vld_vec_27[0];
    assign dep_chan_data_27_26 = out_chan_dep_data_27;
    assign token_27_26 = token_out_vec_27[0];

    // Process: xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split24_proc_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 28, 1, 1) pp_pipeline_accel_hls_deadlock_detect_unit_28 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_28),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_28),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_28),
        .token_in_vec(token_in_vec_28),
        .dl_detect_in(dl_detect_out),
        .origin(origin[28]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_28),
        .out_chan_dep_data(out_chan_dep_data_28),
        .token_out_vec(token_out_vec_28),
        .dl_detect_out(dl_in_vec[28]));

    assign proc_28_data_FIFO_blk[0] = 1'b0;
    assign proc_28_data_PIPO_blk[0] = 1'b0;
    assign proc_28_start_FIFO_blk[0] = 1'b0;
    assign proc_28_TLF_FIFO_blk[0] = 1'b0 | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.p_channel_U.if_empty_n & xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2Axi_Block_split24_proc_U0.ap_idle & ~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.p_channel_U.if_write);
    assign proc_28_input_sync_blk[0] = 1'b0;
    assign proc_28_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_28[0] = dl_detect_out ? proc_dep_vld_vec_28_reg[0] : (proc_28_data_FIFO_blk[0] | proc_28_data_PIPO_blk[0] | proc_28_start_FIFO_blk[0] | proc_28_TLF_FIFO_blk[0] | proc_28_input_sync_blk[0] | proc_28_output_sync_blk[0]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_28_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_28_reg <= proc_dep_vld_vec_28;
        end
    end
    assign in_chan_dep_vld_vec_28[0] = dep_chan_vld_32_28;
    assign in_chan_dep_data_vec_28[32 : 0] = dep_chan_data_32_28;
    assign token_in_vec_28[0] = token_32_28;
    assign dep_chan_vld_28_27 = out_chan_dep_vld_vec_28[0];
    assign dep_chan_data_28_27 = out_chan_dep_data_28;
    assign token_28_27 = token_out_vec_28[0];

    // Process: xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 29, 1, 2) pp_pipeline_accel_hls_deadlock_detect_unit_29 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_29),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_29),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_29),
        .token_in_vec(token_in_vec_29),
        .dl_detect_in(dl_detect_out),
        .origin(origin[29]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_29),
        .out_chan_dep_data(out_chan_dep_data_29),
        .token_out_vec(token_out_vec_29),
        .dl_detect_out(dl_in_vec[29]));

    assign proc_29_data_FIFO_blk[0] = 1'b0 | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.MatStream2AxiStream_U0.ldata1_blk_n);
    assign proc_29_data_PIPO_blk[0] = 1'b0;
    assign proc_29_start_FIFO_blk[0] = 1'b0;
    assign proc_29_TLF_FIFO_blk[0] = 1'b0;
    assign proc_29_input_sync_blk[0] = 1'b0;
    assign proc_29_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_29[0] = dl_detect_out ? proc_dep_vld_vec_29_reg[0] : (proc_29_data_FIFO_blk[0] | proc_29_data_PIPO_blk[0] | proc_29_start_FIFO_blk[0] | proc_29_TLF_FIFO_blk[0] | proc_29_input_sync_blk[0] | proc_29_output_sync_blk[0]);
    assign proc_29_data_FIFO_blk[1] = 1'b0 | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0.rows_blk_n) | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0.cols_blk_n) | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0.stride_blk_n);
    assign proc_29_data_PIPO_blk[1] = 1'b0;
    assign proc_29_start_FIFO_blk[1] = 1'b0 | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.start_for_Mat2AxiStream_U0_U.if_empty_n & xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.ap_idle & ~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.start_for_Mat2AxiStream_U0_U.if_write);
    assign proc_29_TLF_FIFO_blk[1] = 1'b0;
    assign proc_29_input_sync_blk[1] = 1'b0;
    assign proc_29_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_29[1] = dl_detect_out ? proc_dep_vld_vec_29_reg[1] : (proc_29_data_FIFO_blk[1] | proc_29_data_PIPO_blk[1] | proc_29_start_FIFO_blk[1] | proc_29_TLF_FIFO_blk[1] | proc_29_input_sync_blk[1] | proc_29_output_sync_blk[1]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_29_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_29_reg <= proc_dep_vld_vec_29;
        end
    end
    assign in_chan_dep_vld_vec_29[0] = dep_chan_vld_25_29;
    assign in_chan_dep_data_vec_29[32 : 0] = dep_chan_data_25_29;
    assign token_in_vec_29[0] = token_25_29;
    assign dep_chan_vld_29_32 = out_chan_dep_vld_vec_29[0];
    assign dep_chan_data_29_32 = out_chan_dep_data_29;
    assign token_29_32 = token_out_vec_29[0];
    assign dep_chan_vld_29_25 = out_chan_dep_vld_vec_29[1];
    assign dep_chan_data_29_25 = out_chan_dep_data_29;
    assign token_29_25 = token_out_vec_29[1];

    // Process: xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 30, 2, 2) pp_pipeline_accel_hls_deadlock_detect_unit_30 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_30),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_30),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_30),
        .token_in_vec(token_in_vec_30),
        .dl_detect_in(dl_detect_out),
        .origin(origin[30]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_30),
        .out_chan_dep_data(out_chan_dep_data_30),
        .token_out_vec(token_out_vec_30),
        .dl_detect_out(dl_in_vec[30]));

    assign proc_30_data_FIFO_blk[0] = 1'b0 | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0.rows_blk_n) | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0.cols_blk_n) | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0.stride_blk_n);
    assign proc_30_data_PIPO_blk[0] = 1'b0;
    assign proc_30_start_FIFO_blk[0] = 1'b0;
    assign proc_30_TLF_FIFO_blk[0] = 1'b0;
    assign proc_30_input_sync_blk[0] = 1'b0;
    assign proc_30_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_30[0] = dl_detect_out ? proc_dep_vld_vec_30_reg[0] : (proc_30_data_FIFO_blk[0] | proc_30_data_PIPO_blk[0] | proc_30_start_FIFO_blk[0] | proc_30_TLF_FIFO_blk[0] | proc_30_input_sync_blk[0] | proc_30_output_sync_blk[0]);
    assign proc_30_data_FIFO_blk[1] = 1'b0 | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0.rows_out_blk_n) | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0.cols_out_blk_n) | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.last_blk_pxl_width25_U0.stride_out_blk_n);
    assign proc_30_data_PIPO_blk[1] = 1'b0;
    assign proc_30_start_FIFO_blk[1] = 1'b0;
    assign proc_30_TLF_FIFO_blk[1] = 1'b0;
    assign proc_30_input_sync_blk[1] = 1'b0;
    assign proc_30_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_30[1] = dl_detect_out ? proc_dep_vld_vec_30_reg[1] : (proc_30_data_FIFO_blk[1] | proc_30_data_PIPO_blk[1] | proc_30_start_FIFO_blk[1] | proc_30_TLF_FIFO_blk[1] | proc_30_input_sync_blk[1] | proc_30_output_sync_blk[1]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_30_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_30_reg <= proc_dep_vld_vec_30;
        end
    end
    assign in_chan_dep_vld_vec_30[0] = dep_chan_vld_25_30;
    assign in_chan_dep_data_vec_30[32 : 0] = dep_chan_data_25_30;
    assign token_in_vec_30[0] = token_25_30;
    assign in_chan_dep_vld_vec_30[1] = dep_chan_vld_31_30;
    assign in_chan_dep_data_vec_30[65 : 33] = dep_chan_data_31_30;
    assign token_in_vec_30[1] = token_31_30;
    assign dep_chan_vld_30_25 = out_chan_dep_vld_vec_30[0];
    assign dep_chan_data_30_25 = out_chan_dep_data_30;
    assign token_30_25 = token_out_vec_30[0];
    assign dep_chan_vld_30_31 = out_chan_dep_vld_vec_30[1];
    assign dep_chan_data_30_31 = out_chan_dep_data_30;
    assign token_30_31 = token_out_vec_30[1];

    // Process: xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.MatStream2AxiStream_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 31, 2, 2) pp_pipeline_accel_hls_deadlock_detect_unit_31 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_31),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_31),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_31),
        .token_in_vec(token_in_vec_31),
        .dl_detect_in(dl_detect_out),
        .origin(origin[31]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_31),
        .out_chan_dep_data(out_chan_dep_data_31),
        .token_out_vec(token_out_vec_31),
        .dl_detect_out(dl_in_vec[31]));

    assign proc_31_data_FIFO_blk[0] = 1'b0 | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.MatStream2AxiStream_U0.ldata1_blk_n);
    assign proc_31_data_PIPO_blk[0] = 1'b0;
    assign proc_31_start_FIFO_blk[0] = 1'b0;
    assign proc_31_TLF_FIFO_blk[0] = 1'b0;
    assign proc_31_input_sync_blk[0] = 1'b0;
    assign proc_31_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_31[0] = dl_detect_out ? proc_dep_vld_vec_31_reg[0] : (proc_31_data_FIFO_blk[0] | proc_31_data_PIPO_blk[0] | proc_31_start_FIFO_blk[0] | proc_31_TLF_FIFO_blk[0] | proc_31_input_sync_blk[0] | proc_31_output_sync_blk[0]);
    assign proc_31_data_FIFO_blk[1] = 1'b0 | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.MatStream2AxiStream_U0.rows_blk_n) | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.MatStream2AxiStream_U0.cols_bound_per_npc_blk_n) | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.MatStream2AxiStream_U0.stride_blk_n);
    assign proc_31_data_PIPO_blk[1] = 1'b0;
    assign proc_31_start_FIFO_blk[1] = 1'b0;
    assign proc_31_TLF_FIFO_blk[1] = 1'b0 | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.p_channel_U.if_empty_n & xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.MatStream2AxiStream_U0.ap_idle & ~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.Mat2AxiStream_U0.p_channel_U.if_write);
    assign proc_31_input_sync_blk[1] = 1'b0;
    assign proc_31_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_31[1] = dl_detect_out ? proc_dep_vld_vec_31_reg[1] : (proc_31_data_FIFO_blk[1] | proc_31_data_PIPO_blk[1] | proc_31_start_FIFO_blk[1] | proc_31_TLF_FIFO_blk[1] | proc_31_input_sync_blk[1] | proc_31_output_sync_blk[1]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_31_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_31_reg <= proc_dep_vld_vec_31;
        end
    end
    assign in_chan_dep_vld_vec_31[0] = dep_chan_vld_30_31;
    assign in_chan_dep_data_vec_31[32 : 0] = dep_chan_data_30_31;
    assign token_in_vec_31[0] = token_30_31;
    assign in_chan_dep_vld_vec_31[1] = dep_chan_vld_32_31;
    assign in_chan_dep_data_vec_31[65 : 33] = dep_chan_data_32_31;
    assign token_in_vec_31[1] = token_32_31;
    assign dep_chan_vld_31_32 = out_chan_dep_vld_vec_31[0];
    assign dep_chan_data_31_32 = out_chan_dep_data_31;
    assign token_31_32 = token_out_vec_31[0];
    assign dep_chan_vld_31_30 = out_chan_dep_vld_vec_31[1];
    assign dep_chan_data_31_30 = out_chan_dep_data_31;
    assign token_31_30 = token_out_vec_31[1];

    // Process: xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.AxiStream2Axi_U0
    pp_pipeline_accel_hls_deadlock_detect_unit #(33, 32, 3, 3) pp_pipeline_accel_hls_deadlock_detect_unit_32 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_32),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_32),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_32),
        .token_in_vec(token_in_vec_32),
        .dl_detect_in(dl_detect_out),
        .origin(origin[32]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_32),
        .out_chan_dep_data(out_chan_dep_data_32),
        .token_out_vec(token_out_vec_32),
        .dl_detect_out(dl_in_vec[32]));

    assign proc_32_data_FIFO_blk[0] = 1'b0 | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.AxiStream2Axi_U0.ldata1_blk_n);
    assign proc_32_data_PIPO_blk[0] = 1'b0;
    assign proc_32_start_FIFO_blk[0] = 1'b0;
    assign proc_32_TLF_FIFO_blk[0] = 1'b0;
    assign proc_32_input_sync_blk[0] = 1'b0;
    assign proc_32_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_32[0] = dl_detect_out ? proc_dep_vld_vec_32_reg[0] : (proc_32_data_FIFO_blk[0] | proc_32_data_PIPO_blk[0] | proc_32_start_FIFO_blk[0] | proc_32_TLF_FIFO_blk[0] | proc_32_input_sync_blk[0] | proc_32_output_sync_blk[0]);
    assign proc_32_data_FIFO_blk[1] = 1'b0 | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.AxiStream2Axi_U0.dout_blk_n);
    assign proc_32_data_PIPO_blk[1] = 1'b0;
    assign proc_32_start_FIFO_blk[1] = 1'b0;
    assign proc_32_TLF_FIFO_blk[1] = 1'b0;
    assign proc_32_input_sync_blk[1] = 1'b0;
    assign proc_32_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_32[1] = dl_detect_out ? proc_dep_vld_vec_32_reg[1] : (proc_32_data_FIFO_blk[1] | proc_32_data_PIPO_blk[1] | proc_32_start_FIFO_blk[1] | proc_32_TLF_FIFO_blk[1] | proc_32_input_sync_blk[1] | proc_32_output_sync_blk[1]);
    assign proc_32_data_FIFO_blk[2] = 1'b0;
    assign proc_32_data_PIPO_blk[2] = 1'b0;
    assign proc_32_start_FIFO_blk[2] = 1'b0;
    assign proc_32_TLF_FIFO_blk[2] = 1'b0 | (~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.axibound_V_U.if_empty_n & xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.AxiStream2Axi_U0.ap_idle & ~xfMat2Array_64_9_720_720_1_1_U0.grp_Mat2Axi_fu_68.axibound_V_U.if_write);
    assign proc_32_input_sync_blk[2] = 1'b0;
    assign proc_32_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_32[2] = dl_detect_out ? proc_dep_vld_vec_32_reg[2] : (proc_32_data_FIFO_blk[2] | proc_32_data_PIPO_blk[2] | proc_32_start_FIFO_blk[2] | proc_32_TLF_FIFO_blk[2] | proc_32_input_sync_blk[2] | proc_32_output_sync_blk[2]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_32_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_32_reg <= proc_dep_vld_vec_32;
        end
    end
    assign in_chan_dep_vld_vec_32[0] = dep_chan_vld_25_32;
    assign in_chan_dep_data_vec_32[32 : 0] = dep_chan_data_25_32;
    assign token_in_vec_32[0] = token_25_32;
    assign in_chan_dep_vld_vec_32[1] = dep_chan_vld_29_32;
    assign in_chan_dep_data_vec_32[65 : 33] = dep_chan_data_29_32;
    assign token_in_vec_32[1] = token_29_32;
    assign in_chan_dep_vld_vec_32[2] = dep_chan_vld_31_32;
    assign in_chan_dep_data_vec_32[98 : 66] = dep_chan_data_31_32;
    assign token_in_vec_32[2] = token_31_32;
    assign dep_chan_vld_32_31 = out_chan_dep_vld_vec_32[0];
    assign dep_chan_data_32_31 = out_chan_dep_data_32;
    assign token_32_31 = token_out_vec_32[0];
    assign dep_chan_vld_32_25 = out_chan_dep_vld_vec_32[1];
    assign dep_chan_data_32_25 = out_chan_dep_data_32;
    assign token_32_25 = token_out_vec_32[1];
    assign dep_chan_vld_32_28 = out_chan_dep_vld_vec_32[2];
    assign dep_chan_data_32_28 = out_chan_dep_data_32;
    assign token_32_28 = token_out_vec_32[2];


`include "pp_pipeline_accel_hls_deadlock_report_unit.vh"
