// Copyright (C) 2022, Advanced Micro Devices, Inc. All rights reserved.
// SPDX-License-Identifier: MIT
// ==============================================================
// Version: 2022.1
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module pp_pipeline_accel_resize_1_9_2160_3840_720_720_1_9_s (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        p_read,
        p_read1,
        rgb_mat_data83_dout,
        rgb_mat_data83_num_data_valid,
        rgb_mat_data83_fifo_cap,
        rgb_mat_data83_empty_n,
        rgb_mat_data83_read,
        p_read2,
        p_read3,
        resize_out_mat_data84_din,
        resize_out_mat_data84_num_data_valid,
        resize_out_mat_data84_fifo_cap,
        resize_out_mat_data84_full_n,
        resize_out_mat_data84_write,
        resize_out_mat_rows_c_din,
        resize_out_mat_rows_c_num_data_valid,
        resize_out_mat_rows_c_fifo_cap,
        resize_out_mat_rows_c_full_n,
        resize_out_mat_rows_c_write,
        resize_out_mat_cols_c_din,
        resize_out_mat_cols_c_num_data_valid,
        resize_out_mat_cols_c_fifo_cap,
        resize_out_mat_cols_c_full_n,
        resize_out_mat_cols_c_write
);

parameter    ap_ST_fsm_state1 = 2'd1;
parameter    ap_ST_fsm_state2 = 2'd2;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [31:0] p_read;
input  [31:0] p_read1;
input  [23:0] rgb_mat_data83_dout;
input  [1:0] rgb_mat_data83_num_data_valid;
input  [1:0] rgb_mat_data83_fifo_cap;
input   rgb_mat_data83_empty_n;
output   rgb_mat_data83_read;
input  [31:0] p_read2;
input  [31:0] p_read3;
output  [23:0] resize_out_mat_data84_din;
input  [1:0] resize_out_mat_data84_num_data_valid;
input  [1:0] resize_out_mat_data84_fifo_cap;
input   resize_out_mat_data84_full_n;
output   resize_out_mat_data84_write;
output  [31:0] resize_out_mat_rows_c_din;
input  [1:0] resize_out_mat_rows_c_num_data_valid;
input  [1:0] resize_out_mat_rows_c_fifo_cap;
input   resize_out_mat_rows_c_full_n;
output   resize_out_mat_rows_c_write;
output  [31:0] resize_out_mat_cols_c_din;
input  [1:0] resize_out_mat_cols_c_num_data_valid;
input  [1:0] resize_out_mat_cols_c_fifo_cap;
input   resize_out_mat_cols_c_full_n;
output   resize_out_mat_cols_c_write;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg rgb_mat_data83_read;
reg resize_out_mat_data84_write;
reg resize_out_mat_rows_c_write;
reg resize_out_mat_cols_c_write;

reg    ap_done_reg;
(* fsm_encoding = "none" *) reg   [1:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    resize_out_mat_rows_c_blk_n;
reg    resize_out_mat_cols_c_blk_n;
wire    grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_ap_start;
wire    grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_ap_done;
wire    grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_ap_idle;
wire    grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_ap_ready;
wire    grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_rgb_mat_data83_read;
wire   [23:0] grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_resize_out_mat_data84_din;
wire    grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_resize_out_mat_data84_write;
reg    grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_ap_start_reg;
reg    ap_block_state1_ignore_call10;
wire    ap_CS_fsm_state2;
reg    ap_block_state1;
reg   [1:0] ap_NS_fsm;
reg    ap_ST_fsm_state1_blk;
reg    ap_ST_fsm_state2_blk;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 2'd1;
#0 grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_ap_start_reg = 1'b0;
end

pp_pipeline_accel_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_ap_start),
    .ap_done(grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_ap_done),
    .ap_idle(grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_ap_idle),
    .ap_ready(grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_ap_ready),
    .p_read(p_read),
    .p_read1(p_read1),
    .rgb_mat_data83_dout(rgb_mat_data83_dout),
    .rgb_mat_data83_num_data_valid(2'd0),
    .rgb_mat_data83_fifo_cap(2'd0),
    .rgb_mat_data83_empty_n(rgb_mat_data83_empty_n),
    .rgb_mat_data83_read(grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_rgb_mat_data83_read),
    .p_read2(p_read2),
    .p_read3(p_read3),
    .resize_out_mat_data84_din(grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_resize_out_mat_data84_din),
    .resize_out_mat_data84_num_data_valid(2'd0),
    .resize_out_mat_data84_fifo_cap(2'd0),
    .resize_out_mat_data84_full_n(resize_out_mat_data84_full_n),
    .resize_out_mat_data84_write(grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_resize_out_mat_data84_write)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state2))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_ap_start_reg <= 1'b0;
    end else begin
        if ((~((ap_start == 1'b0) | (resize_out_mat_cols_c_full_n == 1'b0) | (resize_out_mat_rows_c_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_ap_start_reg <= 1'b1;
        end else if ((grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_ap_ready == 1'b1)) begin
            grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_ap_start_reg <= 1'b0;
        end
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) | (resize_out_mat_cols_c_full_n == 1'b0) | (resize_out_mat_rows_c_full_n == 1'b0) | (ap_done_reg == 1'b1))) begin
        ap_ST_fsm_state1_blk = 1'b1;
    end else begin
        ap_ST_fsm_state1_blk = 1'b0;
    end
end

always @ (*) begin
    if ((grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_ap_done == 1'b0)) begin
        ap_ST_fsm_state2_blk = 1'b1;
    end else begin
        ap_ST_fsm_state2_blk = 1'b0;
    end
end

always @ (*) begin
    if (((grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        resize_out_mat_cols_c_blk_n = resize_out_mat_cols_c_full_n;
    end else begin
        resize_out_mat_cols_c_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (resize_out_mat_cols_c_full_n == 1'b0) | (resize_out_mat_rows_c_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        resize_out_mat_cols_c_write = 1'b1;
    end else begin
        resize_out_mat_cols_c_write = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        resize_out_mat_data84_write = grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_resize_out_mat_data84_write;
    end else begin
        resize_out_mat_data84_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        resize_out_mat_rows_c_blk_n = resize_out_mat_rows_c_full_n;
    end else begin
        resize_out_mat_rows_c_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (resize_out_mat_cols_c_full_n == 1'b0) | (resize_out_mat_rows_c_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        resize_out_mat_rows_c_write = 1'b1;
    end else begin
        resize_out_mat_rows_c_write = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        rgb_mat_data83_read = grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_rgb_mat_data83_read;
    end else begin
        rgb_mat_data83_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (resize_out_mat_cols_c_full_n == 1'b0) | (resize_out_mat_rows_c_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            if (((grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state2))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (resize_out_mat_cols_c_full_n == 1'b0) | (resize_out_mat_rows_c_full_n == 1'b0) | (ap_done_reg == 1'b1));
end

always @ (*) begin
    ap_block_state1_ignore_call10 = ((ap_start == 1'b0) | (resize_out_mat_cols_c_full_n == 1'b0) | (resize_out_mat_rows_c_full_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_ap_start = grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_ap_start_reg;

assign resize_out_mat_cols_c_din = p_read3;

assign resize_out_mat_data84_din = grp_resizeNNBilinear_9_2160_3840_1_720_720_1_9_s_fu_82_resize_out_mat_data84_din;

assign resize_out_mat_rows_c_din = p_read2;

endmodule //pp_pipeline_accel_resize_1_9_2160_3840_720_720_1_9_s
